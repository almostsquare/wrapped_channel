// This is the unpowered netlist.
module wrapped_channel (active,
    wb_clk_i,
    io_in,
    io_oeb,
    io_out,
    la1_data_in,
    la1_data_out,
    la1_oenb);
 input active;
 input wb_clk_i;
 input [37:0] io_in;
 inout [37:0] io_oeb;
 inout [37:0] io_out;
 input [31:0] la1_data_in;
 inout [31:0] la1_data_out;
 input [31:0] la1_oenb;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire clknet_0_wb_clk_i;
 wire \gps_channel0.ca_full_chip ;
 wire \gps_channel0.ca_gen.g1[10] ;
 wire \gps_channel0.ca_gen.g1[1] ;
 wire \gps_channel0.ca_gen.g1[2] ;
 wire \gps_channel0.ca_gen.g1[3] ;
 wire \gps_channel0.ca_gen.g1[4] ;
 wire \gps_channel0.ca_gen.g1[5] ;
 wire \gps_channel0.ca_gen.g1[6] ;
 wire \gps_channel0.ca_gen.g1[7] ;
 wire \gps_channel0.ca_gen.g1[8] ;
 wire \gps_channel0.ca_gen.g1[9] ;
 wire \gps_channel0.ca_gen.g2[10] ;
 wire \gps_channel0.ca_gen.g2[1] ;
 wire \gps_channel0.ca_gen.g2[2] ;
 wire \gps_channel0.ca_gen.g2[3] ;
 wire \gps_channel0.ca_gen.g2[4] ;
 wire \gps_channel0.ca_gen.g2[5] ;
 wire \gps_channel0.ca_gen.g2[6] ;
 wire \gps_channel0.ca_gen.g2[7] ;
 wire \gps_channel0.ca_gen.g2[8] ;
 wire \gps_channel0.ca_gen.g2[9] ;
 wire \gps_channel0.ca_gen.g2_init[10] ;
 wire \gps_channel0.ca_gen.g2_init[1] ;
 wire \gps_channel0.ca_gen.g2_init[2] ;
 wire \gps_channel0.ca_gen.g2_init[3] ;
 wire \gps_channel0.ca_gen.g2_init[4] ;
 wire \gps_channel0.ca_gen.g2_init[5] ;
 wire \gps_channel0.ca_gen.g2_init[6] ;
 wire \gps_channel0.ca_gen.g2_init[7] ;
 wire \gps_channel0.ca_gen.g2_init[8] ;
 wire \gps_channel0.ca_gen.g2_init[9] ;
 wire \gps_channel0.ca_nco.accumulator[0] ;
 wire \gps_channel0.ca_nco.accumulator[10] ;
 wire \gps_channel0.ca_nco.accumulator[11] ;
 wire \gps_channel0.ca_nco.accumulator[12] ;
 wire \gps_channel0.ca_nco.accumulator[13] ;
 wire \gps_channel0.ca_nco.accumulator[14] ;
 wire \gps_channel0.ca_nco.accumulator[15] ;
 wire \gps_channel0.ca_nco.accumulator[16] ;
 wire \gps_channel0.ca_nco.accumulator[17] ;
 wire \gps_channel0.ca_nco.accumulator[18] ;
 wire \gps_channel0.ca_nco.accumulator[19] ;
 wire \gps_channel0.ca_nco.accumulator[1] ;
 wire \gps_channel0.ca_nco.accumulator[20] ;
 wire \gps_channel0.ca_nco.accumulator[21] ;
 wire \gps_channel0.ca_nco.accumulator[22] ;
 wire \gps_channel0.ca_nco.accumulator[23] ;
 wire \gps_channel0.ca_nco.accumulator[24] ;
 wire \gps_channel0.ca_nco.accumulator[25] ;
 wire \gps_channel0.ca_nco.accumulator[26] ;
 wire \gps_channel0.ca_nco.accumulator[27] ;
 wire \gps_channel0.ca_nco.accumulator[28] ;
 wire \gps_channel0.ca_nco.accumulator[29] ;
 wire \gps_channel0.ca_nco.accumulator[2] ;
 wire \gps_channel0.ca_nco.accumulator[30] ;
 wire \gps_channel0.ca_nco.accumulator[3] ;
 wire \gps_channel0.ca_nco.accumulator[4] ;
 wire \gps_channel0.ca_nco.accumulator[5] ;
 wire \gps_channel0.ca_nco.accumulator[6] ;
 wire \gps_channel0.ca_nco.accumulator[7] ;
 wire \gps_channel0.ca_nco.accumulator[8] ;
 wire \gps_channel0.ca_nco.accumulator[9] ;
 wire \gps_channel0.ca_nco.phase_in[0] ;
 wire \gps_channel0.ca_nco.phase_in[10] ;
 wire \gps_channel0.ca_nco.phase_in[11] ;
 wire \gps_channel0.ca_nco.phase_in[12] ;
 wire \gps_channel0.ca_nco.phase_in[13] ;
 wire \gps_channel0.ca_nco.phase_in[14] ;
 wire \gps_channel0.ca_nco.phase_in[15] ;
 wire \gps_channel0.ca_nco.phase_in[1] ;
 wire \gps_channel0.ca_nco.phase_in[2] ;
 wire \gps_channel0.ca_nco.phase_in[3] ;
 wire \gps_channel0.ca_nco.phase_in[4] ;
 wire \gps_channel0.ca_nco.phase_in[5] ;
 wire \gps_channel0.ca_nco.phase_in[6] ;
 wire \gps_channel0.ca_nco.phase_in[7] ;
 wire \gps_channel0.ca_nco.phase_in[8] ;
 wire \gps_channel0.ca_nco.phase_in[9] ;
 wire \gps_channel0.ca_nco.phase_sync ;
 wire \gps_channel0.ca_nco.step[0] ;
 wire \gps_channel0.ca_nco.step[10] ;
 wire \gps_channel0.ca_nco.step[11] ;
 wire \gps_channel0.ca_nco.step[12] ;
 wire \gps_channel0.ca_nco.step[13] ;
 wire \gps_channel0.ca_nco.step[14] ;
 wire \gps_channel0.ca_nco.step[15] ;
 wire \gps_channel0.ca_nco.step[16] ;
 wire \gps_channel0.ca_nco.step[1] ;
 wire \gps_channel0.ca_nco.step[2] ;
 wire \gps_channel0.ca_nco.step[3] ;
 wire \gps_channel0.ca_nco.step[4] ;
 wire \gps_channel0.ca_nco.step[5] ;
 wire \gps_channel0.ca_nco.step[6] ;
 wire \gps_channel0.ca_nco.step[7] ;
 wire \gps_channel0.ca_nco.step[8] ;
 wire \gps_channel0.ca_nco.step[9] ;
 wire \gps_channel0.lo_i ;
 wire \gps_channel0.lo_nco.accumulator[0] ;
 wire \gps_channel0.lo_nco.accumulator[10] ;
 wire \gps_channel0.lo_nco.accumulator[11] ;
 wire \gps_channel0.lo_nco.accumulator[12] ;
 wire \gps_channel0.lo_nco.accumulator[13] ;
 wire \gps_channel0.lo_nco.accumulator[14] ;
 wire \gps_channel0.lo_nco.accumulator[15] ;
 wire \gps_channel0.lo_nco.accumulator[16] ;
 wire \gps_channel0.lo_nco.accumulator[17] ;
 wire \gps_channel0.lo_nco.accumulator[18] ;
 wire \gps_channel0.lo_nco.accumulator[19] ;
 wire \gps_channel0.lo_nco.accumulator[1] ;
 wire \gps_channel0.lo_nco.accumulator[20] ;
 wire \gps_channel0.lo_nco.accumulator[21] ;
 wire \gps_channel0.lo_nco.accumulator[22] ;
 wire \gps_channel0.lo_nco.accumulator[23] ;
 wire \gps_channel0.lo_nco.accumulator[24] ;
 wire \gps_channel0.lo_nco.accumulator[25] ;
 wire \gps_channel0.lo_nco.accumulator[26] ;
 wire \gps_channel0.lo_nco.accumulator[27] ;
 wire \gps_channel0.lo_nco.accumulator[28] ;
 wire \gps_channel0.lo_nco.accumulator[29] ;
 wire \gps_channel0.lo_nco.accumulator[2] ;
 wire \gps_channel0.lo_nco.accumulator[30] ;
 wire \gps_channel0.lo_nco.accumulator[3] ;
 wire \gps_channel0.lo_nco.accumulator[4] ;
 wire \gps_channel0.lo_nco.accumulator[5] ;
 wire \gps_channel0.lo_nco.accumulator[6] ;
 wire \gps_channel0.lo_nco.accumulator[7] ;
 wire \gps_channel0.lo_nco.accumulator[8] ;
 wire \gps_channel0.lo_nco.accumulator[9] ;
 wire \gps_channel0.lo_nco.phase_in[0] ;
 wire \gps_channel0.lo_nco.phase_in[10] ;
 wire \gps_channel0.lo_nco.phase_in[11] ;
 wire \gps_channel0.lo_nco.phase_in[12] ;
 wire \gps_channel0.lo_nco.phase_in[13] ;
 wire \gps_channel0.lo_nco.phase_in[14] ;
 wire \gps_channel0.lo_nco.phase_in[15] ;
 wire \gps_channel0.lo_nco.phase_in[1] ;
 wire \gps_channel0.lo_nco.phase_in[2] ;
 wire \gps_channel0.lo_nco.phase_in[3] ;
 wire \gps_channel0.lo_nco.phase_in[4] ;
 wire \gps_channel0.lo_nco.phase_in[5] ;
 wire \gps_channel0.lo_nco.phase_in[6] ;
 wire \gps_channel0.lo_nco.phase_in[7] ;
 wire \gps_channel0.lo_nco.phase_in[8] ;
 wire \gps_channel0.lo_nco.phase_in[9] ;
 wire \gps_channel0.lo_nco.phase_sync ;
 wire \gps_channel0.lo_nco.step[0] ;
 wire \gps_channel0.lo_nco.step[10] ;
 wire \gps_channel0.lo_nco.step[11] ;
 wire \gps_channel0.lo_nco.step[12] ;
 wire \gps_channel0.lo_nco.step[13] ;
 wire \gps_channel0.lo_nco.step[14] ;
 wire \gps_channel0.lo_nco.step[15] ;
 wire \gps_channel0.lo_nco.step[16] ;
 wire \gps_channel0.lo_nco.step[1] ;
 wire \gps_channel0.lo_nco.step[2] ;
 wire \gps_channel0.lo_nco.step[3] ;
 wire \gps_channel0.lo_nco.step[4] ;
 wire \gps_channel0.lo_nco.step[5] ;
 wire \gps_channel0.lo_nco.step[6] ;
 wire \gps_channel0.lo_nco.step[7] ;
 wire \gps_channel0.lo_nco.step[8] ;
 wire \gps_channel0.lo_nco.step[9] ;
 wire \gps_channel0.prompt_i ;
 wire \gps_channel0.prompt_q ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire clknet_4_0_0_wb_clk_i;
 wire clknet_4_1_0_wb_clk_i;
 wire clknet_4_2_0_wb_clk_i;
 wire clknet_4_3_0_wb_clk_i;
 wire clknet_4_4_0_wb_clk_i;
 wire clknet_4_5_0_wb_clk_i;
 wire clknet_4_6_0_wb_clk_i;
 wire clknet_4_7_0_wb_clk_i;
 wire clknet_4_8_0_wb_clk_i;
 wire clknet_4_9_0_wb_clk_i;
 wire clknet_4_10_0_wb_clk_i;
 wire clknet_4_11_0_wb_clk_i;
 wire clknet_4_12_0_wb_clk_i;
 wire clknet_4_13_0_wb_clk_i;
 wire clknet_4_14_0_wb_clk_i;
 wire clknet_4_15_0_wb_clk_i;

 sky130_fd_sc_hd__buf_6 _0951_ (.A(net1),
    .X(_0374_));
 sky130_fd_sc_hd__buf_8 _0952_ (.A(_0374_),
    .X(_0375_));
 sky130_fd_sc_hd__buf_8 _0953_ (.A(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__inv_2 _0954_ (.A(_0376_),
    .Y(_0787_));
 sky130_fd_sc_hd__inv_2 _0955_ (.A(_0376_),
    .Y(_0788_));
 sky130_fd_sc_hd__inv_2 _0956_ (.A(_0376_),
    .Y(_0789_));
 sky130_fd_sc_hd__inv_2 _0957_ (.A(_0376_),
    .Y(_0790_));
 sky130_fd_sc_hd__inv_2 _0958_ (.A(_0376_),
    .Y(_0791_));
 sky130_fd_sc_hd__inv_2 _0959_ (.A(_0376_),
    .Y(_0792_));
 sky130_fd_sc_hd__inv_2 _0960_ (.A(_0376_),
    .Y(_0793_));
 sky130_fd_sc_hd__inv_2 _0961_ (.A(_0376_),
    .Y(_0794_));
 sky130_fd_sc_hd__inv_2 _0962_ (.A(_0376_),
    .Y(_0795_));
 sky130_fd_sc_hd__inv_2 _0963_ (.A(_0376_),
    .Y(_0796_));
 sky130_fd_sc_hd__buf_8 _0964_ (.A(_0375_),
    .X(_0377_));
 sky130_fd_sc_hd__inv_2 _0965_ (.A(_0377_),
    .Y(_0797_));
 sky130_fd_sc_hd__inv_2 _0966_ (.A(_0377_),
    .Y(_0798_));
 sky130_fd_sc_hd__inv_2 _0967_ (.A(_0377_),
    .Y(_0799_));
 sky130_fd_sc_hd__inv_2 _0968_ (.A(_0377_),
    .Y(_0800_));
 sky130_fd_sc_hd__inv_2 _0969_ (.A(_0377_),
    .Y(_0801_));
 sky130_fd_sc_hd__inv_2 _0970_ (.A(_0377_),
    .Y(_0802_));
 sky130_fd_sc_hd__inv_2 _0971_ (.A(_0377_),
    .Y(_0803_));
 sky130_fd_sc_hd__inv_2 _0972_ (.A(_0377_),
    .Y(_0804_));
 sky130_fd_sc_hd__inv_2 _0973_ (.A(_0377_),
    .Y(_0805_));
 sky130_fd_sc_hd__inv_2 _0974_ (.A(_0377_),
    .Y(_0806_));
 sky130_fd_sc_hd__buf_8 _0975_ (.A(_0374_),
    .X(_0378_));
 sky130_fd_sc_hd__inv_2 _0976_ (.A(_0378_),
    .Y(_0807_));
 sky130_fd_sc_hd__inv_2 _0977_ (.A(_0378_),
    .Y(_0808_));
 sky130_fd_sc_hd__inv_2 _0978_ (.A(_0378_),
    .Y(_0809_));
 sky130_fd_sc_hd__inv_2 _0979_ (.A(_0378_),
    .Y(_0810_));
 sky130_fd_sc_hd__inv_2 _0980_ (.A(_0378_),
    .Y(_0811_));
 sky130_fd_sc_hd__inv_2 _0981_ (.A(_0378_),
    .Y(_0812_));
 sky130_fd_sc_hd__inv_2 _0982_ (.A(_0378_),
    .Y(_0813_));
 sky130_fd_sc_hd__inv_2 _0983_ (.A(_0378_),
    .Y(_0814_));
 sky130_fd_sc_hd__inv_2 _0984_ (.A(_0378_),
    .Y(_0815_));
 sky130_fd_sc_hd__inv_2 _0985_ (.A(_0378_),
    .Y(_0817_));
 sky130_fd_sc_hd__clkbuf_16 _0986_ (.A(_0374_),
    .X(_0379_));
 sky130_fd_sc_hd__inv_2 _0987_ (.A(_0379_),
    .Y(_0818_));
 sky130_fd_sc_hd__inv_2 _0988_ (.A(_0379_),
    .Y(_0819_));
 sky130_fd_sc_hd__inv_2 _0989_ (.A(_0379_),
    .Y(_0820_));
 sky130_fd_sc_hd__inv_2 _0990_ (.A(_0379_),
    .Y(_0821_));
 sky130_fd_sc_hd__inv_2 _0991_ (.A(_0379_),
    .Y(_0822_));
 sky130_fd_sc_hd__inv_2 _0992_ (.A(_0379_),
    .Y(_0823_));
 sky130_fd_sc_hd__inv_2 _0993_ (.A(_0379_),
    .Y(_0824_));
 sky130_fd_sc_hd__inv_2 _0994_ (.A(_0379_),
    .Y(_0825_));
 sky130_fd_sc_hd__inv_2 _0995_ (.A(_0379_),
    .Y(_0826_));
 sky130_fd_sc_hd__inv_2 _0996_ (.A(_0379_),
    .Y(_0827_));
 sky130_fd_sc_hd__buf_8 _0997_ (.A(_0374_),
    .X(_0380_));
 sky130_fd_sc_hd__inv_2 _0998_ (.A(_0380_),
    .Y(_0828_));
 sky130_fd_sc_hd__inv_2 _0999_ (.A(_0380_),
    .Y(_0829_));
 sky130_fd_sc_hd__inv_2 _1000_ (.A(_0380_),
    .Y(_0830_));
 sky130_fd_sc_hd__inv_2 _1001_ (.A(_0380_),
    .Y(_0831_));
 sky130_fd_sc_hd__inv_2 _1002_ (.A(_0380_),
    .Y(_0832_));
 sky130_fd_sc_hd__inv_2 _1003_ (.A(_0380_),
    .Y(_0833_));
 sky130_fd_sc_hd__inv_2 _1004_ (.A(_0380_),
    .Y(_0834_));
 sky130_fd_sc_hd__inv_2 _1005_ (.A(_0380_),
    .Y(_0835_));
 sky130_fd_sc_hd__inv_2 _1006_ (.A(_0380_),
    .Y(_0836_));
 sky130_fd_sc_hd__inv_2 _1007_ (.A(_0380_),
    .Y(_0837_));
 sky130_fd_sc_hd__buf_8 _1008_ (.A(_0374_),
    .X(_0381_));
 sky130_fd_sc_hd__inv_2 _1009_ (.A(_0381_),
    .Y(_0838_));
 sky130_fd_sc_hd__inv_2 _1010_ (.A(_0381_),
    .Y(_0839_));
 sky130_fd_sc_hd__inv_2 _1011_ (.A(_0381_),
    .Y(_0840_));
 sky130_fd_sc_hd__inv_2 _1012_ (.A(_0381_),
    .Y(_0841_));
 sky130_fd_sc_hd__inv_2 _1013_ (.A(_0381_),
    .Y(_0842_));
 sky130_fd_sc_hd__inv_2 _1014_ (.A(_0381_),
    .Y(_0843_));
 sky130_fd_sc_hd__inv_2 _1015_ (.A(_0381_),
    .Y(_0844_));
 sky130_fd_sc_hd__inv_2 _1016_ (.A(_0381_),
    .Y(_0845_));
 sky130_fd_sc_hd__inv_2 _1017_ (.A(_0381_),
    .Y(_0846_));
 sky130_fd_sc_hd__inv_2 _1018_ (.A(_0381_),
    .Y(_0847_));
 sky130_fd_sc_hd__buf_6 _1019_ (.A(_0374_),
    .X(_0382_));
 sky130_fd_sc_hd__inv_2 _1020_ (.A(_0382_),
    .Y(_0848_));
 sky130_fd_sc_hd__inv_2 _1021_ (.A(_0382_),
    .Y(_0849_));
 sky130_fd_sc_hd__inv_2 _1022_ (.A(_0382_),
    .Y(_0746_));
 sky130_fd_sc_hd__inv_2 _1023_ (.A(_0382_),
    .Y(_0850_));
 sky130_fd_sc_hd__inv_2 _1024_ (.A(_0382_),
    .Y(_0747_));
 sky130_fd_sc_hd__inv_2 _1025_ (.A(_0382_),
    .Y(_0851_));
 sky130_fd_sc_hd__inv_2 _1026_ (.A(_0382_),
    .Y(_0748_));
 sky130_fd_sc_hd__inv_2 _1027_ (.A(_0382_),
    .Y(_0852_));
 sky130_fd_sc_hd__inv_2 _1028_ (.A(_0382_),
    .Y(_0749_));
 sky130_fd_sc_hd__inv_2 _1029_ (.A(_0382_),
    .Y(_0853_));
 sky130_fd_sc_hd__buf_8 _1030_ (.A(_0374_),
    .X(_0383_));
 sky130_fd_sc_hd__inv_2 _1031_ (.A(_0383_),
    .Y(_0750_));
 sky130_fd_sc_hd__inv_2 _1032_ (.A(_0383_),
    .Y(_0751_));
 sky130_fd_sc_hd__inv_2 _1033_ (.A(_0383_),
    .Y(_0752_));
 sky130_fd_sc_hd__inv_2 _1034_ (.A(_0383_),
    .Y(_0753_));
 sky130_fd_sc_hd__inv_2 _1035_ (.A(_0383_),
    .Y(_0754_));
 sky130_fd_sc_hd__inv_2 _1036_ (.A(_0383_),
    .Y(_0755_));
 sky130_fd_sc_hd__inv_2 _1037_ (.A(_0383_),
    .Y(_0756_));
 sky130_fd_sc_hd__inv_2 _1038_ (.A(_0383_),
    .Y(_0757_));
 sky130_fd_sc_hd__inv_2 _1039_ (.A(_0383_),
    .Y(_0758_));
 sky130_fd_sc_hd__inv_2 _1040_ (.A(_0383_),
    .Y(_0759_));
 sky130_fd_sc_hd__buf_8 _1041_ (.A(_0374_),
    .X(_0384_));
 sky130_fd_sc_hd__inv_2 _1042_ (.A(_0384_),
    .Y(_0760_));
 sky130_fd_sc_hd__inv_2 _1043_ (.A(_0384_),
    .Y(_0761_));
 sky130_fd_sc_hd__inv_2 _1044_ (.A(_0384_),
    .Y(_0762_));
 sky130_fd_sc_hd__inv_2 _1045_ (.A(_0384_),
    .Y(_0763_));
 sky130_fd_sc_hd__inv_2 _1046_ (.A(_0384_),
    .Y(_0764_));
 sky130_fd_sc_hd__inv_2 _1047_ (.A(_0384_),
    .Y(_0765_));
 sky130_fd_sc_hd__inv_2 _1048_ (.A(_0384_),
    .Y(_0766_));
 sky130_fd_sc_hd__inv_2 _1049_ (.A(_0384_),
    .Y(_0767_));
 sky130_fd_sc_hd__inv_2 _1050_ (.A(_0384_),
    .Y(_0768_));
 sky130_fd_sc_hd__inv_2 _1051_ (.A(_0384_),
    .Y(_0769_));
 sky130_fd_sc_hd__buf_8 _1052_ (.A(_0374_),
    .X(_0385_));
 sky130_fd_sc_hd__inv_2 _1053_ (.A(_0385_),
    .Y(_0770_));
 sky130_fd_sc_hd__inv_2 _1054_ (.A(_0385_),
    .Y(_0771_));
 sky130_fd_sc_hd__inv_2 _1055_ (.A(_0385_),
    .Y(_0776_));
 sky130_fd_sc_hd__inv_2 _1056_ (.A(_0385_),
    .Y(_0773_));
 sky130_fd_sc_hd__inv_2 _1057_ (.A(_0385_),
    .Y(_0772_));
 sky130_fd_sc_hd__inv_2 _1058_ (.A(_0385_),
    .Y(_0774_));
 sky130_fd_sc_hd__inv_2 _1059_ (.A(_0385_),
    .Y(_0781_));
 sky130_fd_sc_hd__inv_2 _1060_ (.A(_0385_),
    .Y(_0782_));
 sky130_fd_sc_hd__inv_2 _1061_ (.A(_0385_),
    .Y(_0783_));
 sky130_fd_sc_hd__inv_2 _1062_ (.A(_0385_),
    .Y(_0779_));
 sky130_fd_sc_hd__inv_2 _1063_ (.A(_0375_),
    .Y(_0780_));
 sky130_fd_sc_hd__inv_2 _1064_ (.A(_0375_),
    .Y(_0777_));
 sky130_fd_sc_hd__inv_2 _1065_ (.A(_0375_),
    .Y(_0775_));
 sky130_fd_sc_hd__inv_2 _1066_ (.A(_0375_),
    .Y(_0784_));
 sky130_fd_sc_hd__inv_2 _1067_ (.A(_0375_),
    .Y(_0785_));
 sky130_fd_sc_hd__inv_2 _1068_ (.A(_0375_),
    .Y(_0786_));
 sky130_fd_sc_hd__inv_2 _1069_ (.A(_0375_),
    .Y(_0816_));
 sky130_fd_sc_hd__inv_2 _1070_ (.A(_0375_),
    .Y(_0778_));
 sky130_fd_sc_hd__xnor2_1 _1071_ (.A(\gps_channel0.ca_gen.g2[10] ),
    .B(\gps_channel0.ca_gen.g2[9] ),
    .Y(_0386_));
 sky130_fd_sc_hd__xnor2_1 _1072_ (.A(\gps_channel0.ca_gen.g2[3] ),
    .B(\gps_channel0.ca_gen.g2[2] ),
    .Y(_0387_));
 sky130_fd_sc_hd__xor2_1 _1073_ (.A(\gps_channel0.ca_gen.g2[8] ),
    .B(\gps_channel0.ca_gen.g2[6] ),
    .X(_0388_));
 sky130_fd_sc_hd__xnor2_1 _1074_ (.A(_0387_),
    .B(_0388_),
    .Y(_0389_));
 sky130_fd_sc_hd__xnor2_1 _1075_ (.A(_0386_),
    .B(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__clkbuf_4 _1076_ (.A(net22),
    .X(_0391_));
 sky130_fd_sc_hd__mux2_1 _1077_ (.A0(\gps_channel0.ca_gen.g2_init[1] ),
    .A1(_0390_),
    .S(_0391_),
    .X(_0392_));
 sky130_fd_sc_hd__clkbuf_1 _1078_ (.A(_0392_),
    .X(_0000_));
 sky130_fd_sc_hd__mux2_1 _1079_ (.A0(\gps_channel0.ca_gen.g2_init[2] ),
    .A1(\gps_channel0.ca_gen.g2[1] ),
    .S(_0391_),
    .X(_0393_));
 sky130_fd_sc_hd__clkbuf_1 _1080_ (.A(_0393_),
    .X(_0001_));
 sky130_fd_sc_hd__mux2_1 _1081_ (.A0(\gps_channel0.ca_gen.g2_init[3] ),
    .A1(\gps_channel0.ca_gen.g2[2] ),
    .S(_0391_),
    .X(_0394_));
 sky130_fd_sc_hd__clkbuf_1 _1082_ (.A(_0394_),
    .X(_0002_));
 sky130_fd_sc_hd__mux2_1 _1083_ (.A0(\gps_channel0.ca_gen.g2_init[4] ),
    .A1(\gps_channel0.ca_gen.g2[3] ),
    .S(_0391_),
    .X(_0395_));
 sky130_fd_sc_hd__clkbuf_1 _1084_ (.A(_0395_),
    .X(_0003_));
 sky130_fd_sc_hd__mux2_1 _1085_ (.A0(\gps_channel0.ca_gen.g2_init[5] ),
    .A1(\gps_channel0.ca_gen.g2[4] ),
    .S(_0391_),
    .X(_0396_));
 sky130_fd_sc_hd__clkbuf_1 _1086_ (.A(_0396_),
    .X(_0004_));
 sky130_fd_sc_hd__mux2_1 _1087_ (.A0(\gps_channel0.ca_gen.g2_init[6] ),
    .A1(\gps_channel0.ca_gen.g2[5] ),
    .S(_0391_),
    .X(_0397_));
 sky130_fd_sc_hd__clkbuf_1 _1088_ (.A(_0397_),
    .X(_0005_));
 sky130_fd_sc_hd__mux2_1 _1089_ (.A0(\gps_channel0.ca_gen.g2_init[7] ),
    .A1(\gps_channel0.ca_gen.g2[6] ),
    .S(_0391_),
    .X(_0398_));
 sky130_fd_sc_hd__clkbuf_1 _1090_ (.A(_0398_),
    .X(_0006_));
 sky130_fd_sc_hd__mux2_1 _1091_ (.A0(\gps_channel0.ca_gen.g2_init[8] ),
    .A1(\gps_channel0.ca_gen.g2[7] ),
    .S(_0391_),
    .X(_0399_));
 sky130_fd_sc_hd__clkbuf_1 _1092_ (.A(_0399_),
    .X(_0007_));
 sky130_fd_sc_hd__mux2_1 _1093_ (.A0(\gps_channel0.ca_gen.g2_init[9] ),
    .A1(\gps_channel0.ca_gen.g2[8] ),
    .S(_0391_),
    .X(_0400_));
 sky130_fd_sc_hd__clkbuf_1 _1094_ (.A(_0400_),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_1 _1095_ (.A0(\gps_channel0.ca_gen.g2_init[10] ),
    .A1(\gps_channel0.ca_gen.g2[9] ),
    .S(_0391_),
    .X(_0401_));
 sky130_fd_sc_hd__clkbuf_1 _1096_ (.A(_0401_),
    .X(_0009_));
 sky130_fd_sc_hd__xnor2_1 _1097_ (.A(\gps_channel0.ca_gen.g1[10] ),
    .B(net2),
    .Y(_0402_));
 sky130_fd_sc_hd__xor2_1 _1098_ (.A(\gps_channel0.ca_gen.g2[10] ),
    .B(\gps_channel0.lo_i ),
    .X(_0403_));
 sky130_fd_sc_hd__xnor2_1 _1099_ (.A(_0402_),
    .B(_0403_),
    .Y(\gps_channel0.prompt_i ));
 sky130_fd_sc_hd__xor2_1 _1100_ (.A(\gps_channel0.lo_nco.accumulator[30] ),
    .B(\gps_channel0.prompt_i ),
    .X(\gps_channel0.prompt_q ));
 sky130_fd_sc_hd__nand2_1 _1101_ (.A(\gps_channel0.lo_nco.step[0] ),
    .B(net8),
    .Y(_0404_));
 sky130_fd_sc_hd__xnor2_1 _1102_ (.A(\gps_channel0.lo_nco.accumulator[0] ),
    .B(_0404_),
    .Y(_0405_));
 sky130_fd_sc_hd__nor2_4 _1103_ (.A(\gps_channel0.lo_nco.phase_sync ),
    .B(net3),
    .Y(_0406_));
 sky130_fd_sc_hd__mux2_1 _1104_ (.A0(\gps_channel0.lo_nco.phase_in[0] ),
    .A1(_0405_),
    .S(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__clkbuf_1 _1105_ (.A(_0407_),
    .X(_0010_));
 sky130_fd_sc_hd__or2_1 _1106_ (.A(\gps_channel0.lo_nco.phase_sync ),
    .B(net3),
    .X(_0408_));
 sky130_fd_sc_hd__clkbuf_4 _1107_ (.A(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__nor2_4 _1108_ (.A(net8),
    .B(_0409_),
    .Y(_0410_));
 sky130_fd_sc_hd__or2_1 _1109_ (.A(\gps_channel0.lo_nco.step[1] ),
    .B(\gps_channel0.lo_nco.accumulator[1] ),
    .X(_0411_));
 sky130_fd_sc_hd__nand2_1 _1110_ (.A(\gps_channel0.lo_nco.step[1] ),
    .B(\gps_channel0.lo_nco.accumulator[1] ),
    .Y(_0412_));
 sky130_fd_sc_hd__nand4_1 _1111_ (.A(\gps_channel0.lo_nco.step[0] ),
    .B(\gps_channel0.lo_nco.accumulator[0] ),
    .C(_0411_),
    .D(_0412_),
    .Y(_0413_));
 sky130_fd_sc_hd__and2_1 _1112_ (.A(net8),
    .B(_0406_),
    .X(_0414_));
 sky130_fd_sc_hd__a22o_1 _1113_ (.A1(\gps_channel0.lo_nco.step[0] ),
    .A2(\gps_channel0.lo_nco.accumulator[0] ),
    .B1(_0411_),
    .B2(_0412_),
    .X(_0415_));
 sky130_fd_sc_hd__and3_1 _1114_ (.A(_0413_),
    .B(_0414_),
    .C(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__a221o_1 _1115_ (.A1(\gps_channel0.lo_nco.phase_in[1] ),
    .A2(_0409_),
    .B1(_0410_),
    .B2(\gps_channel0.lo_nco.accumulator[1] ),
    .C1(_0416_),
    .X(_0011_));
 sky130_fd_sc_hd__clkbuf_4 _1116_ (.A(_0406_),
    .X(_0417_));
 sky130_fd_sc_hd__or2_1 _1117_ (.A(net8),
    .B(_0409_),
    .X(_0418_));
 sky130_fd_sc_hd__clkbuf_4 _1118_ (.A(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__and2_1 _1119_ (.A(\gps_channel0.lo_nco.step[1] ),
    .B(\gps_channel0.lo_nco.accumulator[1] ),
    .X(_0420_));
 sky130_fd_sc_hd__a31o_1 _1120_ (.A1(\gps_channel0.lo_nco.step[0] ),
    .A2(\gps_channel0.lo_nco.accumulator[0] ),
    .A3(_0411_),
    .B1(_0420_),
    .X(_0421_));
 sky130_fd_sc_hd__nor2_1 _1121_ (.A(\gps_channel0.lo_nco.step[2] ),
    .B(\gps_channel0.lo_nco.accumulator[2] ),
    .Y(_0422_));
 sky130_fd_sc_hd__and2_1 _1122_ (.A(\gps_channel0.lo_nco.step[2] ),
    .B(\gps_channel0.lo_nco.accumulator[2] ),
    .X(_0423_));
 sky130_fd_sc_hd__nor2_2 _1123_ (.A(_0422_),
    .B(_0423_),
    .Y(_0424_));
 sky130_fd_sc_hd__nand2_1 _1124_ (.A(_0421_),
    .B(_0424_),
    .Y(_0425_));
 sky130_fd_sc_hd__or2_1 _1125_ (.A(_0421_),
    .B(_0424_),
    .X(_0426_));
 sky130_fd_sc_hd__nand2_1 _1126_ (.A(net8),
    .B(_0406_),
    .Y(_0427_));
 sky130_fd_sc_hd__clkbuf_4 _1127_ (.A(_0427_),
    .X(_0428_));
 sky130_fd_sc_hd__a21o_1 _1128_ (.A1(_0425_),
    .A2(_0426_),
    .B1(_0428_),
    .X(_0429_));
 sky130_fd_sc_hd__o221a_1 _1129_ (.A1(\gps_channel0.lo_nco.phase_in[2] ),
    .A2(_0417_),
    .B1(_0419_),
    .B2(\gps_channel0.lo_nco.accumulator[2] ),
    .C1(_0429_),
    .X(_0012_));
 sky130_fd_sc_hd__or2_1 _1130_ (.A(\gps_channel0.lo_nco.step[3] ),
    .B(\gps_channel0.lo_nco.accumulator[3] ),
    .X(_0430_));
 sky130_fd_sc_hd__nand2_1 _1131_ (.A(\gps_channel0.lo_nco.step[3] ),
    .B(\gps_channel0.lo_nco.accumulator[3] ),
    .Y(_0431_));
 sky130_fd_sc_hd__nand2_1 _1132_ (.A(_0430_),
    .B(_0431_),
    .Y(_0432_));
 sky130_fd_sc_hd__a21o_1 _1133_ (.A1(_0421_),
    .A2(_0424_),
    .B1(_0423_),
    .X(_0433_));
 sky130_fd_sc_hd__xnor2_1 _1134_ (.A(_0432_),
    .B(_0433_),
    .Y(_0434_));
 sky130_fd_sc_hd__mux2_1 _1135_ (.A0(\gps_channel0.lo_nco.phase_in[3] ),
    .A1(_0434_),
    .S(_0406_),
    .X(_0435_));
 sky130_fd_sc_hd__mux2_1 _1136_ (.A0(\gps_channel0.lo_nco.accumulator[3] ),
    .A1(_0435_),
    .S(_0419_),
    .X(_0436_));
 sky130_fd_sc_hd__clkbuf_1 _1137_ (.A(_0436_),
    .X(_0013_));
 sky130_fd_sc_hd__nand2_1 _1138_ (.A(\gps_channel0.lo_nco.step[4] ),
    .B(\gps_channel0.lo_nco.accumulator[4] ),
    .Y(_0437_));
 sky130_fd_sc_hd__or2_1 _1139_ (.A(\gps_channel0.lo_nco.step[4] ),
    .B(\gps_channel0.lo_nco.accumulator[4] ),
    .X(_0438_));
 sky130_fd_sc_hd__nand2_1 _1140_ (.A(_0437_),
    .B(_0438_),
    .Y(_0439_));
 sky130_fd_sc_hd__and2_1 _1141_ (.A(\gps_channel0.lo_nco.step[3] ),
    .B(\gps_channel0.lo_nco.accumulator[3] ),
    .X(_0440_));
 sky130_fd_sc_hd__and3_1 _1142_ (.A(\gps_channel0.lo_nco.step[2] ),
    .B(\gps_channel0.lo_nco.accumulator[2] ),
    .C(_0430_),
    .X(_0441_));
 sky130_fd_sc_hd__a311oi_4 _1143_ (.A1(_0421_),
    .A2(_0424_),
    .A3(_0430_),
    .B1(_0440_),
    .C1(_0441_),
    .Y(_0442_));
 sky130_fd_sc_hd__nand2_1 _1144_ (.A(_0439_),
    .B(_0442_),
    .Y(_0443_));
 sky130_fd_sc_hd__or2_1 _1145_ (.A(_0439_),
    .B(_0442_),
    .X(_0444_));
 sky130_fd_sc_hd__a21o_1 _1146_ (.A1(_0443_),
    .A2(_0444_),
    .B1(_0428_),
    .X(_0445_));
 sky130_fd_sc_hd__o221a_1 _1147_ (.A1(\gps_channel0.lo_nco.phase_in[4] ),
    .A2(_0417_),
    .B1(_0419_),
    .B2(\gps_channel0.lo_nco.accumulator[4] ),
    .C1(_0445_),
    .X(_0014_));
 sky130_fd_sc_hd__o21a_1 _1148_ (.A1(_0439_),
    .A2(_0442_),
    .B1(_0437_),
    .X(_0446_));
 sky130_fd_sc_hd__or2_1 _1149_ (.A(\gps_channel0.lo_nco.step[5] ),
    .B(\gps_channel0.lo_nco.accumulator[5] ),
    .X(_0447_));
 sky130_fd_sc_hd__nand2_1 _1150_ (.A(\gps_channel0.lo_nco.step[5] ),
    .B(\gps_channel0.lo_nco.accumulator[5] ),
    .Y(_0448_));
 sky130_fd_sc_hd__and2_1 _1151_ (.A(_0447_),
    .B(_0448_),
    .X(_0449_));
 sky130_fd_sc_hd__xnor2_1 _1152_ (.A(_0446_),
    .B(_0449_),
    .Y(_0450_));
 sky130_fd_sc_hd__or2_1 _1153_ (.A(\gps_channel0.lo_nco.phase_in[5] ),
    .B(_0406_),
    .X(_0451_));
 sky130_fd_sc_hd__o221a_1 _1154_ (.A1(\gps_channel0.lo_nco.accumulator[5] ),
    .A2(_0419_),
    .B1(_0450_),
    .B2(_0428_),
    .C1(_0451_),
    .X(_0015_));
 sky130_fd_sc_hd__nand2_1 _1155_ (.A(_0446_),
    .B(_0448_),
    .Y(_0452_));
 sky130_fd_sc_hd__xor2_1 _1156_ (.A(\gps_channel0.lo_nco.step[6] ),
    .B(\gps_channel0.lo_nco.accumulator[6] ),
    .X(_0453_));
 sky130_fd_sc_hd__a21oi_1 _1157_ (.A1(_0447_),
    .A2(_0452_),
    .B1(_0453_),
    .Y(_0454_));
 sky130_fd_sc_hd__a31o_1 _1158_ (.A1(_0447_),
    .A2(_0452_),
    .A3(_0453_),
    .B1(_0427_),
    .X(_0455_));
 sky130_fd_sc_hd__a22oi_1 _1159_ (.A1(\gps_channel0.lo_nco.phase_in[6] ),
    .A2(_0409_),
    .B1(_0410_),
    .B2(\gps_channel0.lo_nco.accumulator[6] ),
    .Y(_0456_));
 sky130_fd_sc_hd__o21ai_1 _1160_ (.A1(_0454_),
    .A2(_0455_),
    .B1(_0456_),
    .Y(_0016_));
 sky130_fd_sc_hd__clkbuf_4 _1161_ (.A(_0410_),
    .X(_0457_));
 sky130_fd_sc_hd__or2_1 _1162_ (.A(\gps_channel0.lo_nco.step[7] ),
    .B(\gps_channel0.lo_nco.accumulator[7] ),
    .X(_0458_));
 sky130_fd_sc_hd__nand2_1 _1163_ (.A(\gps_channel0.lo_nco.step[7] ),
    .B(\gps_channel0.lo_nco.accumulator[7] ),
    .Y(_0459_));
 sky130_fd_sc_hd__a32o_1 _1164_ (.A1(_0447_),
    .A2(_0452_),
    .A3(_0453_),
    .B1(\gps_channel0.lo_nco.accumulator[6] ),
    .B2(\gps_channel0.lo_nco.step[6] ),
    .X(_0460_));
 sky130_fd_sc_hd__a21oi_1 _1165_ (.A1(_0458_),
    .A2(_0459_),
    .B1(_0460_),
    .Y(_0461_));
 sky130_fd_sc_hd__and3_1 _1166_ (.A(_0458_),
    .B(_0459_),
    .C(_0460_),
    .X(_0462_));
 sky130_fd_sc_hd__o21ai_1 _1167_ (.A1(_0461_),
    .A2(_0462_),
    .B1(_0417_),
    .Y(_0463_));
 sky130_fd_sc_hd__o21a_1 _1168_ (.A1(\gps_channel0.lo_nco.phase_in[7] ),
    .A2(_0417_),
    .B1(_0419_),
    .X(_0464_));
 sky130_fd_sc_hd__a22o_1 _1169_ (.A1(\gps_channel0.lo_nco.accumulator[7] ),
    .A2(_0457_),
    .B1(_0463_),
    .B2(_0464_),
    .X(_0017_));
 sky130_fd_sc_hd__and3_1 _1170_ (.A(_0453_),
    .B(_0458_),
    .C(_0459_),
    .X(_0465_));
 sky130_fd_sc_hd__or4bb_1 _1171_ (.A(_0439_),
    .B(_0442_),
    .C_N(_0449_),
    .D_N(_0465_),
    .X(_0466_));
 sky130_fd_sc_hd__nand2_1 _1172_ (.A(_0437_),
    .B(_0448_),
    .Y(_0467_));
 sky130_fd_sc_hd__nand3_1 _1173_ (.A(_0447_),
    .B(_0467_),
    .C(_0465_),
    .Y(_0468_));
 sky130_fd_sc_hd__and3_1 _1174_ (.A(\gps_channel0.lo_nco.step[6] ),
    .B(\gps_channel0.lo_nco.accumulator[6] ),
    .C(_0458_),
    .X(_0469_));
 sky130_fd_sc_hd__a21oi_1 _1175_ (.A1(\gps_channel0.lo_nco.step[7] ),
    .A2(\gps_channel0.lo_nco.accumulator[7] ),
    .B1(_0469_),
    .Y(_0470_));
 sky130_fd_sc_hd__and3_1 _1176_ (.A(_0466_),
    .B(_0468_),
    .C(_0470_),
    .X(_0471_));
 sky130_fd_sc_hd__nand2_1 _1177_ (.A(\gps_channel0.lo_nco.step[8] ),
    .B(\gps_channel0.lo_nco.accumulator[8] ),
    .Y(_0472_));
 sky130_fd_sc_hd__or2_1 _1178_ (.A(\gps_channel0.lo_nco.step[8] ),
    .B(\gps_channel0.lo_nco.accumulator[8] ),
    .X(_0473_));
 sky130_fd_sc_hd__nand2_1 _1179_ (.A(_0472_),
    .B(_0473_),
    .Y(_0474_));
 sky130_fd_sc_hd__nand2_1 _1180_ (.A(_0471_),
    .B(_0474_),
    .Y(_0475_));
 sky130_fd_sc_hd__or2_1 _1181_ (.A(_0471_),
    .B(_0474_),
    .X(_0476_));
 sky130_fd_sc_hd__a21o_1 _1182_ (.A1(_0475_),
    .A2(_0476_),
    .B1(_0428_),
    .X(_0477_));
 sky130_fd_sc_hd__o221a_1 _1183_ (.A1(\gps_channel0.lo_nco.phase_in[8] ),
    .A2(_0417_),
    .B1(_0419_),
    .B2(\gps_channel0.lo_nco.accumulator[8] ),
    .C1(_0477_),
    .X(_0018_));
 sky130_fd_sc_hd__o21ai_1 _1184_ (.A1(_0471_),
    .A2(_0474_),
    .B1(_0472_),
    .Y(_0478_));
 sky130_fd_sc_hd__nor2_1 _1185_ (.A(\gps_channel0.lo_nco.step[9] ),
    .B(\gps_channel0.lo_nco.accumulator[9] ),
    .Y(_0479_));
 sky130_fd_sc_hd__nand2_1 _1186_ (.A(\gps_channel0.lo_nco.step[9] ),
    .B(\gps_channel0.lo_nco.accumulator[9] ),
    .Y(_0480_));
 sky130_fd_sc_hd__or2b_1 _1187_ (.A(_0479_),
    .B_N(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__a21oi_1 _1188_ (.A1(_0478_),
    .A2(_0481_),
    .B1(_0428_),
    .Y(_0482_));
 sky130_fd_sc_hd__o21ai_1 _1189_ (.A1(_0478_),
    .A2(_0481_),
    .B1(_0482_),
    .Y(_0483_));
 sky130_fd_sc_hd__o221a_1 _1190_ (.A1(\gps_channel0.lo_nco.phase_in[9] ),
    .A2(_0417_),
    .B1(_0419_),
    .B2(\gps_channel0.lo_nco.accumulator[9] ),
    .C1(_0483_),
    .X(_0019_));
 sky130_fd_sc_hd__or2_1 _1191_ (.A(\gps_channel0.lo_nco.step[10] ),
    .B(\gps_channel0.lo_nco.accumulator[10] ),
    .X(_0484_));
 sky130_fd_sc_hd__nand2_1 _1192_ (.A(\gps_channel0.lo_nco.step[10] ),
    .B(\gps_channel0.lo_nco.accumulator[10] ),
    .Y(_0485_));
 sky130_fd_sc_hd__nand2_1 _1193_ (.A(_0484_),
    .B(_0485_),
    .Y(_0486_));
 sky130_fd_sc_hd__a21o_1 _1194_ (.A1(_0472_),
    .A2(_0480_),
    .B1(_0479_),
    .X(_0487_));
 sky130_fd_sc_hd__o31a_1 _1195_ (.A1(_0471_),
    .A2(_0474_),
    .A3(_0479_),
    .B1(_0487_),
    .X(_0488_));
 sky130_fd_sc_hd__xnor2_1 _1196_ (.A(_0486_),
    .B(_0488_),
    .Y(_0489_));
 sky130_fd_sc_hd__nor2_1 _1197_ (.A(_0428_),
    .B(_0489_),
    .Y(_0490_));
 sky130_fd_sc_hd__a221o_1 _1198_ (.A1(\gps_channel0.lo_nco.phase_in[10] ),
    .A2(_0409_),
    .B1(_0410_),
    .B2(\gps_channel0.lo_nco.accumulator[10] ),
    .C1(_0490_),
    .X(_0020_));
 sky130_fd_sc_hd__nor2_1 _1199_ (.A(\gps_channel0.lo_nco.step[11] ),
    .B(\gps_channel0.lo_nco.accumulator[11] ),
    .Y(_0491_));
 sky130_fd_sc_hd__and2_1 _1200_ (.A(\gps_channel0.lo_nco.step[11] ),
    .B(\gps_channel0.lo_nco.accumulator[11] ),
    .X(_0492_));
 sky130_fd_sc_hd__nor2_1 _1201_ (.A(_0491_),
    .B(_0492_),
    .Y(_0493_));
 sky130_fd_sc_hd__o21a_1 _1202_ (.A1(_0486_),
    .A2(_0488_),
    .B1(_0485_),
    .X(_0494_));
 sky130_fd_sc_hd__xnor2_1 _1203_ (.A(_0493_),
    .B(_0494_),
    .Y(_0495_));
 sky130_fd_sc_hd__mux2_1 _1204_ (.A0(\gps_channel0.lo_nco.phase_in[11] ),
    .A1(_0495_),
    .S(_0406_),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_1 _1205_ (.A0(\gps_channel0.lo_nco.accumulator[11] ),
    .A1(_0496_),
    .S(_0418_),
    .X(_0497_));
 sky130_fd_sc_hd__clkbuf_1 _1206_ (.A(_0497_),
    .X(_0021_));
 sky130_fd_sc_hd__or3_1 _1207_ (.A(_0486_),
    .B(_0491_),
    .C(_0492_),
    .X(_0498_));
 sky130_fd_sc_hd__or3_1 _1208_ (.A(_0474_),
    .B(_0481_),
    .C(_0498_),
    .X(_0499_));
 sky130_fd_sc_hd__a31o_1 _1209_ (.A1(_0466_),
    .A2(_0468_),
    .A3(_0470_),
    .B1(_0499_),
    .X(_0500_));
 sky130_fd_sc_hd__nand2_1 _1210_ (.A(\gps_channel0.lo_nco.step[11] ),
    .B(\gps_channel0.lo_nco.accumulator[11] ),
    .Y(_0501_));
 sky130_fd_sc_hd__o221a_1 _1211_ (.A1(_0485_),
    .A2(_0491_),
    .B1(_0498_),
    .B2(_0487_),
    .C1(_0501_),
    .X(_0502_));
 sky130_fd_sc_hd__nand2_1 _1212_ (.A(\gps_channel0.lo_nco.step[12] ),
    .B(\gps_channel0.lo_nco.accumulator[12] ),
    .Y(_0503_));
 sky130_fd_sc_hd__or2_1 _1213_ (.A(\gps_channel0.lo_nco.step[12] ),
    .B(\gps_channel0.lo_nco.accumulator[12] ),
    .X(_0504_));
 sky130_fd_sc_hd__nand2_1 _1214_ (.A(_0503_),
    .B(_0504_),
    .Y(_0505_));
 sky130_fd_sc_hd__nand3_1 _1215_ (.A(_0500_),
    .B(_0502_),
    .C(_0505_),
    .Y(_0506_));
 sky130_fd_sc_hd__a21o_1 _1216_ (.A1(_0500_),
    .A2(_0502_),
    .B1(_0505_),
    .X(_0507_));
 sky130_fd_sc_hd__a21o_1 _1217_ (.A1(_0506_),
    .A2(_0507_),
    .B1(_0428_),
    .X(_0508_));
 sky130_fd_sc_hd__o221a_1 _1218_ (.A1(\gps_channel0.lo_nco.phase_in[12] ),
    .A2(_0417_),
    .B1(_0419_),
    .B2(\gps_channel0.lo_nco.accumulator[12] ),
    .C1(_0508_),
    .X(_0022_));
 sky130_fd_sc_hd__nand2_1 _1219_ (.A(_0503_),
    .B(_0507_),
    .Y(_0509_));
 sky130_fd_sc_hd__nor2_1 _1220_ (.A(\gps_channel0.lo_nco.step[13] ),
    .B(\gps_channel0.lo_nco.accumulator[13] ),
    .Y(_0510_));
 sky130_fd_sc_hd__nand2_1 _1221_ (.A(\gps_channel0.lo_nco.step[13] ),
    .B(\gps_channel0.lo_nco.accumulator[13] ),
    .Y(_0511_));
 sky130_fd_sc_hd__or2b_1 _1222_ (.A(_0510_),
    .B_N(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__xnor2_1 _1223_ (.A(_0509_),
    .B(_0512_),
    .Y(_0513_));
 sky130_fd_sc_hd__or2_1 _1224_ (.A(\gps_channel0.lo_nco.phase_in[13] ),
    .B(_0406_),
    .X(_0514_));
 sky130_fd_sc_hd__o221a_1 _1225_ (.A1(\gps_channel0.lo_nco.accumulator[13] ),
    .A2(_0419_),
    .B1(_0513_),
    .B2(_0428_),
    .C1(_0514_),
    .X(_0023_));
 sky130_fd_sc_hd__clkbuf_4 _1226_ (.A(_0414_),
    .X(_0515_));
 sky130_fd_sc_hd__and3_1 _1227_ (.A(_0503_),
    .B(_0507_),
    .C(_0511_),
    .X(_0516_));
 sky130_fd_sc_hd__or2_1 _1228_ (.A(\gps_channel0.lo_nco.step[14] ),
    .B(\gps_channel0.lo_nco.accumulator[14] ),
    .X(_0517_));
 sky130_fd_sc_hd__nand2_1 _1229_ (.A(\gps_channel0.lo_nco.step[14] ),
    .B(\gps_channel0.lo_nco.accumulator[14] ),
    .Y(_0518_));
 sky130_fd_sc_hd__nand2_1 _1230_ (.A(_0517_),
    .B(_0518_),
    .Y(_0519_));
 sky130_fd_sc_hd__o21ai_1 _1231_ (.A1(_0510_),
    .A2(_0516_),
    .B1(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__or3_1 _1232_ (.A(_0510_),
    .B(_0516_),
    .C(_0519_),
    .X(_0521_));
 sky130_fd_sc_hd__a22o_1 _1233_ (.A1(\gps_channel0.lo_nco.phase_in[14] ),
    .A2(_0409_),
    .B1(_0410_),
    .B2(\gps_channel0.lo_nco.accumulator[14] ),
    .X(_0522_));
 sky130_fd_sc_hd__a31o_1 _1234_ (.A1(_0515_),
    .A2(_0520_),
    .A3(_0521_),
    .B1(_0522_),
    .X(_0024_));
 sky130_fd_sc_hd__nor2_1 _1235_ (.A(\gps_channel0.lo_nco.step[15] ),
    .B(\gps_channel0.lo_nco.accumulator[15] ),
    .Y(_0523_));
 sky130_fd_sc_hd__nand2_1 _1236_ (.A(\gps_channel0.lo_nco.step[15] ),
    .B(\gps_channel0.lo_nco.accumulator[15] ),
    .Y(_0524_));
 sky130_fd_sc_hd__and2b_1 _1237_ (.A_N(_0523_),
    .B(_0524_),
    .X(_0525_));
 sky130_fd_sc_hd__o31a_1 _1238_ (.A1(_0510_),
    .A2(_0516_),
    .A3(_0519_),
    .B1(_0518_),
    .X(_0526_));
 sky130_fd_sc_hd__xor2_1 _1239_ (.A(_0525_),
    .B(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__nand2_1 _1240_ (.A(_0417_),
    .B(_0527_),
    .Y(_0528_));
 sky130_fd_sc_hd__o21a_1 _1241_ (.A1(\gps_channel0.lo_nco.phase_in[15] ),
    .A2(_0417_),
    .B1(_0419_),
    .X(_0529_));
 sky130_fd_sc_hd__a22o_1 _1242_ (.A1(\gps_channel0.lo_nco.accumulator[15] ),
    .A2(_0457_),
    .B1(_0528_),
    .B2(_0529_),
    .X(_0025_));
 sky130_fd_sc_hd__nor2_1 _1243_ (.A(\gps_channel0.ca_nco.step[11] ),
    .B(\gps_channel0.ca_nco.accumulator[11] ),
    .Y(_0530_));
 sky130_fd_sc_hd__nand2_1 _1244_ (.A(\gps_channel0.ca_nco.step[10] ),
    .B(\gps_channel0.ca_nco.accumulator[10] ),
    .Y(_0531_));
 sky130_fd_sc_hd__or2_1 _1245_ (.A(\gps_channel0.ca_nco.step[10] ),
    .B(\gps_channel0.ca_nco.accumulator[10] ),
    .X(_0532_));
 sky130_fd_sc_hd__nand2_1 _1246_ (.A(_0531_),
    .B(_0532_),
    .Y(_0533_));
 sky130_fd_sc_hd__nand2_1 _1247_ (.A(\gps_channel0.ca_nco.step[11] ),
    .B(\gps_channel0.ca_nco.accumulator[11] ),
    .Y(_0534_));
 sky130_fd_sc_hd__or3b_1 _1248_ (.A(_0530_),
    .B(_0533_),
    .C_N(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__nand2_1 _1249_ (.A(\gps_channel0.ca_nco.step[9] ),
    .B(\gps_channel0.ca_nco.accumulator[9] ),
    .Y(_0536_));
 sky130_fd_sc_hd__nand2_1 _1250_ (.A(\gps_channel0.ca_nco.step[8] ),
    .B(\gps_channel0.ca_nco.accumulator[8] ),
    .Y(_0537_));
 sky130_fd_sc_hd__nor2_1 _1251_ (.A(\gps_channel0.ca_nco.step[9] ),
    .B(\gps_channel0.ca_nco.accumulator[9] ),
    .Y(_0538_));
 sky130_fd_sc_hd__a21o_1 _1252_ (.A1(_0536_),
    .A2(_0537_),
    .B1(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__o221a_1 _1253_ (.A1(_0530_),
    .A2(_0531_),
    .B1(_0535_),
    .B2(_0539_),
    .C1(_0534_),
    .X(_0540_));
 sky130_fd_sc_hd__nand2_1 _1254_ (.A(\gps_channel0.ca_nco.step[3] ),
    .B(\gps_channel0.ca_nco.accumulator[3] ),
    .Y(_0541_));
 sky130_fd_sc_hd__nand2_1 _1255_ (.A(\gps_channel0.ca_nco.step[2] ),
    .B(\gps_channel0.ca_nco.accumulator[2] ),
    .Y(_0542_));
 sky130_fd_sc_hd__or2_1 _1256_ (.A(\gps_channel0.ca_nco.step[2] ),
    .B(\gps_channel0.ca_nco.accumulator[2] ),
    .X(_0543_));
 sky130_fd_sc_hd__nand2_1 _1257_ (.A(_0542_),
    .B(_0543_),
    .Y(_0544_));
 sky130_fd_sc_hd__xor2_1 _1258_ (.A(\gps_channel0.ca_nco.step[1] ),
    .B(\gps_channel0.ca_nco.accumulator[1] ),
    .X(_0545_));
 sky130_fd_sc_hd__and2_1 _1259_ (.A(\gps_channel0.ca_nco.step[0] ),
    .B(\gps_channel0.ca_nco.accumulator[0] ),
    .X(_0546_));
 sky130_fd_sc_hd__and2_1 _1260_ (.A(\gps_channel0.ca_nco.step[1] ),
    .B(\gps_channel0.ca_nco.accumulator[1] ),
    .X(_0547_));
 sky130_fd_sc_hd__a21oi_1 _1261_ (.A1(_0545_),
    .A2(_0546_),
    .B1(_0547_),
    .Y(_0548_));
 sky130_fd_sc_hd__o21a_1 _1262_ (.A1(_0544_),
    .A2(_0548_),
    .B1(_0542_),
    .X(_0549_));
 sky130_fd_sc_hd__nand2_1 _1263_ (.A(\gps_channel0.ca_nco.step[4] ),
    .B(\gps_channel0.ca_nco.accumulator[4] ),
    .Y(_0550_));
 sky130_fd_sc_hd__or2_1 _1264_ (.A(\gps_channel0.ca_nco.step[4] ),
    .B(\gps_channel0.ca_nco.accumulator[4] ),
    .X(_0551_));
 sky130_fd_sc_hd__nand2_1 _1265_ (.A(_0550_),
    .B(_0551_),
    .Y(_0552_));
 sky130_fd_sc_hd__nor2_1 _1266_ (.A(\gps_channel0.ca_nco.step[3] ),
    .B(\gps_channel0.ca_nco.accumulator[3] ),
    .Y(_0553_));
 sky130_fd_sc_hd__nor2_1 _1267_ (.A(\gps_channel0.ca_nco.step[5] ),
    .B(\gps_channel0.ca_nco.accumulator[5] ),
    .Y(_0554_));
 sky130_fd_sc_hd__nand2_1 _1268_ (.A(\gps_channel0.ca_nco.step[5] ),
    .B(\gps_channel0.ca_nco.accumulator[5] ),
    .Y(_0555_));
 sky130_fd_sc_hd__or2b_1 _1269_ (.A(_0554_),
    .B_N(_0555_),
    .X(_0556_));
 sky130_fd_sc_hd__a2111o_1 _1270_ (.A1(_0541_),
    .A2(_0549_),
    .B1(_0552_),
    .C1(_0553_),
    .D1(_0556_),
    .X(_0557_));
 sky130_fd_sc_hd__nor2_1 _1271_ (.A(\gps_channel0.ca_nco.step[7] ),
    .B(\gps_channel0.ca_nco.accumulator[7] ),
    .Y(_0558_));
 sky130_fd_sc_hd__nand2_1 _1272_ (.A(\gps_channel0.ca_nco.step[6] ),
    .B(\gps_channel0.ca_nco.accumulator[6] ),
    .Y(_0559_));
 sky130_fd_sc_hd__a21o_1 _1273_ (.A1(_0555_),
    .A2(_0550_),
    .B1(_0554_),
    .X(_0560_));
 sky130_fd_sc_hd__nand2_1 _1274_ (.A(\gps_channel0.ca_nco.step[7] ),
    .B(\gps_channel0.ca_nco.accumulator[7] ),
    .Y(_0561_));
 sky130_fd_sc_hd__o211a_1 _1275_ (.A1(_0558_),
    .A2(_0559_),
    .B1(_0560_),
    .C1(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__inv_2 _1276_ (.A(\gps_channel0.ca_nco.step[6] ),
    .Y(_0563_));
 sky130_fd_sc_hd__inv_2 _1277_ (.A(\gps_channel0.ca_nco.accumulator[6] ),
    .Y(_0564_));
 sky130_fd_sc_hd__a31o_1 _1278_ (.A1(_0563_),
    .A2(_0564_),
    .A3(_0561_),
    .B1(_0558_),
    .X(_0565_));
 sky130_fd_sc_hd__or2_1 _1279_ (.A(\gps_channel0.ca_nco.step[8] ),
    .B(\gps_channel0.ca_nco.accumulator[8] ),
    .X(_0566_));
 sky130_fd_sc_hd__nand2_1 _1280_ (.A(_0537_),
    .B(_0566_),
    .Y(_0567_));
 sky130_fd_sc_hd__or3b_1 _1281_ (.A(_0538_),
    .B(_0567_),
    .C_N(_0536_),
    .X(_0568_));
 sky130_fd_sc_hd__a2111o_1 _1282_ (.A1(_0557_),
    .A2(_0562_),
    .B1(_0565_),
    .C1(_0535_),
    .D1(_0568_),
    .X(_0569_));
 sky130_fd_sc_hd__nand2_1 _1283_ (.A(\gps_channel0.ca_nco.step[12] ),
    .B(\gps_channel0.ca_nco.accumulator[12] ),
    .Y(_0570_));
 sky130_fd_sc_hd__or2_1 _1284_ (.A(\gps_channel0.ca_nco.step[12] ),
    .B(\gps_channel0.ca_nco.accumulator[12] ),
    .X(_0571_));
 sky130_fd_sc_hd__nand2_1 _1285_ (.A(_0570_),
    .B(_0571_),
    .Y(_0572_));
 sky130_fd_sc_hd__a21o_1 _1286_ (.A1(_0540_),
    .A2(_0569_),
    .B1(_0572_),
    .X(_0573_));
 sky130_fd_sc_hd__and2_1 _1287_ (.A(\gps_channel0.ca_nco.step[15] ),
    .B(\gps_channel0.ca_nco.accumulator[15] ),
    .X(_0574_));
 sky130_fd_sc_hd__nor2_1 _1288_ (.A(\gps_channel0.ca_nco.step[15] ),
    .B(\gps_channel0.ca_nco.accumulator[15] ),
    .Y(_0575_));
 sky130_fd_sc_hd__nand2_1 _1289_ (.A(\gps_channel0.ca_nco.step[14] ),
    .B(\gps_channel0.ca_nco.accumulator[14] ),
    .Y(_0576_));
 sky130_fd_sc_hd__or2_1 _1290_ (.A(\gps_channel0.ca_nco.step[14] ),
    .B(\gps_channel0.ca_nco.accumulator[14] ),
    .X(_0577_));
 sky130_fd_sc_hd__nand2_1 _1291_ (.A(_0576_),
    .B(_0577_),
    .Y(_0578_));
 sky130_fd_sc_hd__or3_1 _1292_ (.A(_0574_),
    .B(_0575_),
    .C(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__nor2_1 _1293_ (.A(\gps_channel0.ca_nco.step[13] ),
    .B(\gps_channel0.ca_nco.accumulator[13] ),
    .Y(_0580_));
 sky130_fd_sc_hd__nand2_1 _1294_ (.A(\gps_channel0.ca_nco.step[13] ),
    .B(\gps_channel0.ca_nco.accumulator[13] ),
    .Y(_0581_));
 sky130_fd_sc_hd__and2b_1 _1295_ (.A_N(_0580_),
    .B(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__or2b_1 _1296_ (.A(_0579_),
    .B_N(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__a211o_1 _1297_ (.A1(_0570_),
    .A2(_0581_),
    .B1(_0580_),
    .C1(_0579_),
    .X(_0584_));
 sky130_fd_sc_hd__o21ba_1 _1298_ (.A1(_0575_),
    .A2(_0576_),
    .B1_N(_0574_),
    .X(_0585_));
 sky130_fd_sc_hd__o211ai_4 _1299_ (.A1(_0573_),
    .A2(_0583_),
    .B1(_0584_),
    .C1(_0585_),
    .Y(_0586_));
 sky130_fd_sc_hd__clkbuf_4 _1300_ (.A(\gps_channel0.ca_nco.step[16] ),
    .X(_0587_));
 sky130_fd_sc_hd__nor2_1 _1301_ (.A(_0587_),
    .B(\gps_channel0.ca_nco.accumulator[16] ),
    .Y(_0588_));
 sky130_fd_sc_hd__and2_1 _1302_ (.A(_0587_),
    .B(\gps_channel0.ca_nco.accumulator[16] ),
    .X(_0589_));
 sky130_fd_sc_hd__nor2_1 _1303_ (.A(_0588_),
    .B(_0589_),
    .Y(_0590_));
 sky130_fd_sc_hd__and2_1 _1304_ (.A(_0586_),
    .B(_0590_),
    .X(_0591_));
 sky130_fd_sc_hd__or2_1 _1305_ (.A(\gps_channel0.ca_nco.phase_sync ),
    .B(net3),
    .X(_0592_));
 sky130_fd_sc_hd__buf_2 _1306_ (.A(_0592_),
    .X(_0593_));
 sky130_fd_sc_hd__nor2_2 _1307_ (.A(net19),
    .B(_0593_),
    .Y(_0594_));
 sky130_fd_sc_hd__nor2_1 _1308_ (.A(_0593_),
    .B(_0594_),
    .Y(_0595_));
 sky130_fd_sc_hd__clkbuf_4 _1309_ (.A(_0595_),
    .X(_0596_));
 sky130_fd_sc_hd__clkbuf_4 _1310_ (.A(_0596_),
    .X(_0597_));
 sky130_fd_sc_hd__o21ai_1 _1311_ (.A1(_0586_),
    .A2(_0590_),
    .B1(_0597_),
    .Y(_0598_));
 sky130_fd_sc_hd__clkbuf_4 _1312_ (.A(_0594_),
    .X(_0599_));
 sky130_fd_sc_hd__a2bb2o_1 _1313_ (.A1_N(_0591_),
    .A2_N(_0598_),
    .B1(\gps_channel0.ca_nco.accumulator[16] ),
    .B2(_0599_),
    .X(_0026_));
 sky130_fd_sc_hd__xor2_1 _1314_ (.A(_0587_),
    .B(\gps_channel0.ca_nco.accumulator[17] ),
    .X(_0600_));
 sky130_fd_sc_hd__or3_1 _1315_ (.A(_0589_),
    .B(_0591_),
    .C(_0600_),
    .X(_0601_));
 sky130_fd_sc_hd__o21ai_1 _1316_ (.A1(_0589_),
    .A2(_0591_),
    .B1(_0600_),
    .Y(_0602_));
 sky130_fd_sc_hd__a32o_1 _1317_ (.A1(_0597_),
    .A2(_0601_),
    .A3(_0602_),
    .B1(_0599_),
    .B2(\gps_channel0.ca_nco.accumulator[17] ),
    .X(_0027_));
 sky130_fd_sc_hd__nand2_1 _1318_ (.A(_0591_),
    .B(_0600_),
    .Y(_0603_));
 sky130_fd_sc_hd__clkbuf_4 _1319_ (.A(_0587_),
    .X(_0604_));
 sky130_fd_sc_hd__o21ai_1 _1320_ (.A1(\gps_channel0.ca_nco.accumulator[16] ),
    .A2(\gps_channel0.ca_nco.accumulator[17] ),
    .B1(_0604_),
    .Y(_0605_));
 sky130_fd_sc_hd__nand2_1 _1321_ (.A(_0587_),
    .B(\gps_channel0.ca_nco.accumulator[18] ),
    .Y(_0606_));
 sky130_fd_sc_hd__or2_1 _1322_ (.A(_0587_),
    .B(\gps_channel0.ca_nco.accumulator[18] ),
    .X(_0607_));
 sky130_fd_sc_hd__and2_1 _1323_ (.A(_0606_),
    .B(_0607_),
    .X(_0608_));
 sky130_fd_sc_hd__a21bo_1 _1324_ (.A1(_0603_),
    .A2(_0605_),
    .B1_N(_0608_),
    .X(_0609_));
 sky130_fd_sc_hd__nand3b_1 _1325_ (.A_N(_0608_),
    .B(_0603_),
    .C(_0605_),
    .Y(_0610_));
 sky130_fd_sc_hd__buf_4 _1326_ (.A(_0594_),
    .X(_0611_));
 sky130_fd_sc_hd__a32o_1 _1327_ (.A1(_0597_),
    .A2(_0609_),
    .A3(_0610_),
    .B1(_0611_),
    .B2(\gps_channel0.ca_nco.accumulator[18] ),
    .X(_0028_));
 sky130_fd_sc_hd__xnor2_1 _1328_ (.A(_0587_),
    .B(\gps_channel0.ca_nco.accumulator[19] ),
    .Y(_0612_));
 sky130_fd_sc_hd__a21oi_1 _1329_ (.A1(_0606_),
    .A2(_0609_),
    .B1(_0612_),
    .Y(_0613_));
 sky130_fd_sc_hd__clkinv_2 _1330_ (.A(_0595_),
    .Y(_0614_));
 sky130_fd_sc_hd__a31o_1 _1331_ (.A1(_0606_),
    .A2(_0609_),
    .A3(_0612_),
    .B1(_0614_),
    .X(_0615_));
 sky130_fd_sc_hd__a2bb2o_1 _1332_ (.A1_N(_0613_),
    .A2_N(_0615_),
    .B1(\gps_channel0.ca_nco.accumulator[19] ),
    .B2(_0599_),
    .X(_0029_));
 sky130_fd_sc_hd__or2_1 _1333_ (.A(\gps_channel0.ca_nco.step[16] ),
    .B(\gps_channel0.ca_nco.accumulator[20] ),
    .X(_0616_));
 sky130_fd_sc_hd__nand2_1 _1334_ (.A(\gps_channel0.ca_nco.step[16] ),
    .B(\gps_channel0.ca_nco.accumulator[20] ),
    .Y(_0617_));
 sky130_fd_sc_hd__nand2_1 _1335_ (.A(_0616_),
    .B(_0617_),
    .Y(_0618_));
 sky130_fd_sc_hd__clkinv_2 _1336_ (.A(_0612_),
    .Y(_0619_));
 sky130_fd_sc_hd__and4_1 _1337_ (.A(_0590_),
    .B(_0600_),
    .C(_0608_),
    .D(_0619_),
    .X(_0620_));
 sky130_fd_sc_hd__o41a_1 _1338_ (.A1(\gps_channel0.ca_nco.accumulator[16] ),
    .A2(\gps_channel0.ca_nco.accumulator[17] ),
    .A3(\gps_channel0.ca_nco.accumulator[18] ),
    .A4(\gps_channel0.ca_nco.accumulator[19] ),
    .B1(_0587_),
    .X(_0621_));
 sky130_fd_sc_hd__a21oi_1 _1339_ (.A1(_0586_),
    .A2(_0620_),
    .B1(_0621_),
    .Y(_0622_));
 sky130_fd_sc_hd__or2_1 _1340_ (.A(_0618_),
    .B(_0622_),
    .X(_0623_));
 sky130_fd_sc_hd__nand2_1 _1341_ (.A(_0618_),
    .B(_0622_),
    .Y(_0624_));
 sky130_fd_sc_hd__a32o_1 _1342_ (.A1(_0597_),
    .A2(_0623_),
    .A3(_0624_),
    .B1(_0611_),
    .B2(\gps_channel0.ca_nco.accumulator[20] ),
    .X(_0030_));
 sky130_fd_sc_hd__xnor2_1 _1343_ (.A(\gps_channel0.ca_nco.step[16] ),
    .B(\gps_channel0.ca_nco.accumulator[21] ),
    .Y(_0625_));
 sky130_fd_sc_hd__o21a_1 _1344_ (.A1(_0618_),
    .A2(_0622_),
    .B1(_0617_),
    .X(_0626_));
 sky130_fd_sc_hd__xor2_1 _1345_ (.A(_0625_),
    .B(_0626_),
    .X(_0627_));
 sky130_fd_sc_hd__a22o_1 _1346_ (.A1(\gps_channel0.ca_nco.accumulator[21] ),
    .A2(_0599_),
    .B1(_0597_),
    .B2(_0627_),
    .X(_0031_));
 sky130_fd_sc_hd__or3_1 _1347_ (.A(_0618_),
    .B(_0622_),
    .C(_0625_),
    .X(_0628_));
 sky130_fd_sc_hd__o21ai_1 _1348_ (.A1(\gps_channel0.ca_nco.accumulator[20] ),
    .A2(\gps_channel0.ca_nco.accumulator[21] ),
    .B1(_0604_),
    .Y(_0629_));
 sky130_fd_sc_hd__nand2_1 _1349_ (.A(\gps_channel0.ca_nco.step[16] ),
    .B(\gps_channel0.ca_nco.accumulator[22] ),
    .Y(_0630_));
 sky130_fd_sc_hd__or2_1 _1350_ (.A(\gps_channel0.ca_nco.step[16] ),
    .B(\gps_channel0.ca_nco.accumulator[22] ),
    .X(_0631_));
 sky130_fd_sc_hd__nand2_1 _1351_ (.A(_0630_),
    .B(_0631_),
    .Y(_0632_));
 sky130_fd_sc_hd__a21o_1 _1352_ (.A1(_0628_),
    .A2(_0629_),
    .B1(_0632_),
    .X(_0633_));
 sky130_fd_sc_hd__a31oi_1 _1353_ (.A1(_0632_),
    .A2(_0628_),
    .A3(_0629_),
    .B1(_0614_),
    .Y(_0634_));
 sky130_fd_sc_hd__a22o_1 _1354_ (.A1(\gps_channel0.ca_nco.accumulator[22] ),
    .A2(_0599_),
    .B1(_0633_),
    .B2(_0634_),
    .X(_0032_));
 sky130_fd_sc_hd__xor2_1 _1355_ (.A(\gps_channel0.ca_nco.step[16] ),
    .B(\gps_channel0.ca_nco.accumulator[23] ),
    .X(_0635_));
 sky130_fd_sc_hd__inv_2 _1356_ (.A(_0635_),
    .Y(_0636_));
 sky130_fd_sc_hd__a21o_1 _1357_ (.A1(_0630_),
    .A2(_0633_),
    .B1(_0636_),
    .X(_0637_));
 sky130_fd_sc_hd__nand3_1 _1358_ (.A(_0630_),
    .B(_0633_),
    .C(_0636_),
    .Y(_0638_));
 sky130_fd_sc_hd__a32o_1 _1359_ (.A1(_0597_),
    .A2(_0637_),
    .A3(_0638_),
    .B1(_0611_),
    .B2(\gps_channel0.ca_nco.accumulator[23] ),
    .X(_0033_));
 sky130_fd_sc_hd__inv_2 _1360_ (.A(_0621_),
    .Y(_0639_));
 sky130_fd_sc_hd__or4_1 _1361_ (.A(_0618_),
    .B(_0625_),
    .C(_0632_),
    .D(_0636_),
    .X(_0640_));
 sky130_fd_sc_hd__inv_2 _1362_ (.A(_0640_),
    .Y(_0641_));
 sky130_fd_sc_hd__o41a_1 _1363_ (.A1(\gps_channel0.ca_nco.accumulator[20] ),
    .A2(\gps_channel0.ca_nco.accumulator[21] ),
    .A3(\gps_channel0.ca_nco.accumulator[22] ),
    .A4(\gps_channel0.ca_nco.accumulator[23] ),
    .B1(_0587_),
    .X(_0642_));
 sky130_fd_sc_hd__a31oi_1 _1364_ (.A1(_0586_),
    .A2(_0620_),
    .A3(_0641_),
    .B1(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__and2_1 _1365_ (.A(_0639_),
    .B(_0643_),
    .X(_0644_));
 sky130_fd_sc_hd__xnor2_1 _1366_ (.A(_0604_),
    .B(\gps_channel0.ca_nco.accumulator[24] ),
    .Y(_0645_));
 sky130_fd_sc_hd__nand2_1 _1367_ (.A(_0644_),
    .B(_0645_),
    .Y(_0646_));
 sky130_fd_sc_hd__o21a_1 _1368_ (.A1(_0644_),
    .A2(_0645_),
    .B1(_0597_),
    .X(_0647_));
 sky130_fd_sc_hd__a22o_1 _1369_ (.A1(\gps_channel0.ca_nco.accumulator[24] ),
    .A2(_0599_),
    .B1(_0646_),
    .B2(_0647_),
    .X(_0034_));
 sky130_fd_sc_hd__xor2_1 _1370_ (.A(_0587_),
    .B(\gps_channel0.ca_nco.accumulator[25] ),
    .X(_0648_));
 sky130_fd_sc_hd__a2bb2o_1 _1371_ (.A1_N(_0644_),
    .A2_N(_0645_),
    .B1(_0604_),
    .B2(\gps_channel0.ca_nco.accumulator[24] ),
    .X(_0649_));
 sky130_fd_sc_hd__nand2_1 _1372_ (.A(_0648_),
    .B(_0649_),
    .Y(_0650_));
 sky130_fd_sc_hd__o21a_1 _1373_ (.A1(_0648_),
    .A2(_0649_),
    .B1(_0596_),
    .X(_0651_));
 sky130_fd_sc_hd__a22o_1 _1374_ (.A1(\gps_channel0.ca_nco.accumulator[25] ),
    .A2(_0599_),
    .B1(_0650_),
    .B2(_0651_),
    .X(_0035_));
 sky130_fd_sc_hd__inv_2 _1375_ (.A(_0648_),
    .Y(_0652_));
 sky130_fd_sc_hd__a211o_1 _1376_ (.A1(_0639_),
    .A2(_0643_),
    .B1(_0645_),
    .C1(_0652_),
    .X(_0653_));
 sky130_fd_sc_hd__o21ai_2 _1377_ (.A1(\gps_channel0.ca_nco.accumulator[24] ),
    .A2(\gps_channel0.ca_nco.accumulator[25] ),
    .B1(_0604_),
    .Y(_0654_));
 sky130_fd_sc_hd__or2_1 _1378_ (.A(_0604_),
    .B(\gps_channel0.ca_nco.accumulator[26] ),
    .X(_0655_));
 sky130_fd_sc_hd__nand2_1 _1379_ (.A(_0604_),
    .B(\gps_channel0.ca_nco.accumulator[26] ),
    .Y(_0656_));
 sky130_fd_sc_hd__nand2_1 _1380_ (.A(_0655_),
    .B(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__a21o_1 _1381_ (.A1(_0653_),
    .A2(_0654_),
    .B1(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__nand3_1 _1382_ (.A(_0657_),
    .B(_0653_),
    .C(_0654_),
    .Y(_0659_));
 sky130_fd_sc_hd__a32o_1 _1383_ (.A1(_0597_),
    .A2(_0658_),
    .A3(_0659_),
    .B1(_0611_),
    .B2(\gps_channel0.ca_nco.accumulator[26] ),
    .X(_0036_));
 sky130_fd_sc_hd__xnor2_1 _1384_ (.A(_0604_),
    .B(\gps_channel0.ca_nco.accumulator[27] ),
    .Y(_0660_));
 sky130_fd_sc_hd__nand3_1 _1385_ (.A(_0656_),
    .B(_0658_),
    .C(_0660_),
    .Y(_0661_));
 sky130_fd_sc_hd__a21o_1 _1386_ (.A1(_0656_),
    .A2(_0658_),
    .B1(_0660_),
    .X(_0662_));
 sky130_fd_sc_hd__a32o_1 _1387_ (.A1(_0597_),
    .A2(_0661_),
    .A3(_0662_),
    .B1(_0611_),
    .B2(\gps_channel0.ca_nco.accumulator[27] ),
    .X(_0037_));
 sky130_fd_sc_hd__or2_1 _1388_ (.A(_0657_),
    .B(_0660_),
    .X(_0663_));
 sky130_fd_sc_hd__o21ai_1 _1389_ (.A1(\gps_channel0.ca_nco.accumulator[26] ),
    .A2(\gps_channel0.ca_nco.accumulator[27] ),
    .B1(_0604_),
    .Y(_0664_));
 sky130_fd_sc_hd__o211ai_4 _1390_ (.A1(_0653_),
    .A2(_0663_),
    .B1(_0664_),
    .C1(_0654_),
    .Y(_0665_));
 sky130_fd_sc_hd__clkbuf_4 _1391_ (.A(_0593_),
    .X(_0666_));
 sky130_fd_sc_hd__a31oi_1 _1392_ (.A1(net19),
    .A2(\gps_channel0.ca_nco.accumulator[28] ),
    .A3(_0665_),
    .B1(_0666_),
    .Y(_0667_));
 sky130_fd_sc_hd__a21o_1 _1393_ (.A1(_0596_),
    .A2(_0665_),
    .B1(\gps_channel0.ca_nco.accumulator[28] ),
    .X(_0668_));
 sky130_fd_sc_hd__and2_1 _1394_ (.A(_0667_),
    .B(_0668_),
    .X(_0669_));
 sky130_fd_sc_hd__clkbuf_1 _1395_ (.A(_0669_),
    .X(_0038_));
 sky130_fd_sc_hd__and3_1 _1396_ (.A(\gps_channel0.ca_nco.accumulator[28] ),
    .B(_0596_),
    .C(_0665_),
    .X(_0670_));
 sky130_fd_sc_hd__mux2_1 _1397_ (.A0(_0670_),
    .A1(_0667_),
    .S(\gps_channel0.ca_nco.accumulator[29] ),
    .X(_0671_));
 sky130_fd_sc_hd__clkbuf_1 _1398_ (.A(_0671_),
    .X(_0039_));
 sky130_fd_sc_hd__and2_1 _1399_ (.A(\gps_channel0.ca_nco.accumulator[28] ),
    .B(\gps_channel0.ca_nco.accumulator[29] ),
    .X(_0672_));
 sky130_fd_sc_hd__a21oi_1 _1400_ (.A1(_0665_),
    .A2(_0672_),
    .B1(\gps_channel0.ca_nco.accumulator[30] ),
    .Y(_0673_));
 sky130_fd_sc_hd__a31o_1 _1401_ (.A1(\gps_channel0.ca_nco.accumulator[30] ),
    .A2(_0665_),
    .A3(_0672_),
    .B1(_0614_),
    .X(_0674_));
 sky130_fd_sc_hd__a2bb2o_1 _1402_ (.A1_N(_0673_),
    .A2_N(_0674_),
    .B1(\gps_channel0.ca_nco.accumulator[30] ),
    .B2(_0599_),
    .X(_0040_));
 sky130_fd_sc_hd__or2_1 _1403_ (.A(net19),
    .B(_0593_),
    .X(_0675_));
 sky130_fd_sc_hd__buf_4 _1404_ (.A(_0675_),
    .X(_0676_));
 sky130_fd_sc_hd__and2_1 _1405_ (.A(net28),
    .B(_0676_),
    .X(_0677_));
 sky130_fd_sc_hd__and4_1 _1406_ (.A(\gps_channel0.ca_nco.accumulator[30] ),
    .B(_0596_),
    .C(_0665_),
    .D(_0672_),
    .X(_0678_));
 sky130_fd_sc_hd__o2bb2a_1 _1407_ (.A1_N(_0674_),
    .A2_N(_0677_),
    .B1(_0678_),
    .B2(net28),
    .X(_0041_));
 sky130_fd_sc_hd__nor2_1 _1408_ (.A(\gps_channel0.ca_nco.step[0] ),
    .B(\gps_channel0.ca_nco.accumulator[0] ),
    .Y(_0679_));
 sky130_fd_sc_hd__nor2_1 _1409_ (.A(_0546_),
    .B(_0679_),
    .Y(_0680_));
 sky130_fd_sc_hd__a22o_1 _1410_ (.A1(\gps_channel0.ca_nco.phase_in[0] ),
    .A2(_0666_),
    .B1(_0594_),
    .B2(\gps_channel0.ca_nco.accumulator[0] ),
    .X(_0681_));
 sky130_fd_sc_hd__a21o_1 _1411_ (.A1(_0597_),
    .A2(_0680_),
    .B1(_0681_),
    .X(_0042_));
 sky130_fd_sc_hd__a21oi_1 _1412_ (.A1(_0545_),
    .A2(_0546_),
    .B1(_0614_),
    .Y(_0682_));
 sky130_fd_sc_hd__o21a_1 _1413_ (.A1(_0545_),
    .A2(_0546_),
    .B1(_0682_),
    .X(_0683_));
 sky130_fd_sc_hd__a221o_1 _1414_ (.A1(\gps_channel0.ca_nco.phase_in[1] ),
    .A2(_0666_),
    .B1(_0611_),
    .B2(\gps_channel0.ca_nco.accumulator[1] ),
    .C1(_0683_),
    .X(_0043_));
 sky130_fd_sc_hd__xor2_1 _1415_ (.A(_0544_),
    .B(_0548_),
    .X(_0684_));
 sky130_fd_sc_hd__nor2_4 _1416_ (.A(\gps_channel0.ca_nco.phase_sync ),
    .B(net3),
    .Y(_0685_));
 sky130_fd_sc_hd__mux2_1 _1417_ (.A0(\gps_channel0.ca_nco.phase_in[2] ),
    .A1(_0684_),
    .S(_0685_),
    .X(_0686_));
 sky130_fd_sc_hd__mux2_1 _1418_ (.A0(\gps_channel0.ca_nco.accumulator[2] ),
    .A1(_0686_),
    .S(_0676_),
    .X(_0687_));
 sky130_fd_sc_hd__clkbuf_1 _1419_ (.A(_0687_),
    .X(_0044_));
 sky130_fd_sc_hd__and2_1 _1420_ (.A(\gps_channel0.ca_nco.step[3] ),
    .B(\gps_channel0.ca_nco.accumulator[3] ),
    .X(_0688_));
 sky130_fd_sc_hd__o21ai_1 _1421_ (.A1(_0553_),
    .A2(_0688_),
    .B1(_0549_),
    .Y(_0689_));
 sky130_fd_sc_hd__o311a_1 _1422_ (.A1(_0553_),
    .A2(_0688_),
    .A3(_0549_),
    .B1(_0596_),
    .C1(_0689_),
    .X(_0690_));
 sky130_fd_sc_hd__a221o_1 _1423_ (.A1(\gps_channel0.ca_nco.phase_in[3] ),
    .A2(_0666_),
    .B1(_0611_),
    .B2(\gps_channel0.ca_nco.accumulator[3] ),
    .C1(_0690_),
    .X(_0045_));
 sky130_fd_sc_hd__a21oi_1 _1424_ (.A1(_0541_),
    .A2(_0549_),
    .B1(_0553_),
    .Y(_0691_));
 sky130_fd_sc_hd__xnor2_1 _1425_ (.A(_0691_),
    .B(_0552_),
    .Y(_0692_));
 sky130_fd_sc_hd__mux2_1 _1426_ (.A0(\gps_channel0.ca_nco.phase_in[4] ),
    .A1(_0692_),
    .S(_0685_),
    .X(_0693_));
 sky130_fd_sc_hd__mux2_1 _1427_ (.A0(\gps_channel0.ca_nco.accumulator[4] ),
    .A1(_0693_),
    .S(_0676_),
    .X(_0694_));
 sky130_fd_sc_hd__clkbuf_1 _1428_ (.A(_0694_),
    .X(_0046_));
 sky130_fd_sc_hd__a21bo_1 _1429_ (.A1(_0691_),
    .A2(_0551_),
    .B1_N(_0550_),
    .X(_0695_));
 sky130_fd_sc_hd__xnor2_1 _1430_ (.A(_0556_),
    .B(_0695_),
    .Y(_0696_));
 sky130_fd_sc_hd__mux2_1 _1431_ (.A0(\gps_channel0.ca_nco.phase_in[5] ),
    .A1(_0696_),
    .S(_0685_),
    .X(_0697_));
 sky130_fd_sc_hd__mux2_1 _1432_ (.A0(\gps_channel0.ca_nco.accumulator[5] ),
    .A1(_0697_),
    .S(_0676_),
    .X(_0698_));
 sky130_fd_sc_hd__clkbuf_1 _1433_ (.A(_0698_),
    .X(_0047_));
 sky130_fd_sc_hd__or2_1 _1434_ (.A(\gps_channel0.ca_nco.step[6] ),
    .B(\gps_channel0.ca_nco.accumulator[6] ),
    .X(_0699_));
 sky130_fd_sc_hd__nand2_1 _1435_ (.A(_0559_),
    .B(_0699_),
    .Y(_0700_));
 sky130_fd_sc_hd__and3_1 _1436_ (.A(_0557_),
    .B(_0560_),
    .C(_0700_),
    .X(_0701_));
 sky130_fd_sc_hd__a21o_1 _1437_ (.A1(_0557_),
    .A2(_0560_),
    .B1(_0700_),
    .X(_0702_));
 sky130_fd_sc_hd__and3b_1 _1438_ (.A_N(_0701_),
    .B(_0702_),
    .C(_0596_),
    .X(_0703_));
 sky130_fd_sc_hd__a221o_1 _1439_ (.A1(\gps_channel0.ca_nco.phase_in[6] ),
    .A2(_0666_),
    .B1(_0611_),
    .B2(\gps_channel0.ca_nco.accumulator[6] ),
    .C1(_0703_),
    .X(_0048_));
 sky130_fd_sc_hd__clkinv_2 _1440_ (.A(_0558_),
    .Y(_0704_));
 sky130_fd_sc_hd__and2_1 _1441_ (.A(_0561_),
    .B(_0704_),
    .X(_0705_));
 sky130_fd_sc_hd__a21oi_1 _1442_ (.A1(_0559_),
    .A2(_0702_),
    .B1(_0705_),
    .Y(_0706_));
 sky130_fd_sc_hd__a31o_1 _1443_ (.A1(_0559_),
    .A2(_0705_),
    .A3(_0702_),
    .B1(_0593_),
    .X(_0707_));
 sky130_fd_sc_hd__o22a_1 _1444_ (.A1(\gps_channel0.ca_nco.phase_in[7] ),
    .A2(_0685_),
    .B1(_0706_),
    .B2(_0707_),
    .X(_0708_));
 sky130_fd_sc_hd__mux2_1 _1445_ (.A0(\gps_channel0.ca_nco.accumulator[7] ),
    .A1(_0708_),
    .S(_0676_),
    .X(_0709_));
 sky130_fd_sc_hd__clkbuf_1 _1446_ (.A(_0709_),
    .X(_0049_));
 sky130_fd_sc_hd__a21o_1 _1447_ (.A1(_0557_),
    .A2(_0562_),
    .B1(_0565_),
    .X(_0710_));
 sky130_fd_sc_hd__nor2_1 _1448_ (.A(_0710_),
    .B(_0567_),
    .Y(_0711_));
 sky130_fd_sc_hd__nand2_1 _1449_ (.A(_0710_),
    .B(_0567_),
    .Y(_0712_));
 sky130_fd_sc_hd__and3b_1 _1450_ (.A_N(_0711_),
    .B(_0596_),
    .C(_0712_),
    .X(_0713_));
 sky130_fd_sc_hd__a221o_1 _1451_ (.A1(\gps_channel0.ca_nco.phase_in[8] ),
    .A2(_0666_),
    .B1(_0611_),
    .B2(\gps_channel0.ca_nco.accumulator[8] ),
    .C1(_0713_),
    .X(_0050_));
 sky130_fd_sc_hd__and2b_1 _1452_ (.A_N(_0538_),
    .B(_0536_),
    .X(_0714_));
 sky130_fd_sc_hd__o21ai_1 _1453_ (.A1(_0710_),
    .A2(_0567_),
    .B1(_0537_),
    .Y(_0715_));
 sky130_fd_sc_hd__xor2_1 _1454_ (.A(_0714_),
    .B(_0715_),
    .X(_0716_));
 sky130_fd_sc_hd__mux2_1 _1455_ (.A0(\gps_channel0.ca_nco.phase_in[9] ),
    .A1(_0716_),
    .S(_0685_),
    .X(_0717_));
 sky130_fd_sc_hd__mux2_1 _1456_ (.A0(\gps_channel0.ca_nco.accumulator[9] ),
    .A1(_0717_),
    .S(_0676_),
    .X(_0718_));
 sky130_fd_sc_hd__clkbuf_1 _1457_ (.A(_0718_),
    .X(_0051_));
 sky130_fd_sc_hd__nand2_1 _1458_ (.A(_0714_),
    .B(_0711_),
    .Y(_0719_));
 sky130_fd_sc_hd__and3_1 _1459_ (.A(_0719_),
    .B(_0539_),
    .C(_0533_),
    .X(_0720_));
 sky130_fd_sc_hd__a21o_1 _1460_ (.A1(_0719_),
    .A2(_0539_),
    .B1(_0533_),
    .X(_0721_));
 sky130_fd_sc_hd__and3b_1 _1461_ (.A_N(_0720_),
    .B(_0721_),
    .C(_0596_),
    .X(_0722_));
 sky130_fd_sc_hd__a221o_1 _1462_ (.A1(\gps_channel0.ca_nco.phase_in[10] ),
    .A2(_0666_),
    .B1(_0611_),
    .B2(\gps_channel0.ca_nco.accumulator[10] ),
    .C1(_0722_),
    .X(_0052_));
 sky130_fd_sc_hd__and2b_1 _1463_ (.A_N(_0530_),
    .B(_0534_),
    .X(_0723_));
 sky130_fd_sc_hd__a21oi_1 _1464_ (.A1(_0531_),
    .A2(_0721_),
    .B1(_0723_),
    .Y(_0724_));
 sky130_fd_sc_hd__a31o_1 _1465_ (.A1(_0531_),
    .A2(_0723_),
    .A3(_0721_),
    .B1(_0593_),
    .X(_0725_));
 sky130_fd_sc_hd__o22a_1 _1466_ (.A1(\gps_channel0.ca_nco.phase_in[11] ),
    .A2(_0685_),
    .B1(_0724_),
    .B2(_0725_),
    .X(_0726_));
 sky130_fd_sc_hd__mux2_1 _1467_ (.A0(\gps_channel0.ca_nco.accumulator[11] ),
    .A1(_0726_),
    .S(_0676_),
    .X(_0727_));
 sky130_fd_sc_hd__clkbuf_1 _1468_ (.A(_0727_),
    .X(_0053_));
 sky130_fd_sc_hd__and3_1 _1469_ (.A(_0540_),
    .B(_0569_),
    .C(_0572_),
    .X(_0728_));
 sky130_fd_sc_hd__or3b_1 _1470_ (.A(_0614_),
    .B(_0728_),
    .C_N(_0573_),
    .X(_0729_));
 sky130_fd_sc_hd__a22oi_1 _1471_ (.A1(\gps_channel0.ca_nco.phase_in[12] ),
    .A2(_0666_),
    .B1(_0594_),
    .B2(\gps_channel0.ca_nco.accumulator[12] ),
    .Y(_0730_));
 sky130_fd_sc_hd__nand2_1 _1472_ (.A(_0729_),
    .B(_0730_),
    .Y(_0054_));
 sky130_fd_sc_hd__and3_1 _1473_ (.A(_0570_),
    .B(_0573_),
    .C(_0582_),
    .X(_0731_));
 sky130_fd_sc_hd__a21oi_1 _1474_ (.A1(_0570_),
    .A2(_0573_),
    .B1(_0582_),
    .Y(_0732_));
 sky130_fd_sc_hd__or3_1 _1475_ (.A(_0666_),
    .B(_0731_),
    .C(_0732_),
    .X(_0733_));
 sky130_fd_sc_hd__a21o_1 _1476_ (.A1(\gps_channel0.ca_nco.phase_in[13] ),
    .A2(_0666_),
    .B1(_0596_),
    .X(_0734_));
 sky130_fd_sc_hd__a22o_1 _1477_ (.A1(\gps_channel0.ca_nco.accumulator[13] ),
    .A2(_0599_),
    .B1(_0733_),
    .B2(_0734_),
    .X(_0055_));
 sky130_fd_sc_hd__a31o_1 _1478_ (.A1(_0570_),
    .A2(_0573_),
    .A3(_0581_),
    .B1(_0580_),
    .X(_0735_));
 sky130_fd_sc_hd__or2_1 _1479_ (.A(_0578_),
    .B(_0735_),
    .X(_0736_));
 sky130_fd_sc_hd__nand2_1 _1480_ (.A(_0578_),
    .B(_0735_),
    .Y(_0737_));
 sky130_fd_sc_hd__and2_1 _1481_ (.A(\gps_channel0.ca_nco.phase_in[14] ),
    .B(_0593_),
    .X(_0738_));
 sky130_fd_sc_hd__a31o_1 _1482_ (.A1(_0685_),
    .A2(_0736_),
    .A3(_0737_),
    .B1(_0738_),
    .X(_0739_));
 sky130_fd_sc_hd__mux2_1 _1483_ (.A0(\gps_channel0.ca_nco.accumulator[14] ),
    .A1(_0739_),
    .S(_0676_),
    .X(_0740_));
 sky130_fd_sc_hd__clkbuf_1 _1484_ (.A(_0740_),
    .X(_0056_));
 sky130_fd_sc_hd__nor2_1 _1485_ (.A(_0574_),
    .B(_0575_),
    .Y(_0741_));
 sky130_fd_sc_hd__a21oi_1 _1486_ (.A1(_0576_),
    .A2(_0736_),
    .B1(_0741_),
    .Y(_0742_));
 sky130_fd_sc_hd__a31o_1 _1487_ (.A1(_0741_),
    .A2(_0576_),
    .A3(_0736_),
    .B1(_0593_),
    .X(_0743_));
 sky130_fd_sc_hd__or2_1 _1488_ (.A(_0742_),
    .B(_0743_),
    .X(_0744_));
 sky130_fd_sc_hd__o21a_1 _1489_ (.A1(\gps_channel0.ca_nco.phase_in[15] ),
    .A2(_0685_),
    .B1(_0676_),
    .X(_0745_));
 sky130_fd_sc_hd__a22o_1 _1490_ (.A1(\gps_channel0.ca_nco.accumulator[15] ),
    .A2(_0599_),
    .B1(_0744_),
    .B2(_0745_),
    .X(_0057_));
 sky130_fd_sc_hd__clkinv_2 _1491_ (.A(net24),
    .Y(_0162_));
 sky130_fd_sc_hd__or2_1 _1492_ (.A(net25),
    .B(net23),
    .X(_0163_));
 sky130_fd_sc_hd__or2_1 _1493_ (.A(_0162_),
    .B(_0163_),
    .X(_0164_));
 sky130_fd_sc_hd__clkbuf_2 _1494_ (.A(_0164_),
    .X(_0165_));
 sky130_fd_sc_hd__clkbuf_4 _1495_ (.A(_0165_),
    .X(_0166_));
 sky130_fd_sc_hd__nor2_4 _1496_ (.A(_0162_),
    .B(_0163_),
    .Y(_0167_));
 sky130_fd_sc_hd__clkbuf_4 _1497_ (.A(_0167_),
    .X(_0168_));
 sky130_fd_sc_hd__buf_2 _1498_ (.A(net3),
    .X(_0169_));
 sky130_fd_sc_hd__o21ba_1 _1499_ (.A1(\gps_channel0.lo_nco.phase_in[0] ),
    .A2(_0168_),
    .B1_N(_0169_),
    .X(_0170_));
 sky130_fd_sc_hd__o21a_1 _1500_ (.A1(net4),
    .A2(_0166_),
    .B1(_0170_),
    .X(_0058_));
 sky130_fd_sc_hd__o21ba_1 _1501_ (.A1(\gps_channel0.lo_nco.phase_in[1] ),
    .A2(_0168_),
    .B1_N(_0169_),
    .X(_0171_));
 sky130_fd_sc_hd__o21a_1 _1502_ (.A1(net5),
    .A2(_0166_),
    .B1(_0171_),
    .X(_0059_));
 sky130_fd_sc_hd__o21ba_1 _1503_ (.A1(\gps_channel0.lo_nco.phase_in[2] ),
    .A2(_0168_),
    .B1_N(_0169_),
    .X(_0172_));
 sky130_fd_sc_hd__o21a_1 _1504_ (.A1(net6),
    .A2(_0166_),
    .B1(_0172_),
    .X(_0060_));
 sky130_fd_sc_hd__o21ba_1 _1505_ (.A1(\gps_channel0.lo_nco.phase_in[3] ),
    .A2(_0168_),
    .B1_N(_0169_),
    .X(_0173_));
 sky130_fd_sc_hd__o21a_1 _1506_ (.A1(net7),
    .A2(_0166_),
    .B1(_0173_),
    .X(_0061_));
 sky130_fd_sc_hd__buf_2 _1507_ (.A(net3),
    .X(_0174_));
 sky130_fd_sc_hd__buf_2 _1508_ (.A(_0174_),
    .X(_0175_));
 sky130_fd_sc_hd__o21ba_1 _1509_ (.A1(\gps_channel0.lo_nco.phase_in[4] ),
    .A2(_0168_),
    .B1_N(_0175_),
    .X(_0176_));
 sky130_fd_sc_hd__o21a_1 _1510_ (.A1(net9),
    .A2(_0166_),
    .B1(_0176_),
    .X(_0062_));
 sky130_fd_sc_hd__o21ba_1 _1511_ (.A1(\gps_channel0.lo_nco.phase_in[5] ),
    .A2(_0168_),
    .B1_N(_0175_),
    .X(_0177_));
 sky130_fd_sc_hd__o21a_1 _1512_ (.A1(net10),
    .A2(_0166_),
    .B1(_0177_),
    .X(_0063_));
 sky130_fd_sc_hd__o21ba_1 _1513_ (.A1(\gps_channel0.lo_nco.phase_in[6] ),
    .A2(_0168_),
    .B1_N(_0175_),
    .X(_0178_));
 sky130_fd_sc_hd__o21a_1 _1514_ (.A1(net11),
    .A2(_0166_),
    .B1(_0178_),
    .X(_0064_));
 sky130_fd_sc_hd__o21ba_1 _1515_ (.A1(\gps_channel0.lo_nco.phase_in[7] ),
    .A2(_0168_),
    .B1_N(_0175_),
    .X(_0179_));
 sky130_fd_sc_hd__o21a_1 _1516_ (.A1(net12),
    .A2(_0166_),
    .B1(_0179_),
    .X(_0065_));
 sky130_fd_sc_hd__o21ba_1 _1517_ (.A1(\gps_channel0.lo_nco.phase_in[8] ),
    .A2(_0168_),
    .B1_N(_0175_),
    .X(_0180_));
 sky130_fd_sc_hd__o21a_1 _1518_ (.A1(net13),
    .A2(_0166_),
    .B1(_0180_),
    .X(_0066_));
 sky130_fd_sc_hd__o21ba_1 _1519_ (.A1(\gps_channel0.lo_nco.phase_in[9] ),
    .A2(_0167_),
    .B1_N(_0175_),
    .X(_0181_));
 sky130_fd_sc_hd__o21a_1 _1520_ (.A1(net14),
    .A2(_0166_),
    .B1(_0181_),
    .X(_0067_));
 sky130_fd_sc_hd__o21ba_1 _1521_ (.A1(\gps_channel0.lo_nco.phase_in[10] ),
    .A2(_0167_),
    .B1_N(_0175_),
    .X(_0182_));
 sky130_fd_sc_hd__o21a_1 _1522_ (.A1(net15),
    .A2(_0165_),
    .B1(_0182_),
    .X(_0068_));
 sky130_fd_sc_hd__o21ba_1 _1523_ (.A1(\gps_channel0.lo_nco.phase_in[11] ),
    .A2(_0167_),
    .B1_N(_0175_),
    .X(_0183_));
 sky130_fd_sc_hd__o21a_1 _1524_ (.A1(net16),
    .A2(_0165_),
    .B1(_0183_),
    .X(_0069_));
 sky130_fd_sc_hd__o21ba_1 _1525_ (.A1(\gps_channel0.lo_nco.phase_in[12] ),
    .A2(_0167_),
    .B1_N(_0175_),
    .X(_0184_));
 sky130_fd_sc_hd__o21a_1 _1526_ (.A1(net17),
    .A2(_0165_),
    .B1(_0184_),
    .X(_0070_));
 sky130_fd_sc_hd__o21ba_1 _1527_ (.A1(\gps_channel0.lo_nco.phase_in[13] ),
    .A2(_0167_),
    .B1_N(_0175_),
    .X(_0185_));
 sky130_fd_sc_hd__o21a_1 _1528_ (.A1(net18),
    .A2(_0165_),
    .B1(_0185_),
    .X(_0071_));
 sky130_fd_sc_hd__buf_2 _1529_ (.A(net3),
    .X(_0186_));
 sky130_fd_sc_hd__o21ba_1 _1530_ (.A1(\gps_channel0.lo_nco.phase_in[14] ),
    .A2(_0167_),
    .B1_N(_0186_),
    .X(_0187_));
 sky130_fd_sc_hd__o21a_1 _1531_ (.A1(net20),
    .A2(_0165_),
    .B1(_0187_),
    .X(_0072_));
 sky130_fd_sc_hd__o21ba_1 _1532_ (.A1(\gps_channel0.lo_nco.phase_in[15] ),
    .A2(_0167_),
    .B1_N(_0186_),
    .X(_0188_));
 sky130_fd_sc_hd__o21a_1 _1533_ (.A1(net21),
    .A2(_0165_),
    .B1(_0188_),
    .X(_0073_));
 sky130_fd_sc_hd__inv_2 _1534_ (.A(\gps_channel0.ca_gen.g1[10] ),
    .Y(_0189_));
 sky130_fd_sc_hd__clkbuf_2 _1535_ (.A(net22),
    .X(_0190_));
 sky130_fd_sc_hd__o21ai_1 _1536_ (.A1(\gps_channel0.ca_gen.g1[3] ),
    .A2(_0189_),
    .B1(_0190_),
    .Y(_0191_));
 sky130_fd_sc_hd__a21o_1 _1537_ (.A1(\gps_channel0.ca_gen.g1[3] ),
    .A2(_0189_),
    .B1(_0191_),
    .X(_0074_));
 sky130_fd_sc_hd__or2b_1 _1538_ (.A(\gps_channel0.ca_gen.g1[1] ),
    .B_N(_0190_),
    .X(_0192_));
 sky130_fd_sc_hd__clkbuf_1 _1539_ (.A(_0192_),
    .X(_0075_));
 sky130_fd_sc_hd__or2b_1 _1540_ (.A(\gps_channel0.ca_gen.g1[2] ),
    .B_N(_0190_),
    .X(_0193_));
 sky130_fd_sc_hd__clkbuf_1 _1541_ (.A(_0193_),
    .X(_0076_));
 sky130_fd_sc_hd__or2b_1 _1542_ (.A(\gps_channel0.ca_gen.g1[3] ),
    .B_N(_0190_),
    .X(_0194_));
 sky130_fd_sc_hd__clkbuf_1 _1543_ (.A(_0194_),
    .X(_0077_));
 sky130_fd_sc_hd__or2b_1 _1544_ (.A(\gps_channel0.ca_gen.g1[4] ),
    .B_N(_0190_),
    .X(_0195_));
 sky130_fd_sc_hd__clkbuf_1 _1545_ (.A(_0195_),
    .X(_0078_));
 sky130_fd_sc_hd__or2b_1 _1546_ (.A(\gps_channel0.ca_gen.g1[5] ),
    .B_N(_0190_),
    .X(_0196_));
 sky130_fd_sc_hd__clkbuf_1 _1547_ (.A(_0196_),
    .X(_0079_));
 sky130_fd_sc_hd__or2b_1 _1548_ (.A(\gps_channel0.ca_gen.g1[6] ),
    .B_N(_0190_),
    .X(_0197_));
 sky130_fd_sc_hd__clkbuf_1 _1549_ (.A(_0197_),
    .X(_0080_));
 sky130_fd_sc_hd__or2b_1 _1550_ (.A(\gps_channel0.ca_gen.g1[7] ),
    .B_N(_0190_),
    .X(_0198_));
 sky130_fd_sc_hd__clkbuf_1 _1551_ (.A(_0198_),
    .X(_0081_));
 sky130_fd_sc_hd__or2b_1 _1552_ (.A(\gps_channel0.ca_gen.g1[8] ),
    .B_N(_0190_),
    .X(_0199_));
 sky130_fd_sc_hd__clkbuf_1 _1553_ (.A(_0199_),
    .X(_0082_));
 sky130_fd_sc_hd__or2b_1 _1554_ (.A(\gps_channel0.ca_gen.g1[9] ),
    .B_N(_0190_),
    .X(_0200_));
 sky130_fd_sc_hd__clkbuf_1 _1555_ (.A(_0200_),
    .X(_0083_));
 sky130_fd_sc_hd__or2b_1 _1556_ (.A(_0519_),
    .B_N(_0525_),
    .X(_0201_));
 sky130_fd_sc_hd__or3_1 _1557_ (.A(_0505_),
    .B(_0512_),
    .C(_0201_),
    .X(_0202_));
 sky130_fd_sc_hd__a21o_1 _1558_ (.A1(_0500_),
    .A2(_0502_),
    .B1(_0202_),
    .X(_0203_));
 sky130_fd_sc_hd__a21o_1 _1559_ (.A1(_0503_),
    .A2(_0511_),
    .B1(_0510_),
    .X(_0204_));
 sky130_fd_sc_hd__o221a_1 _1560_ (.A1(_0518_),
    .A2(_0523_),
    .B1(_0201_),
    .B2(_0204_),
    .C1(_0524_),
    .X(_0205_));
 sky130_fd_sc_hd__and2_1 _1561_ (.A(_0203_),
    .B(_0205_),
    .X(_0206_));
 sky130_fd_sc_hd__clkbuf_4 _1562_ (.A(\gps_channel0.lo_nco.step[16] ),
    .X(_0207_));
 sky130_fd_sc_hd__nand2_1 _1563_ (.A(_0207_),
    .B(\gps_channel0.lo_nco.accumulator[16] ),
    .Y(_0208_));
 sky130_fd_sc_hd__or2_1 _1564_ (.A(\gps_channel0.lo_nco.step[16] ),
    .B(\gps_channel0.lo_nco.accumulator[16] ),
    .X(_0209_));
 sky130_fd_sc_hd__nand2_1 _1565_ (.A(_0208_),
    .B(_0209_),
    .Y(_0210_));
 sky130_fd_sc_hd__xor2_1 _1566_ (.A(_0206_),
    .B(_0210_),
    .X(_0211_));
 sky130_fd_sc_hd__a22o_1 _1567_ (.A1(\gps_channel0.lo_nco.accumulator[16] ),
    .A2(_0457_),
    .B1(_0211_),
    .B2(_0515_),
    .X(_0084_));
 sky130_fd_sc_hd__xor2_1 _1568_ (.A(_0207_),
    .B(\gps_channel0.lo_nco.accumulator[17] ),
    .X(_0212_));
 sky130_fd_sc_hd__o21a_1 _1569_ (.A1(_0206_),
    .A2(_0210_),
    .B1(_0208_),
    .X(_0213_));
 sky130_fd_sc_hd__xnor2_1 _1570_ (.A(_0212_),
    .B(_0213_),
    .Y(_0214_));
 sky130_fd_sc_hd__a22o_1 _1571_ (.A1(\gps_channel0.lo_nco.accumulator[17] ),
    .A2(_0457_),
    .B1(_0214_),
    .B2(_0515_),
    .X(_0085_));
 sky130_fd_sc_hd__nand2_1 _1572_ (.A(_0207_),
    .B(\gps_channel0.lo_nco.accumulator[18] ),
    .Y(_0215_));
 sky130_fd_sc_hd__or2_1 _1573_ (.A(_0207_),
    .B(\gps_channel0.lo_nco.accumulator[18] ),
    .X(_0216_));
 sky130_fd_sc_hd__nand2_1 _1574_ (.A(_0215_),
    .B(_0216_),
    .Y(_0217_));
 sky130_fd_sc_hd__buf_2 _1575_ (.A(_0207_),
    .X(_0218_));
 sky130_fd_sc_hd__o21ai_1 _1576_ (.A1(\gps_channel0.lo_nco.accumulator[16] ),
    .A2(\gps_channel0.lo_nco.accumulator[17] ),
    .B1(_0218_),
    .Y(_0219_));
 sky130_fd_sc_hd__or2b_1 _1577_ (.A(_0210_),
    .B_N(_0212_),
    .X(_0220_));
 sky130_fd_sc_hd__or2_1 _1578_ (.A(_0206_),
    .B(_0220_),
    .X(_0221_));
 sky130_fd_sc_hd__nand3_1 _1579_ (.A(_0217_),
    .B(_0219_),
    .C(_0221_),
    .Y(_0222_));
 sky130_fd_sc_hd__a21o_1 _1580_ (.A1(_0219_),
    .A2(_0221_),
    .B1(_0217_),
    .X(_0223_));
 sky130_fd_sc_hd__a32o_1 _1581_ (.A1(_0515_),
    .A2(_0222_),
    .A3(_0223_),
    .B1(_0457_),
    .B2(\gps_channel0.lo_nco.accumulator[18] ),
    .X(_0086_));
 sky130_fd_sc_hd__xor2_1 _1582_ (.A(_0207_),
    .B(\gps_channel0.lo_nco.accumulator[19] ),
    .X(_0224_));
 sky130_fd_sc_hd__inv_2 _1583_ (.A(_0224_),
    .Y(_0225_));
 sky130_fd_sc_hd__nand3_1 _1584_ (.A(_0215_),
    .B(_0223_),
    .C(_0225_),
    .Y(_0226_));
 sky130_fd_sc_hd__a21o_1 _1585_ (.A1(_0215_),
    .A2(_0223_),
    .B1(_0225_),
    .X(_0227_));
 sky130_fd_sc_hd__a32o_1 _1586_ (.A1(_0515_),
    .A2(_0226_),
    .A3(_0227_),
    .B1(_0457_),
    .B2(\gps_channel0.lo_nco.accumulator[19] ),
    .X(_0087_));
 sky130_fd_sc_hd__o41a_1 _1587_ (.A1(\gps_channel0.lo_nco.accumulator[16] ),
    .A2(\gps_channel0.lo_nco.accumulator[17] ),
    .A3(\gps_channel0.lo_nco.accumulator[18] ),
    .A4(\gps_channel0.lo_nco.accumulator[19] ),
    .B1(_0218_),
    .X(_0228_));
 sky130_fd_sc_hd__a2111oi_4 _1588_ (.A1(_0203_),
    .A2(_0205_),
    .B1(_0217_),
    .C1(_0220_),
    .D1(_0225_),
    .Y(_0229_));
 sky130_fd_sc_hd__nor2_1 _1589_ (.A(_0218_),
    .B(\gps_channel0.lo_nco.accumulator[20] ),
    .Y(_0230_));
 sky130_fd_sc_hd__and2_1 _1590_ (.A(_0207_),
    .B(\gps_channel0.lo_nco.accumulator[20] ),
    .X(_0231_));
 sky130_fd_sc_hd__nor2_1 _1591_ (.A(_0230_),
    .B(_0231_),
    .Y(_0232_));
 sky130_fd_sc_hd__o21a_1 _1592_ (.A1(_0228_),
    .A2(_0229_),
    .B1(_0232_),
    .X(_0233_));
 sky130_fd_sc_hd__nor3_1 _1593_ (.A(_0232_),
    .B(_0228_),
    .C(_0229_),
    .Y(_0234_));
 sky130_fd_sc_hd__nor2_1 _1594_ (.A(_0233_),
    .B(_0234_),
    .Y(_0235_));
 sky130_fd_sc_hd__a22o_1 _1595_ (.A1(\gps_channel0.lo_nco.accumulator[20] ),
    .A2(_0457_),
    .B1(_0235_),
    .B2(_0515_),
    .X(_0088_));
 sky130_fd_sc_hd__xor2_1 _1596_ (.A(_0218_),
    .B(\gps_channel0.lo_nco.accumulator[21] ),
    .X(_0236_));
 sky130_fd_sc_hd__or3_1 _1597_ (.A(_0231_),
    .B(_0233_),
    .C(_0236_),
    .X(_0237_));
 sky130_fd_sc_hd__o21ai_1 _1598_ (.A1(_0231_),
    .A2(_0233_),
    .B1(_0236_),
    .Y(_0238_));
 sky130_fd_sc_hd__a32o_1 _1599_ (.A1(_0515_),
    .A2(_0237_),
    .A3(_0238_),
    .B1(_0410_),
    .B2(\gps_channel0.lo_nco.accumulator[21] ),
    .X(_0089_));
 sky130_fd_sc_hd__o21a_1 _1600_ (.A1(\gps_channel0.lo_nco.accumulator[20] ),
    .A2(\gps_channel0.lo_nco.accumulator[21] ),
    .B1(_0218_),
    .X(_0239_));
 sky130_fd_sc_hd__and2_1 _1601_ (.A(_0233_),
    .B(_0236_),
    .X(_0240_));
 sky130_fd_sc_hd__or2_1 _1602_ (.A(_0207_),
    .B(\gps_channel0.lo_nco.accumulator[22] ),
    .X(_0241_));
 sky130_fd_sc_hd__nand2_1 _1603_ (.A(_0207_),
    .B(\gps_channel0.lo_nco.accumulator[22] ),
    .Y(_0242_));
 sky130_fd_sc_hd__and2_1 _1604_ (.A(_0241_),
    .B(_0242_),
    .X(_0243_));
 sky130_fd_sc_hd__o21ai_1 _1605_ (.A1(_0239_),
    .A2(_0240_),
    .B1(_0243_),
    .Y(_0244_));
 sky130_fd_sc_hd__o31a_1 _1606_ (.A1(_0243_),
    .A2(_0239_),
    .A3(_0240_),
    .B1(_0515_),
    .X(_0245_));
 sky130_fd_sc_hd__a22o_1 _1607_ (.A1(\gps_channel0.lo_nco.accumulator[22] ),
    .A2(_0457_),
    .B1(_0244_),
    .B2(_0245_),
    .X(_0090_));
 sky130_fd_sc_hd__xnor2_1 _1608_ (.A(_0207_),
    .B(\gps_channel0.lo_nco.accumulator[23] ),
    .Y(_0246_));
 sky130_fd_sc_hd__a21oi_1 _1609_ (.A1(_0242_),
    .A2(_0244_),
    .B1(_0246_),
    .Y(_0247_));
 sky130_fd_sc_hd__a31o_1 _1610_ (.A1(_0242_),
    .A2(_0244_),
    .A3(_0246_),
    .B1(_0428_),
    .X(_0248_));
 sky130_fd_sc_hd__a2bb2o_1 _1611_ (.A1_N(_0247_),
    .A2_N(_0248_),
    .B1(\gps_channel0.lo_nco.accumulator[23] ),
    .B2(_0457_),
    .X(_0091_));
 sky130_fd_sc_hd__and3b_1 _1612_ (.A_N(_0246_),
    .B(_0242_),
    .C(_0241_),
    .X(_0249_));
 sky130_fd_sc_hd__and3_1 _1613_ (.A(_0232_),
    .B(_0236_),
    .C(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__o21a_1 _1614_ (.A1(\gps_channel0.lo_nco.accumulator[22] ),
    .A2(\gps_channel0.lo_nco.accumulator[23] ),
    .B1(_0218_),
    .X(_0251_));
 sky130_fd_sc_hd__or3_1 _1615_ (.A(_0228_),
    .B(_0239_),
    .C(_0251_),
    .X(_0252_));
 sky130_fd_sc_hd__a21o_1 _1616_ (.A1(_0229_),
    .A2(_0250_),
    .B1(_0252_),
    .X(_0253_));
 sky130_fd_sc_hd__nand2_1 _1617_ (.A(_0218_),
    .B(\gps_channel0.lo_nco.accumulator[24] ),
    .Y(_0254_));
 sky130_fd_sc_hd__or2_1 _1618_ (.A(_0218_),
    .B(\gps_channel0.lo_nco.accumulator[24] ),
    .X(_0255_));
 sky130_fd_sc_hd__nand3_1 _1619_ (.A(_0253_),
    .B(_0254_),
    .C(_0255_),
    .Y(_0256_));
 sky130_fd_sc_hd__a21o_1 _1620_ (.A1(_0254_),
    .A2(_0255_),
    .B1(_0253_),
    .X(_0257_));
 sky130_fd_sc_hd__a32o_1 _1621_ (.A1(_0515_),
    .A2(_0256_),
    .A3(_0257_),
    .B1(_0410_),
    .B2(\gps_channel0.lo_nco.accumulator[24] ),
    .X(_0092_));
 sky130_fd_sc_hd__a221o_1 _1622_ (.A1(_0218_),
    .A2(\gps_channel0.lo_nco.accumulator[24] ),
    .B1(_0229_),
    .B2(_0250_),
    .C1(_0252_),
    .X(_0258_));
 sky130_fd_sc_hd__and3_1 _1623_ (.A(\gps_channel0.lo_nco.accumulator[25] ),
    .B(_0255_),
    .C(_0258_),
    .X(_0259_));
 sky130_fd_sc_hd__nand2_1 _1624_ (.A(net8),
    .B(_0259_),
    .Y(_0260_));
 sky130_fd_sc_hd__a31o_1 _1625_ (.A1(net8),
    .A2(_0255_),
    .A3(_0258_),
    .B1(\gps_channel0.lo_nco.accumulator[25] ),
    .X(_0261_));
 sky130_fd_sc_hd__and3_1 _1626_ (.A(_0417_),
    .B(_0260_),
    .C(_0261_),
    .X(_0262_));
 sky130_fd_sc_hd__clkbuf_1 _1627_ (.A(_0262_),
    .X(_0093_));
 sky130_fd_sc_hd__a31oi_1 _1628_ (.A1(net8),
    .A2(\gps_channel0.lo_nco.accumulator[26] ),
    .A3(_0259_),
    .B1(_0409_),
    .Y(_0263_));
 sky130_fd_sc_hd__a21o_1 _1629_ (.A1(_0414_),
    .A2(_0259_),
    .B1(\gps_channel0.lo_nco.accumulator[26] ),
    .X(_0264_));
 sky130_fd_sc_hd__and2_1 _1630_ (.A(_0263_),
    .B(_0264_),
    .X(_0265_));
 sky130_fd_sc_hd__clkbuf_1 _1631_ (.A(_0265_),
    .X(_0094_));
 sky130_fd_sc_hd__and3_1 _1632_ (.A(\gps_channel0.lo_nco.accumulator[26] ),
    .B(_0414_),
    .C(_0259_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _1633_ (.A0(_0266_),
    .A1(_0263_),
    .S(\gps_channel0.lo_nco.accumulator[27] ),
    .X(_0267_));
 sky130_fd_sc_hd__clkbuf_1 _1634_ (.A(_0267_),
    .X(_0095_));
 sky130_fd_sc_hd__and3_1 _1635_ (.A(\gps_channel0.lo_nco.accumulator[26] ),
    .B(\gps_channel0.lo_nco.accumulator[27] ),
    .C(_0259_),
    .X(_0268_));
 sky130_fd_sc_hd__a31oi_1 _1636_ (.A1(net8),
    .A2(\gps_channel0.lo_nco.accumulator[28] ),
    .A3(_0268_),
    .B1(_0409_),
    .Y(_0269_));
 sky130_fd_sc_hd__a21o_1 _1637_ (.A1(_0414_),
    .A2(_0268_),
    .B1(\gps_channel0.lo_nco.accumulator[28] ),
    .X(_0270_));
 sky130_fd_sc_hd__and2_1 _1638_ (.A(_0269_),
    .B(_0270_),
    .X(_0271_));
 sky130_fd_sc_hd__clkbuf_1 _1639_ (.A(_0271_),
    .X(_0096_));
 sky130_fd_sc_hd__and3_1 _1640_ (.A(\gps_channel0.lo_nco.accumulator[28] ),
    .B(_0414_),
    .C(_0268_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _1641_ (.A0(_0272_),
    .A1(_0269_),
    .S(\gps_channel0.lo_nco.accumulator[29] ),
    .X(_0273_));
 sky130_fd_sc_hd__clkbuf_1 _1642_ (.A(_0273_),
    .X(_0097_));
 sky130_fd_sc_hd__and2_1 _1643_ (.A(\gps_channel0.lo_nco.accumulator[28] ),
    .B(\gps_channel0.lo_nco.accumulator[29] ),
    .X(_0274_));
 sky130_fd_sc_hd__a21o_1 _1644_ (.A1(_0268_),
    .A2(_0274_),
    .B1(\gps_channel0.lo_nco.accumulator[30] ),
    .X(_0275_));
 sky130_fd_sc_hd__a31oi_1 _1645_ (.A1(\gps_channel0.lo_nco.accumulator[30] ),
    .A2(_0268_),
    .A3(_0274_),
    .B1(_0428_),
    .Y(_0276_));
 sky130_fd_sc_hd__a22o_1 _1646_ (.A1(\gps_channel0.lo_nco.accumulator[30] ),
    .A2(_0457_),
    .B1(_0275_),
    .B2(_0276_),
    .X(_0098_));
 sky130_fd_sc_hd__inv_2 _1647_ (.A(\gps_channel0.lo_i ),
    .Y(_0277_));
 sky130_fd_sc_hd__a41o_1 _1648_ (.A1(\gps_channel0.lo_nco.accumulator[30] ),
    .A2(_0515_),
    .A3(_0268_),
    .A4(_0274_),
    .B1(\gps_channel0.lo_i ),
    .X(_0278_));
 sky130_fd_sc_hd__o31a_1 _1649_ (.A1(_0277_),
    .A2(_0410_),
    .A3(_0276_),
    .B1(_0278_),
    .X(_0099_));
 sky130_fd_sc_hd__and3_1 _1650_ (.A(net25),
    .B(net23),
    .C(_0162_),
    .X(_0279_));
 sky130_fd_sc_hd__clkbuf_4 _1651_ (.A(_0279_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _1652_ (.A0(\gps_channel0.ca_gen.g2_init[1] ),
    .A1(net4),
    .S(_0280_),
    .X(_0281_));
 sky130_fd_sc_hd__or2_1 _1653_ (.A(_0169_),
    .B(_0281_),
    .X(_0282_));
 sky130_fd_sc_hd__clkbuf_1 _1654_ (.A(_0282_),
    .X(_0100_));
 sky130_fd_sc_hd__clkbuf_4 _1655_ (.A(_0174_),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _1656_ (.A0(\gps_channel0.ca_gen.g2_init[2] ),
    .A1(net5),
    .S(_0280_),
    .X(_0284_));
 sky130_fd_sc_hd__and2b_1 _1657_ (.A_N(_0283_),
    .B(_0284_),
    .X(_0285_));
 sky130_fd_sc_hd__clkbuf_1 _1658_ (.A(_0285_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _1659_ (.A0(\gps_channel0.ca_gen.g2_init[3] ),
    .A1(net6),
    .S(_0280_),
    .X(_0286_));
 sky130_fd_sc_hd__and2b_1 _1660_ (.A_N(_0283_),
    .B(_0286_),
    .X(_0287_));
 sky130_fd_sc_hd__clkbuf_1 _1661_ (.A(_0287_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _1662_ (.A0(\gps_channel0.ca_gen.g2_init[4] ),
    .A1(net7),
    .S(_0280_),
    .X(_0288_));
 sky130_fd_sc_hd__and2b_1 _1663_ (.A_N(_0283_),
    .B(_0288_),
    .X(_0289_));
 sky130_fd_sc_hd__clkbuf_1 _1664_ (.A(_0289_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _1665_ (.A0(\gps_channel0.ca_gen.g2_init[5] ),
    .A1(net9),
    .S(_0280_),
    .X(_0290_));
 sky130_fd_sc_hd__and2b_1 _1666_ (.A_N(_0283_),
    .B(_0290_),
    .X(_0291_));
 sky130_fd_sc_hd__clkbuf_1 _1667_ (.A(_0291_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _1668_ (.A0(\gps_channel0.ca_gen.g2_init[6] ),
    .A1(net10),
    .S(_0280_),
    .X(_0292_));
 sky130_fd_sc_hd__or2_1 _1669_ (.A(_0169_),
    .B(_0292_),
    .X(_0293_));
 sky130_fd_sc_hd__clkbuf_1 _1670_ (.A(_0293_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _1671_ (.A0(\gps_channel0.ca_gen.g2_init[7] ),
    .A1(net11),
    .S(_0280_),
    .X(_0294_));
 sky130_fd_sc_hd__or2_1 _1672_ (.A(_0169_),
    .B(_0294_),
    .X(_0295_));
 sky130_fd_sc_hd__clkbuf_1 _1673_ (.A(_0295_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _1674_ (.A0(\gps_channel0.ca_gen.g2_init[8] ),
    .A1(net12),
    .S(_0280_),
    .X(_0296_));
 sky130_fd_sc_hd__and2b_1 _1675_ (.A_N(_0169_),
    .B(_0296_),
    .X(_0297_));
 sky130_fd_sc_hd__clkbuf_1 _1676_ (.A(_0297_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _1677_ (.A0(\gps_channel0.ca_gen.g2_init[9] ),
    .A1(net13),
    .S(_0280_),
    .X(_0298_));
 sky130_fd_sc_hd__or2_1 _1678_ (.A(_0169_),
    .B(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__clkbuf_1 _1679_ (.A(_0299_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _1680_ (.A0(\gps_channel0.ca_gen.g2_init[10] ),
    .A1(net14),
    .S(_0280_),
    .X(_0300_));
 sky130_fd_sc_hd__and2b_1 _1681_ (.A_N(_0169_),
    .B(_0300_),
    .X(_0301_));
 sky130_fd_sc_hd__clkbuf_1 _1682_ (.A(_0301_),
    .X(_0109_));
 sky130_fd_sc_hd__inv_2 _1683_ (.A(net25),
    .Y(_0302_));
 sky130_fd_sc_hd__mux2_1 _1684_ (.A0(_0302_),
    .A1(net23),
    .S(_0162_),
    .X(_0303_));
 sky130_fd_sc_hd__and3b_2 _1685_ (.A_N(net23),
    .B(_0162_),
    .C(net25),
    .X(_0304_));
 sky130_fd_sc_hd__clkbuf_4 _1686_ (.A(_0304_),
    .X(_0305_));
 sky130_fd_sc_hd__a21oi_1 _1687_ (.A1(\gps_channel0.ca_nco.phase_sync ),
    .A2(_0303_),
    .B1(_0305_),
    .Y(_0306_));
 sky130_fd_sc_hd__nor2_1 _1688_ (.A(_0283_),
    .B(_0306_),
    .Y(_0110_));
 sky130_fd_sc_hd__o211a_1 _1689_ (.A1(_0302_),
    .A2(_0162_),
    .B1(_0163_),
    .C1(\gps_channel0.lo_nco.phase_sync ),
    .X(_0307_));
 sky130_fd_sc_hd__o21ba_1 _1690_ (.A1(_0168_),
    .A2(_0307_),
    .B1_N(_0283_),
    .X(_0111_));
 sky130_fd_sc_hd__and3_1 _1691_ (.A(_0302_),
    .B(net23),
    .C(_0162_),
    .X(_0308_));
 sky130_fd_sc_hd__clkbuf_2 _1692_ (.A(_0308_),
    .X(_0309_));
 sky130_fd_sc_hd__clkbuf_4 _1693_ (.A(_0309_),
    .X(_0310_));
 sky130_fd_sc_hd__or3b_1 _1694_ (.A(net25),
    .B(net24),
    .C_N(net23),
    .X(_0311_));
 sky130_fd_sc_hd__buf_2 _1695_ (.A(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__clkbuf_4 _1696_ (.A(_0312_),
    .X(_0313_));
 sky130_fd_sc_hd__o21ba_1 _1697_ (.A1(net4),
    .A2(_0313_),
    .B1_N(_0186_),
    .X(_0314_));
 sky130_fd_sc_hd__o21a_1 _1698_ (.A1(\gps_channel0.lo_nco.step[0] ),
    .A2(_0310_),
    .B1(_0314_),
    .X(_0112_));
 sky130_fd_sc_hd__o21ba_1 _1699_ (.A1(net5),
    .A2(_0313_),
    .B1_N(_0186_),
    .X(_0315_));
 sky130_fd_sc_hd__o21a_1 _1700_ (.A1(\gps_channel0.lo_nco.step[1] ),
    .A2(_0310_),
    .B1(_0315_),
    .X(_0113_));
 sky130_fd_sc_hd__o21ba_1 _1701_ (.A1(net6),
    .A2(_0313_),
    .B1_N(_0186_),
    .X(_0316_));
 sky130_fd_sc_hd__o21a_1 _1702_ (.A1(\gps_channel0.lo_nco.step[2] ),
    .A2(_0310_),
    .B1(_0316_),
    .X(_0114_));
 sky130_fd_sc_hd__o21ba_1 _1703_ (.A1(net7),
    .A2(_0313_),
    .B1_N(_0186_),
    .X(_0317_));
 sky130_fd_sc_hd__o21a_1 _1704_ (.A1(\gps_channel0.lo_nco.step[3] ),
    .A2(_0310_),
    .B1(_0317_),
    .X(_0115_));
 sky130_fd_sc_hd__o21ba_1 _1705_ (.A1(net9),
    .A2(_0313_),
    .B1_N(_0186_),
    .X(_0318_));
 sky130_fd_sc_hd__o21a_1 _1706_ (.A1(\gps_channel0.lo_nco.step[4] ),
    .A2(_0310_),
    .B1(_0318_),
    .X(_0116_));
 sky130_fd_sc_hd__o21ba_1 _1707_ (.A1(net10),
    .A2(_0313_),
    .B1_N(_0186_),
    .X(_0319_));
 sky130_fd_sc_hd__o21a_1 _1708_ (.A1(\gps_channel0.lo_nco.step[5] ),
    .A2(_0310_),
    .B1(_0319_),
    .X(_0117_));
 sky130_fd_sc_hd__o21ba_1 _1709_ (.A1(net11),
    .A2(_0313_),
    .B1_N(_0186_),
    .X(_0320_));
 sky130_fd_sc_hd__o21a_1 _1710_ (.A1(\gps_channel0.lo_nco.step[6] ),
    .A2(_0310_),
    .B1(_0320_),
    .X(_0118_));
 sky130_fd_sc_hd__o21ba_1 _1711_ (.A1(net12),
    .A2(_0313_),
    .B1_N(_0186_),
    .X(_0321_));
 sky130_fd_sc_hd__o21a_1 _1712_ (.A1(\gps_channel0.lo_nco.step[7] ),
    .A2(_0310_),
    .B1(_0321_),
    .X(_0119_));
 sky130_fd_sc_hd__buf_2 _1713_ (.A(net3),
    .X(_0322_));
 sky130_fd_sc_hd__o21ba_1 _1714_ (.A1(net13),
    .A2(_0313_),
    .B1_N(_0322_),
    .X(_0323_));
 sky130_fd_sc_hd__o21a_1 _1715_ (.A1(\gps_channel0.lo_nco.step[8] ),
    .A2(_0310_),
    .B1(_0323_),
    .X(_0120_));
 sky130_fd_sc_hd__o21ba_1 _1716_ (.A1(net14),
    .A2(_0312_),
    .B1_N(_0322_),
    .X(_0324_));
 sky130_fd_sc_hd__o21a_1 _1717_ (.A1(\gps_channel0.lo_nco.step[9] ),
    .A2(_0310_),
    .B1(_0324_),
    .X(_0121_));
 sky130_fd_sc_hd__o21ba_1 _1718_ (.A1(net15),
    .A2(_0312_),
    .B1_N(_0322_),
    .X(_0325_));
 sky130_fd_sc_hd__o21a_1 _1719_ (.A1(\gps_channel0.lo_nco.step[10] ),
    .A2(_0309_),
    .B1(_0325_),
    .X(_0122_));
 sky130_fd_sc_hd__o21ba_1 _1720_ (.A1(net16),
    .A2(_0312_),
    .B1_N(_0322_),
    .X(_0326_));
 sky130_fd_sc_hd__o21a_1 _1721_ (.A1(\gps_channel0.lo_nco.step[11] ),
    .A2(_0309_),
    .B1(_0326_),
    .X(_0123_));
 sky130_fd_sc_hd__o21ba_1 _1722_ (.A1(net17),
    .A2(_0312_),
    .B1_N(_0322_),
    .X(_0327_));
 sky130_fd_sc_hd__o21a_1 _1723_ (.A1(\gps_channel0.lo_nco.step[12] ),
    .A2(_0309_),
    .B1(_0327_),
    .X(_0124_));
 sky130_fd_sc_hd__o21ba_1 _1724_ (.A1(net18),
    .A2(_0312_),
    .B1_N(_0322_),
    .X(_0328_));
 sky130_fd_sc_hd__o21a_1 _1725_ (.A1(\gps_channel0.lo_nco.step[13] ),
    .A2(_0309_),
    .B1(_0328_),
    .X(_0125_));
 sky130_fd_sc_hd__o21ba_1 _1726_ (.A1(net20),
    .A2(_0312_),
    .B1_N(_0322_),
    .X(_0329_));
 sky130_fd_sc_hd__o21a_1 _1727_ (.A1(\gps_channel0.lo_nco.step[14] ),
    .A2(_0309_),
    .B1(_0329_),
    .X(_0126_));
 sky130_fd_sc_hd__o21ba_1 _1728_ (.A1(net21),
    .A2(_0312_),
    .B1_N(_0322_),
    .X(_0330_));
 sky130_fd_sc_hd__o21a_1 _1729_ (.A1(\gps_channel0.lo_nco.step[15] ),
    .A2(_0309_),
    .B1(_0330_),
    .X(_0127_));
 sky130_fd_sc_hd__a21o_1 _1730_ (.A1(_0218_),
    .A2(_0313_),
    .B1(_0283_),
    .X(_0128_));
 sky130_fd_sc_hd__or3b_1 _1731_ (.A(_0162_),
    .B(net25),
    .C_N(net23),
    .X(_0331_));
 sky130_fd_sc_hd__clkbuf_4 _1732_ (.A(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__clkbuf_4 _1733_ (.A(_0332_),
    .X(_0333_));
 sky130_fd_sc_hd__and3_2 _1734_ (.A(_0302_),
    .B(net23),
    .C(net24),
    .X(_0334_));
 sky130_fd_sc_hd__clkbuf_4 _1735_ (.A(_0334_),
    .X(_0335_));
 sky130_fd_sc_hd__o21ba_1 _1736_ (.A1(\gps_channel0.ca_nco.step[0] ),
    .A2(_0335_),
    .B1_N(_0322_),
    .X(_0336_));
 sky130_fd_sc_hd__o21a_1 _1737_ (.A1(net4),
    .A2(_0333_),
    .B1(_0336_),
    .X(_0129_));
 sky130_fd_sc_hd__o21ba_1 _1738_ (.A1(\gps_channel0.ca_nco.step[1] ),
    .A2(_0335_),
    .B1_N(_0322_),
    .X(_0337_));
 sky130_fd_sc_hd__o21a_1 _1739_ (.A1(net5),
    .A2(_0333_),
    .B1(_0337_),
    .X(_0130_));
 sky130_fd_sc_hd__buf_2 _1740_ (.A(net3),
    .X(_0338_));
 sky130_fd_sc_hd__o21ba_1 _1741_ (.A1(\gps_channel0.ca_nco.step[2] ),
    .A2(_0335_),
    .B1_N(_0338_),
    .X(_0339_));
 sky130_fd_sc_hd__o21a_1 _1742_ (.A1(net6),
    .A2(_0333_),
    .B1(_0339_),
    .X(_0131_));
 sky130_fd_sc_hd__o21ba_1 _1743_ (.A1(\gps_channel0.ca_nco.step[3] ),
    .A2(_0335_),
    .B1_N(_0338_),
    .X(_0340_));
 sky130_fd_sc_hd__o21a_1 _1744_ (.A1(net7),
    .A2(_0333_),
    .B1(_0340_),
    .X(_0132_));
 sky130_fd_sc_hd__o21ba_1 _1745_ (.A1(\gps_channel0.ca_nco.step[4] ),
    .A2(_0335_),
    .B1_N(_0338_),
    .X(_0341_));
 sky130_fd_sc_hd__o21a_1 _1746_ (.A1(net9),
    .A2(_0333_),
    .B1(_0341_),
    .X(_0133_));
 sky130_fd_sc_hd__o21ba_1 _1747_ (.A1(\gps_channel0.ca_nco.step[5] ),
    .A2(_0335_),
    .B1_N(_0338_),
    .X(_0342_));
 sky130_fd_sc_hd__o21a_1 _1748_ (.A1(net10),
    .A2(_0333_),
    .B1(_0342_),
    .X(_0134_));
 sky130_fd_sc_hd__a21oi_1 _1749_ (.A1(_0563_),
    .A2(_0332_),
    .B1(_0283_),
    .Y(_0343_));
 sky130_fd_sc_hd__o21a_1 _1750_ (.A1(net11),
    .A2(_0333_),
    .B1(_0343_),
    .X(_0135_));
 sky130_fd_sc_hd__o21ba_1 _1751_ (.A1(\gps_channel0.ca_nco.step[7] ),
    .A2(_0335_),
    .B1_N(_0338_),
    .X(_0344_));
 sky130_fd_sc_hd__o21a_1 _1752_ (.A1(net12),
    .A2(_0333_),
    .B1(_0344_),
    .X(_0136_));
 sky130_fd_sc_hd__o21ba_1 _1753_ (.A1(\gps_channel0.ca_nco.step[8] ),
    .A2(_0335_),
    .B1_N(_0338_),
    .X(_0345_));
 sky130_fd_sc_hd__o21a_1 _1754_ (.A1(net13),
    .A2(_0333_),
    .B1(_0345_),
    .X(_0137_));
 sky130_fd_sc_hd__o21ba_1 _1755_ (.A1(\gps_channel0.ca_nco.step[9] ),
    .A2(_0335_),
    .B1_N(_0338_),
    .X(_0346_));
 sky130_fd_sc_hd__o21a_1 _1756_ (.A1(net14),
    .A2(_0333_),
    .B1(_0346_),
    .X(_0138_));
 sky130_fd_sc_hd__o21ba_1 _1757_ (.A1(\gps_channel0.ca_nco.step[10] ),
    .A2(_0335_),
    .B1_N(_0338_),
    .X(_0347_));
 sky130_fd_sc_hd__o21a_1 _1758_ (.A1(net15),
    .A2(_0332_),
    .B1(_0347_),
    .X(_0139_));
 sky130_fd_sc_hd__o21ba_1 _1759_ (.A1(\gps_channel0.ca_nco.step[11] ),
    .A2(_0334_),
    .B1_N(_0338_),
    .X(_0348_));
 sky130_fd_sc_hd__o21a_1 _1760_ (.A1(net16),
    .A2(_0332_),
    .B1(_0348_),
    .X(_0140_));
 sky130_fd_sc_hd__o21ba_1 _1761_ (.A1(\gps_channel0.ca_nco.step[12] ),
    .A2(_0334_),
    .B1_N(_0338_),
    .X(_0349_));
 sky130_fd_sc_hd__o21a_1 _1762_ (.A1(net17),
    .A2(_0332_),
    .B1(_0349_),
    .X(_0141_));
 sky130_fd_sc_hd__buf_2 _1763_ (.A(net3),
    .X(_0350_));
 sky130_fd_sc_hd__o21ba_1 _1764_ (.A1(\gps_channel0.ca_nco.step[13] ),
    .A2(_0334_),
    .B1_N(_0350_),
    .X(_0351_));
 sky130_fd_sc_hd__o21a_1 _1765_ (.A1(net18),
    .A2(_0332_),
    .B1(_0351_),
    .X(_0142_));
 sky130_fd_sc_hd__o21ba_1 _1766_ (.A1(\gps_channel0.ca_nco.step[14] ),
    .A2(_0334_),
    .B1_N(_0350_),
    .X(_0352_));
 sky130_fd_sc_hd__o21a_1 _1767_ (.A1(net20),
    .A2(_0332_),
    .B1(_0352_),
    .X(_0143_));
 sky130_fd_sc_hd__o21ba_1 _1768_ (.A1(\gps_channel0.ca_nco.step[15] ),
    .A2(_0334_),
    .B1_N(_0350_),
    .X(_0353_));
 sky130_fd_sc_hd__o21a_1 _1769_ (.A1(net21),
    .A2(_0332_),
    .B1(_0353_),
    .X(_0144_));
 sky130_fd_sc_hd__a21o_1 _1770_ (.A1(_0604_),
    .A2(_0332_),
    .B1(_0283_),
    .X(_0145_));
 sky130_fd_sc_hd__or3_1 _1771_ (.A(_0302_),
    .B(net23),
    .C(net24),
    .X(_0354_));
 sky130_fd_sc_hd__buf_2 _1772_ (.A(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__clkbuf_4 _1773_ (.A(_0355_),
    .X(_0356_));
 sky130_fd_sc_hd__o21ba_1 _1774_ (.A1(\gps_channel0.ca_nco.phase_in[0] ),
    .A2(_0305_),
    .B1_N(_0350_),
    .X(_0357_));
 sky130_fd_sc_hd__o21a_1 _1775_ (.A1(net4),
    .A2(_0356_),
    .B1(_0357_),
    .X(_0146_));
 sky130_fd_sc_hd__o21ba_1 _1776_ (.A1(\gps_channel0.ca_nco.phase_in[1] ),
    .A2(_0305_),
    .B1_N(_0350_),
    .X(_0358_));
 sky130_fd_sc_hd__o21a_1 _1777_ (.A1(net5),
    .A2(_0356_),
    .B1(_0358_),
    .X(_0147_));
 sky130_fd_sc_hd__o21ba_1 _1778_ (.A1(\gps_channel0.ca_nco.phase_in[2] ),
    .A2(_0305_),
    .B1_N(_0350_),
    .X(_0359_));
 sky130_fd_sc_hd__o21a_1 _1779_ (.A1(net6),
    .A2(_0356_),
    .B1(_0359_),
    .X(_0148_));
 sky130_fd_sc_hd__o21ba_1 _1780_ (.A1(\gps_channel0.ca_nco.phase_in[3] ),
    .A2(_0305_),
    .B1_N(_0350_),
    .X(_0360_));
 sky130_fd_sc_hd__o21a_1 _1781_ (.A1(net7),
    .A2(_0356_),
    .B1(_0360_),
    .X(_0149_));
 sky130_fd_sc_hd__o21ba_1 _1782_ (.A1(\gps_channel0.ca_nco.phase_in[4] ),
    .A2(_0305_),
    .B1_N(_0350_),
    .X(_0361_));
 sky130_fd_sc_hd__o21a_1 _1783_ (.A1(net9),
    .A2(_0356_),
    .B1(_0361_),
    .X(_0150_));
 sky130_fd_sc_hd__o21ba_1 _1784_ (.A1(\gps_channel0.ca_nco.phase_in[5] ),
    .A2(_0305_),
    .B1_N(_0350_),
    .X(_0362_));
 sky130_fd_sc_hd__o21a_1 _1785_ (.A1(net10),
    .A2(_0356_),
    .B1(_0362_),
    .X(_0151_));
 sky130_fd_sc_hd__inv_2 _1786_ (.A(\gps_channel0.ca_nco.phase_in[6] ),
    .Y(_0363_));
 sky130_fd_sc_hd__a21oi_1 _1787_ (.A1(_0363_),
    .A2(_0355_),
    .B1(_0283_),
    .Y(_0364_));
 sky130_fd_sc_hd__o21a_1 _1788_ (.A1(net11),
    .A2(_0356_),
    .B1(_0364_),
    .X(_0152_));
 sky130_fd_sc_hd__o21ba_1 _1789_ (.A1(\gps_channel0.ca_nco.phase_in[7] ),
    .A2(_0305_),
    .B1_N(_0350_),
    .X(_0365_));
 sky130_fd_sc_hd__o21a_1 _1790_ (.A1(net12),
    .A2(_0356_),
    .B1(_0365_),
    .X(_0153_));
 sky130_fd_sc_hd__o21ba_1 _1791_ (.A1(\gps_channel0.ca_nco.phase_in[8] ),
    .A2(_0305_),
    .B1_N(_0174_),
    .X(_0366_));
 sky130_fd_sc_hd__o21a_1 _1792_ (.A1(net13),
    .A2(_0356_),
    .B1(_0366_),
    .X(_0154_));
 sky130_fd_sc_hd__o21ba_1 _1793_ (.A1(\gps_channel0.ca_nco.phase_in[9] ),
    .A2(_0305_),
    .B1_N(_0174_),
    .X(_0367_));
 sky130_fd_sc_hd__o21a_1 _1794_ (.A1(net14),
    .A2(_0356_),
    .B1(_0367_),
    .X(_0155_));
 sky130_fd_sc_hd__o21ba_1 _1795_ (.A1(\gps_channel0.ca_nco.phase_in[10] ),
    .A2(_0304_),
    .B1_N(_0174_),
    .X(_0368_));
 sky130_fd_sc_hd__o21a_1 _1796_ (.A1(net15),
    .A2(_0355_),
    .B1(_0368_),
    .X(_0156_));
 sky130_fd_sc_hd__o21ba_1 _1797_ (.A1(\gps_channel0.ca_nco.phase_in[11] ),
    .A2(_0304_),
    .B1_N(_0174_),
    .X(_0369_));
 sky130_fd_sc_hd__o21a_1 _1798_ (.A1(net16),
    .A2(_0355_),
    .B1(_0369_),
    .X(_0157_));
 sky130_fd_sc_hd__o21ba_1 _1799_ (.A1(\gps_channel0.ca_nco.phase_in[12] ),
    .A2(_0304_),
    .B1_N(_0174_),
    .X(_0370_));
 sky130_fd_sc_hd__o21a_1 _1800_ (.A1(net17),
    .A2(_0355_),
    .B1(_0370_),
    .X(_0158_));
 sky130_fd_sc_hd__o21ba_1 _1801_ (.A1(\gps_channel0.ca_nco.phase_in[13] ),
    .A2(_0304_),
    .B1_N(_0174_),
    .X(_0371_));
 sky130_fd_sc_hd__o21a_1 _1802_ (.A1(net18),
    .A2(_0355_),
    .B1(_0371_),
    .X(_0159_));
 sky130_fd_sc_hd__o21ba_1 _1803_ (.A1(\gps_channel0.ca_nco.phase_in[14] ),
    .A2(_0304_),
    .B1_N(_0174_),
    .X(_0372_));
 sky130_fd_sc_hd__o21a_1 _1804_ (.A1(net20),
    .A2(_0355_),
    .B1(_0372_),
    .X(_0160_));
 sky130_fd_sc_hd__o21ba_1 _1805_ (.A1(\gps_channel0.ca_nco.phase_in[15] ),
    .A2(_0304_),
    .B1_N(_0174_),
    .X(_0373_));
 sky130_fd_sc_hd__o21a_1 _1806_ (.A1(net21),
    .A2(_0355_),
    .B1(_0373_),
    .X(_0161_));
 sky130_fd_sc_hd__dfxtp_1 _1807_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0010_),
    .Q(\gps_channel0.lo_nco.accumulator[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1808_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0011_),
    .Q(\gps_channel0.lo_nco.accumulator[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1809_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0012_),
    .Q(\gps_channel0.lo_nco.accumulator[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1810_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0013_),
    .Q(\gps_channel0.lo_nco.accumulator[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1811_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0014_),
    .Q(\gps_channel0.lo_nco.accumulator[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1812_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0015_),
    .Q(\gps_channel0.lo_nco.accumulator[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1813_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0016_),
    .Q(\gps_channel0.lo_nco.accumulator[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1814_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0017_),
    .Q(\gps_channel0.lo_nco.accumulator[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1815_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0018_),
    .Q(\gps_channel0.lo_nco.accumulator[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1816_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0019_),
    .Q(\gps_channel0.lo_nco.accumulator[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1817_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0020_),
    .Q(\gps_channel0.lo_nco.accumulator[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1818_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0021_),
    .Q(\gps_channel0.lo_nco.accumulator[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1819_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0022_),
    .Q(\gps_channel0.lo_nco.accumulator[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1820_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0023_),
    .Q(\gps_channel0.lo_nco.accumulator[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1821_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0024_),
    .Q(\gps_channel0.lo_nco.accumulator[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1822_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0025_),
    .Q(\gps_channel0.lo_nco.accumulator[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1823_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0026_),
    .Q(\gps_channel0.ca_nco.accumulator[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1824_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0027_),
    .Q(\gps_channel0.ca_nco.accumulator[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1825_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0028_),
    .Q(\gps_channel0.ca_nco.accumulator[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1826_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0029_),
    .Q(\gps_channel0.ca_nco.accumulator[19] ));
 sky130_fd_sc_hd__dfxtp_1 _1827_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0030_),
    .Q(\gps_channel0.ca_nco.accumulator[20] ));
 sky130_fd_sc_hd__dfxtp_1 _1828_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0031_),
    .Q(\gps_channel0.ca_nco.accumulator[21] ));
 sky130_fd_sc_hd__dfxtp_1 _1829_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0032_),
    .Q(\gps_channel0.ca_nco.accumulator[22] ));
 sky130_fd_sc_hd__dfxtp_1 _1830_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0033_),
    .Q(\gps_channel0.ca_nco.accumulator[23] ));
 sky130_fd_sc_hd__dfxtp_1 _1831_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0034_),
    .Q(\gps_channel0.ca_nco.accumulator[24] ));
 sky130_fd_sc_hd__dfxtp_1 _1832_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0035_),
    .Q(\gps_channel0.ca_nco.accumulator[25] ));
 sky130_fd_sc_hd__dfxtp_1 _1833_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0036_),
    .Q(\gps_channel0.ca_nco.accumulator[26] ));
 sky130_fd_sc_hd__dfxtp_1 _1834_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0037_),
    .Q(\gps_channel0.ca_nco.accumulator[27] ));
 sky130_fd_sc_hd__dfxtp_1 _1835_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0038_),
    .Q(\gps_channel0.ca_nco.accumulator[28] ));
 sky130_fd_sc_hd__dfxtp_1 _1836_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0039_),
    .Q(\gps_channel0.ca_nco.accumulator[29] ));
 sky130_fd_sc_hd__dfxtp_1 _1837_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0040_),
    .Q(\gps_channel0.ca_nco.accumulator[30] ));
 sky130_fd_sc_hd__dfxtp_1 _1838_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0041_),
    .Q(\gps_channel0.ca_full_chip ));
 sky130_fd_sc_hd__dfxtp_1 _1839_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0042_),
    .Q(\gps_channel0.ca_nco.accumulator[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1840_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0043_),
    .Q(\gps_channel0.ca_nco.accumulator[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1841_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0044_),
    .Q(\gps_channel0.ca_nco.accumulator[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1842_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0045_),
    .Q(\gps_channel0.ca_nco.accumulator[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1843_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0046_),
    .Q(\gps_channel0.ca_nco.accumulator[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1844_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0047_),
    .Q(\gps_channel0.ca_nco.accumulator[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1845_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0048_),
    .Q(\gps_channel0.ca_nco.accumulator[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1846_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0049_),
    .Q(\gps_channel0.ca_nco.accumulator[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1847_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0050_),
    .Q(\gps_channel0.ca_nco.accumulator[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1848_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0051_),
    .Q(\gps_channel0.ca_nco.accumulator[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1849_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0052_),
    .Q(\gps_channel0.ca_nco.accumulator[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1850_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0053_),
    .Q(\gps_channel0.ca_nco.accumulator[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1851_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0054_),
    .Q(\gps_channel0.ca_nco.accumulator[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1852_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0055_),
    .Q(\gps_channel0.ca_nco.accumulator[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1853_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0056_),
    .Q(\gps_channel0.ca_nco.accumulator[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1854_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0057_),
    .Q(\gps_channel0.ca_nco.accumulator[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1855_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0058_),
    .Q(\gps_channel0.lo_nco.phase_in[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1856_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0059_),
    .Q(\gps_channel0.lo_nco.phase_in[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1857_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0060_),
    .Q(\gps_channel0.lo_nco.phase_in[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1858_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0061_),
    .Q(\gps_channel0.lo_nco.phase_in[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1859_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0062_),
    .Q(\gps_channel0.lo_nco.phase_in[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1860_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0063_),
    .Q(\gps_channel0.lo_nco.phase_in[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1861_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0064_),
    .Q(\gps_channel0.lo_nco.phase_in[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1862_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0065_),
    .Q(\gps_channel0.lo_nco.phase_in[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1863_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0066_),
    .Q(\gps_channel0.lo_nco.phase_in[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1864_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0067_),
    .Q(\gps_channel0.lo_nco.phase_in[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1865_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0068_),
    .Q(\gps_channel0.lo_nco.phase_in[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1866_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0069_),
    .Q(\gps_channel0.lo_nco.phase_in[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1867_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0070_),
    .Q(\gps_channel0.lo_nco.phase_in[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1868_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0071_),
    .Q(\gps_channel0.lo_nco.phase_in[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1869_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0072_),
    .Q(\gps_channel0.lo_nco.phase_in[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1870_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0073_),
    .Q(\gps_channel0.lo_nco.phase_in[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1871_ (.CLK(net27),
    .D(_0000_),
    .Q(\gps_channel0.ca_gen.g2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1872_ (.CLK(net27),
    .D(_0001_),
    .Q(\gps_channel0.ca_gen.g2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1873_ (.CLK(net27),
    .D(_0002_),
    .Q(\gps_channel0.ca_gen.g2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1874_ (.CLK(net27),
    .D(_0003_),
    .Q(\gps_channel0.ca_gen.g2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1875_ (.CLK(net26),
    .D(_0004_),
    .Q(\gps_channel0.ca_gen.g2[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1876_ (.CLK(net26),
    .D(_0005_),
    .Q(\gps_channel0.ca_gen.g2[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1877_ (.CLK(net26),
    .D(_0006_),
    .Q(\gps_channel0.ca_gen.g2[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1878_ (.CLK(net27),
    .D(_0007_),
    .Q(\gps_channel0.ca_gen.g2[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1879_ (.CLK(net26),
    .D(_0008_),
    .Q(\gps_channel0.ca_gen.g2[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1880_ (.CLK(net26),
    .D(_0009_),
    .Q(\gps_channel0.ca_gen.g2[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1881_ (.CLK(net28),
    .D(_0074_),
    .Q(\gps_channel0.ca_gen.g1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1882_ (.CLK(net28),
    .D(_0075_),
    .Q(\gps_channel0.ca_gen.g1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1883_ (.CLK(net28),
    .D(_0076_),
    .Q(\gps_channel0.ca_gen.g1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1884_ (.CLK(net28),
    .D(_0077_),
    .Q(\gps_channel0.ca_gen.g1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1885_ (.CLK(net28),
    .D(_0078_),
    .Q(\gps_channel0.ca_gen.g1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1886_ (.CLK(net28),
    .D(_0079_),
    .Q(\gps_channel0.ca_gen.g1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1887_ (.CLK(net26),
    .D(_0080_),
    .Q(\gps_channel0.ca_gen.g1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1888_ (.CLK(net26),
    .D(_0081_),
    .Q(\gps_channel0.ca_gen.g1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1889_ (.CLK(net26),
    .D(_0082_),
    .Q(\gps_channel0.ca_gen.g1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1890_ (.CLK(net26),
    .D(_0083_),
    .Q(\gps_channel0.ca_gen.g1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1891_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0084_),
    .Q(\gps_channel0.lo_nco.accumulator[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1892_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0085_),
    .Q(\gps_channel0.lo_nco.accumulator[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1893_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0086_),
    .Q(\gps_channel0.lo_nco.accumulator[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1894_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0087_),
    .Q(\gps_channel0.lo_nco.accumulator[19] ));
 sky130_fd_sc_hd__dfxtp_1 _1895_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0088_),
    .Q(\gps_channel0.lo_nco.accumulator[20] ));
 sky130_fd_sc_hd__dfxtp_1 _1896_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0089_),
    .Q(\gps_channel0.lo_nco.accumulator[21] ));
 sky130_fd_sc_hd__dfxtp_1 _1897_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0090_),
    .Q(\gps_channel0.lo_nco.accumulator[22] ));
 sky130_fd_sc_hd__dfxtp_1 _1898_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0091_),
    .Q(\gps_channel0.lo_nco.accumulator[23] ));
 sky130_fd_sc_hd__dfxtp_1 _1899_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0092_),
    .Q(\gps_channel0.lo_nco.accumulator[24] ));
 sky130_fd_sc_hd__dfxtp_1 _1900_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0093_),
    .Q(\gps_channel0.lo_nco.accumulator[25] ));
 sky130_fd_sc_hd__dfxtp_1 _1901_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0094_),
    .Q(\gps_channel0.lo_nco.accumulator[26] ));
 sky130_fd_sc_hd__dfxtp_1 _1902_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0095_),
    .Q(\gps_channel0.lo_nco.accumulator[27] ));
 sky130_fd_sc_hd__dfxtp_1 _1903_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0096_),
    .Q(\gps_channel0.lo_nco.accumulator[28] ));
 sky130_fd_sc_hd__dfxtp_1 _1904_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0097_),
    .Q(\gps_channel0.lo_nco.accumulator[29] ));
 sky130_fd_sc_hd__dfxtp_2 _1905_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0098_),
    .Q(\gps_channel0.lo_nco.accumulator[30] ));
 sky130_fd_sc_hd__dfxtp_4 _1906_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0099_),
    .Q(\gps_channel0.lo_i ));
 sky130_fd_sc_hd__dfxtp_1 _1907_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0100_),
    .Q(\gps_channel0.ca_gen.g2_init[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1908_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0101_),
    .Q(\gps_channel0.ca_gen.g2_init[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1909_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0102_),
    .Q(\gps_channel0.ca_gen.g2_init[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1910_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0103_),
    .Q(\gps_channel0.ca_gen.g2_init[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1911_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0104_),
    .Q(\gps_channel0.ca_gen.g2_init[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1912_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0105_),
    .Q(\gps_channel0.ca_gen.g2_init[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1913_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0106_),
    .Q(\gps_channel0.ca_gen.g2_init[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1914_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0107_),
    .Q(\gps_channel0.ca_gen.g2_init[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1915_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0108_),
    .Q(\gps_channel0.ca_gen.g2_init[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1916_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0109_),
    .Q(\gps_channel0.ca_gen.g2_init[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1917_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0110_),
    .Q(\gps_channel0.ca_nco.phase_sync ));
 sky130_fd_sc_hd__dfxtp_1 _1918_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0111_),
    .Q(\gps_channel0.lo_nco.phase_sync ));
 sky130_fd_sc_hd__dfxtp_1 _1919_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0112_),
    .Q(\gps_channel0.lo_nco.step[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1920_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0113_),
    .Q(\gps_channel0.lo_nco.step[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1921_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0114_),
    .Q(\gps_channel0.lo_nco.step[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1922_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0115_),
    .Q(\gps_channel0.lo_nco.step[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1923_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0116_),
    .Q(\gps_channel0.lo_nco.step[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1924_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0117_),
    .Q(\gps_channel0.lo_nco.step[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1925_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0118_),
    .Q(\gps_channel0.lo_nco.step[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1926_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0119_),
    .Q(\gps_channel0.lo_nco.step[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1927_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0120_),
    .Q(\gps_channel0.lo_nco.step[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1928_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0121_),
    .Q(\gps_channel0.lo_nco.step[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1929_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0122_),
    .Q(\gps_channel0.lo_nco.step[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1930_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0123_),
    .Q(\gps_channel0.lo_nco.step[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1931_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0124_),
    .Q(\gps_channel0.lo_nco.step[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1932_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0125_),
    .Q(\gps_channel0.lo_nco.step[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1933_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0126_),
    .Q(\gps_channel0.lo_nco.step[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1934_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0127_),
    .Q(\gps_channel0.lo_nco.step[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1935_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0128_),
    .Q(\gps_channel0.lo_nco.step[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1936_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0129_),
    .Q(\gps_channel0.ca_nco.step[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1937_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0130_),
    .Q(\gps_channel0.ca_nco.step[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1938_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0131_),
    .Q(\gps_channel0.ca_nco.step[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1939_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0132_),
    .Q(\gps_channel0.ca_nco.step[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1940_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0133_),
    .Q(\gps_channel0.ca_nco.step[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1941_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0134_),
    .Q(\gps_channel0.ca_nco.step[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1942_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0135_),
    .Q(\gps_channel0.ca_nco.step[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1943_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0136_),
    .Q(\gps_channel0.ca_nco.step[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1944_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0137_),
    .Q(\gps_channel0.ca_nco.step[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1945_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0138_),
    .Q(\gps_channel0.ca_nco.step[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1946_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0139_),
    .Q(\gps_channel0.ca_nco.step[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1947_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0140_),
    .Q(\gps_channel0.ca_nco.step[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1948_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0141_),
    .Q(\gps_channel0.ca_nco.step[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1949_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0142_),
    .Q(\gps_channel0.ca_nco.step[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1950_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0143_),
    .Q(\gps_channel0.ca_nco.step[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1951_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0144_),
    .Q(\gps_channel0.ca_nco.step[15] ));
 sky130_fd_sc_hd__dfxtp_2 _1952_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0145_),
    .Q(\gps_channel0.ca_nco.step[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1953_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0146_),
    .Q(\gps_channel0.ca_nco.phase_in[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1954_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0147_),
    .Q(\gps_channel0.ca_nco.phase_in[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1955_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0148_),
    .Q(\gps_channel0.ca_nco.phase_in[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1956_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0149_),
    .Q(\gps_channel0.ca_nco.phase_in[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1957_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0150_),
    .Q(\gps_channel0.ca_nco.phase_in[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1958_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0151_),
    .Q(\gps_channel0.ca_nco.phase_in[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1959_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0152_),
    .Q(\gps_channel0.ca_nco.phase_in[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1960_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0153_),
    .Q(\gps_channel0.ca_nco.phase_in[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1961_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0154_),
    .Q(\gps_channel0.ca_nco.phase_in[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1962_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0155_),
    .Q(\gps_channel0.ca_nco.phase_in[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1963_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0156_),
    .Q(\gps_channel0.ca_nco.phase_in[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1964_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0157_),
    .Q(\gps_channel0.ca_nco.phase_in[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1965_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0158_),
    .Q(\gps_channel0.ca_nco.phase_in[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1966_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0159_),
    .Q(\gps_channel0.ca_nco.phase_in[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1967_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0160_),
    .Q(\gps_channel0.ca_nco.phase_in[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1968_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0161_),
    .Q(\gps_channel0.ca_nco.phase_in[15] ));
 sky130_fd_sc_hd__conb_1 _2067__30 (.LO(net30));
 sky130_fd_sc_hd__conb_1 _2068__31 (.LO(net31));
 sky130_fd_sc_hd__conb_1 _2069__32 (.LO(net32));
 sky130_fd_sc_hd__conb_1 _2070__33 (.LO(net33));
 sky130_fd_sc_hd__conb_1 _2071__34 (.LO(net34));
 sky130_fd_sc_hd__conb_1 _2072__35 (.LO(net35));
 sky130_fd_sc_hd__conb_1 _2082__36 (.LO(net36));
 sky130_fd_sc_hd__conb_1 _2083__37 (.LO(net37));
 sky130_fd_sc_hd__conb_1 _2084__38 (.LO(net38));
 sky130_fd_sc_hd__conb_1 _2085__39 (.LO(net39));
 sky130_fd_sc_hd__conb_1 _2086__40 (.LO(net40));
 sky130_fd_sc_hd__conb_1 _2087__41 (.LO(net41));
 sky130_fd_sc_hd__conb_1 _2088__42 (.LO(net42));
 sky130_fd_sc_hd__conb_1 _2089__43 (.LO(net43));
 sky130_fd_sc_hd__conb_1 _2090__44 (.LO(net44));
 sky130_fd_sc_hd__conb_1 _2091__45 (.LO(net45));
 sky130_fd_sc_hd__conb_1 _2092__46 (.LO(net46));
 sky130_fd_sc_hd__conb_1 _2093__47 (.LO(net47));
 sky130_fd_sc_hd__conb_1 _2094__48 (.LO(net48));
 sky130_fd_sc_hd__conb_1 _2095__49 (.LO(net49));
 sky130_fd_sc_hd__conb_1 _2096__50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 _2097__51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 _2098__52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 _2099__53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 _2100__54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 _2101__55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 _2102__56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 _2103__57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 _2104__58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 _2105__59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 _2106__60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 _2107__61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 _2108__62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 _2109__63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 _2110__64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 _2111__65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 _2112__66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 _2113__67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 _2114__68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 _2115__69 (.LO(net69));
 sky130_fd_sc_hd__conb_1 _2116__70 (.LO(net70));
 sky130_fd_sc_hd__conb_1 _2118__71 (.LO(net71));
 sky130_fd_sc_hd__conb_1 _2120__72 (.LO(net72));
 sky130_fd_sc_hd__conb_1 _2121__73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 _2122__74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 _2123__75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 _2124__76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 _2125__77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 _2126__78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 _2127__79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 _2128__80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 _2129__81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 _2130__82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 _2131__83 (.LO(net83));
 sky130_fd_sc_hd__conb_1 _2132__84 (.LO(net84));
 sky130_fd_sc_hd__conb_1 _2133__85 (.LO(net85));
 sky130_fd_sc_hd__conb_1 _2134__86 (.LO(net86));
 sky130_fd_sc_hd__conb_1 _2135__87 (.LO(net87));
 sky130_fd_sc_hd__conb_1 _2136__88 (.LO(net88));
 sky130_fd_sc_hd__conb_1 _2137__89 (.LO(net89));
 sky130_fd_sc_hd__conb_1 _2138__90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 _2139__91 (.LO(net91));
 sky130_fd_sc_hd__conb_1 _2140__92 (.LO(net92));
 sky130_fd_sc_hd__conb_1 _2141__93 (.LO(net93));
 sky130_fd_sc_hd__conb_1 _2142__94 (.LO(net94));
 sky130_fd_sc_hd__conb_1 _2143__95 (.LO(net95));
 sky130_fd_sc_hd__conb_1 _2144__96 (.LO(net96));
 sky130_fd_sc_hd__conb_1 _2145__97 (.LO(net97));
 sky130_fd_sc_hd__conb_1 _2146__98 (.LO(net98));
 sky130_fd_sc_hd__conb_1 _2147__99 (.LO(net99));
 sky130_fd_sc_hd__conb_1 _2148__100 (.LO(net100));
 sky130_fd_sc_hd__conb_1 _2149__101 (.LO(net101));
 sky130_fd_sc_hd__conb_1 _2150__102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 _2151__103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 _2152__104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 _2153__105 (.LO(net105));
 sky130_fd_sc_hd__conb_1 _2154__106 (.LO(net106));
 sky130_fd_sc_hd__conb_1 _2155__107 (.LO(net107));
 sky130_fd_sc_hd__conb_1 _2156__108 (.LO(net108));
 sky130_fd_sc_hd__conb_1 _2157__109 (.LO(net109));
 sky130_fd_sc_hd__conb_1 _2158__110 (.LO(net110));
 sky130_fd_sc_hd__conb_1 _2159__111 (.LO(net111));
 sky130_fd_sc_hd__conb_1 _2160__112 (.LO(net112));
 sky130_fd_sc_hd__conb_1 _2161__113 (.LO(net113));
 sky130_fd_sc_hd__conb_1 _2162__114 (.LO(net114));
 sky130_fd_sc_hd__conb_1 _2163__115 (.LO(net115));
 sky130_fd_sc_hd__conb_1 _2164__116 (.LO(net116));
 sky130_fd_sc_hd__conb_1 _2165__117 (.LO(net117));
 sky130_fd_sc_hd__conb_1 _2166__118 (.LO(net118));
 sky130_fd_sc_hd__conb_1 _2167__119 (.LO(net119));
 sky130_fd_sc_hd__conb_1 _2168__120 (.LO(net120));
 sky130_fd_sc_hd__conb_1 _2169__121 (.LO(net121));
 sky130_fd_sc_hd__conb_1 _2170__122 (.LO(net122));
 sky130_fd_sc_hd__conb_1 _2171__123 (.LO(net123));
 sky130_fd_sc_hd__conb_1 _2172__124 (.LO(net124));
 sky130_fd_sc_hd__conb_1 _2173__125 (.LO(net125));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__ebufn_8 _2066_ (.A(net29),
    .TE_B(_0746_),
    .Z(la1_data_out[0]));
 sky130_fd_sc_hd__ebufn_8 _2067_ (.A(net30),
    .TE_B(_0747_),
    .Z(la1_data_out[1]));
 sky130_fd_sc_hd__ebufn_8 _2068_ (.A(net31),
    .TE_B(_0748_),
    .Z(la1_data_out[2]));
 sky130_fd_sc_hd__ebufn_8 _2069_ (.A(net32),
    .TE_B(_0749_),
    .Z(la1_data_out[3]));
 sky130_fd_sc_hd__ebufn_8 _2070_ (.A(net33),
    .TE_B(_0750_),
    .Z(la1_data_out[4]));
 sky130_fd_sc_hd__ebufn_8 _2071_ (.A(net34),
    .TE_B(_0751_),
    .Z(la1_data_out[5]));
 sky130_fd_sc_hd__ebufn_8 _2072_ (.A(net35),
    .TE_B(_0752_),
    .Z(la1_data_out[6]));
 sky130_fd_sc_hd__ebufn_8 _2073_ (.A(\gps_channel0.prompt_q ),
    .TE_B(_0753_),
    .Z(la1_data_out[7]));
 sky130_fd_sc_hd__ebufn_8 _2074_ (.A(\gps_channel0.lo_nco.accumulator[28] ),
    .TE_B(_0754_),
    .Z(la1_data_out[8]));
 sky130_fd_sc_hd__ebufn_8 _2075_ (.A(\gps_channel0.lo_nco.accumulator[29] ),
    .TE_B(_0755_),
    .Z(la1_data_out[9]));
 sky130_fd_sc_hd__ebufn_8 _2076_ (.A(\gps_channel0.lo_nco.accumulator[30] ),
    .TE_B(_0756_),
    .Z(la1_data_out[10]));
 sky130_fd_sc_hd__ebufn_8 _2077_ (.A(\gps_channel0.lo_i ),
    .TE_B(_0757_),
    .Z(la1_data_out[11]));
 sky130_fd_sc_hd__ebufn_8 _2078_ (.A(\gps_channel0.ca_nco.accumulator[28] ),
    .TE_B(_0758_),
    .Z(la1_data_out[12]));
 sky130_fd_sc_hd__ebufn_8 _2079_ (.A(\gps_channel0.ca_nco.accumulator[29] ),
    .TE_B(_0759_),
    .Z(la1_data_out[13]));
 sky130_fd_sc_hd__ebufn_8 _2080_ (.A(\gps_channel0.ca_nco.accumulator[30] ),
    .TE_B(_0760_),
    .Z(la1_data_out[14]));
 sky130_fd_sc_hd__ebufn_8 _2081_ (.A(net26),
    .TE_B(_0761_),
    .Z(la1_data_out[15]));
 sky130_fd_sc_hd__ebufn_8 _2082_ (.A(net36),
    .TE_B(_0762_),
    .Z(la1_data_out[16]));
 sky130_fd_sc_hd__ebufn_8 _2083_ (.A(net37),
    .TE_B(_0763_),
    .Z(la1_data_out[17]));
 sky130_fd_sc_hd__ebufn_8 _2084_ (.A(net38),
    .TE_B(_0764_),
    .Z(la1_data_out[18]));
 sky130_fd_sc_hd__ebufn_8 _2085_ (.A(net39),
    .TE_B(_0765_),
    .Z(la1_data_out[19]));
 sky130_fd_sc_hd__ebufn_8 _2086_ (.A(net40),
    .TE_B(_0766_),
    .Z(la1_data_out[20]));
 sky130_fd_sc_hd__ebufn_8 _2087_ (.A(net41),
    .TE_B(_0767_),
    .Z(la1_data_out[21]));
 sky130_fd_sc_hd__ebufn_8 _2088_ (.A(net42),
    .TE_B(_0768_),
    .Z(la1_data_out[22]));
 sky130_fd_sc_hd__ebufn_8 _2089_ (.A(net43),
    .TE_B(_0769_),
    .Z(la1_data_out[23]));
 sky130_fd_sc_hd__ebufn_8 _2090_ (.A(net44),
    .TE_B(_0770_),
    .Z(la1_data_out[24]));
 sky130_fd_sc_hd__ebufn_8 _2091_ (.A(net45),
    .TE_B(_0771_),
    .Z(la1_data_out[25]));
 sky130_fd_sc_hd__ebufn_8 _2092_ (.A(net46),
    .TE_B(_0772_),
    .Z(la1_data_out[26]));
 sky130_fd_sc_hd__ebufn_8 _2093_ (.A(net47),
    .TE_B(_0773_),
    .Z(la1_data_out[27]));
 sky130_fd_sc_hd__ebufn_8 _2094_ (.A(net48),
    .TE_B(_0774_),
    .Z(la1_data_out[28]));
 sky130_fd_sc_hd__ebufn_8 _2095_ (.A(net49),
    .TE_B(_0775_),
    .Z(la1_data_out[29]));
 sky130_fd_sc_hd__ebufn_8 _2096_ (.A(net50),
    .TE_B(_0776_),
    .Z(la1_data_out[30]));
 sky130_fd_sc_hd__ebufn_8 _2097_ (.A(net51),
    .TE_B(_0777_),
    .Z(la1_data_out[31]));
 sky130_fd_sc_hd__ebufn_8 _2098_ (.A(net52),
    .TE_B(_0778_),
    .Z(io_out[0]));
 sky130_fd_sc_hd__ebufn_8 _2099_ (.A(net53),
    .TE_B(_0779_),
    .Z(io_out[1]));
 sky130_fd_sc_hd__ebufn_8 _2100_ (.A(net54),
    .TE_B(_0780_),
    .Z(io_out[2]));
 sky130_fd_sc_hd__ebufn_8 _2101_ (.A(net55),
    .TE_B(_0781_),
    .Z(io_out[3]));
 sky130_fd_sc_hd__ebufn_8 _2102_ (.A(net56),
    .TE_B(_0782_),
    .Z(io_out[4]));
 sky130_fd_sc_hd__ebufn_8 _2103_ (.A(net57),
    .TE_B(_0783_),
    .Z(io_out[5]));
 sky130_fd_sc_hd__ebufn_8 _2104_ (.A(net58),
    .TE_B(_0784_),
    .Z(io_out[6]));
 sky130_fd_sc_hd__ebufn_8 _2105_ (.A(net59),
    .TE_B(_0785_),
    .Z(io_out[7]));
 sky130_fd_sc_hd__ebufn_8 _2106_ (.A(net60),
    .TE_B(_0786_),
    .Z(io_out[8]));
 sky130_fd_sc_hd__ebufn_8 _2107_ (.A(net61),
    .TE_B(_0787_),
    .Z(io_out[9]));
 sky130_fd_sc_hd__ebufn_8 _2108_ (.A(net62),
    .TE_B(_0788_),
    .Z(io_out[10]));
 sky130_fd_sc_hd__ebufn_8 _2109_ (.A(net63),
    .TE_B(_0789_),
    .Z(io_out[11]));
 sky130_fd_sc_hd__ebufn_8 _2110_ (.A(net64),
    .TE_B(_0790_),
    .Z(io_out[12]));
 sky130_fd_sc_hd__ebufn_8 _2111_ (.A(net65),
    .TE_B(_0791_),
    .Z(io_out[13]));
 sky130_fd_sc_hd__ebufn_8 _2112_ (.A(net66),
    .TE_B(_0792_),
    .Z(io_out[14]));
 sky130_fd_sc_hd__ebufn_8 _2113_ (.A(net67),
    .TE_B(_0793_),
    .Z(io_out[15]));
 sky130_fd_sc_hd__ebufn_8 _2114_ (.A(net68),
    .TE_B(_0794_),
    .Z(io_out[16]));
 sky130_fd_sc_hd__ebufn_8 _2115_ (.A(net69),
    .TE_B(_0795_),
    .Z(io_out[17]));
 sky130_fd_sc_hd__ebufn_8 _2116_ (.A(net70),
    .TE_B(_0796_),
    .Z(io_out[18]));
 sky130_fd_sc_hd__ebufn_8 _2117_ (.A(\gps_channel0.lo_i ),
    .TE_B(_0797_),
    .Z(io_out[19]));
 sky130_fd_sc_hd__ebufn_8 _2118_ (.A(net71),
    .TE_B(_0798_),
    .Z(io_out[20]));
 sky130_fd_sc_hd__ebufn_8 _2119_ (.A(\gps_channel0.prompt_i ),
    .TE_B(_0799_),
    .Z(io_out[21]));
 sky130_fd_sc_hd__ebufn_8 _2120_ (.A(net72),
    .TE_B(_0800_),
    .Z(io_out[22]));
 sky130_fd_sc_hd__ebufn_8 _2121_ (.A(net73),
    .TE_B(_0801_),
    .Z(io_out[23]));
 sky130_fd_sc_hd__ebufn_8 _2122_ (.A(net74),
    .TE_B(_0802_),
    .Z(io_out[24]));
 sky130_fd_sc_hd__ebufn_8 _2123_ (.A(net75),
    .TE_B(_0803_),
    .Z(io_out[25]));
 sky130_fd_sc_hd__ebufn_8 _2124_ (.A(net76),
    .TE_B(_0804_),
    .Z(io_out[26]));
 sky130_fd_sc_hd__ebufn_8 _2125_ (.A(net77),
    .TE_B(_0805_),
    .Z(io_out[27]));
 sky130_fd_sc_hd__ebufn_8 _2126_ (.A(net78),
    .TE_B(_0806_),
    .Z(io_out[28]));
 sky130_fd_sc_hd__ebufn_8 _2127_ (.A(net79),
    .TE_B(_0807_),
    .Z(io_out[29]));
 sky130_fd_sc_hd__ebufn_8 _2128_ (.A(net80),
    .TE_B(_0808_),
    .Z(io_out[30]));
 sky130_fd_sc_hd__ebufn_8 _2129_ (.A(net81),
    .TE_B(_0809_),
    .Z(io_out[31]));
 sky130_fd_sc_hd__ebufn_8 _2130_ (.A(net82),
    .TE_B(_0810_),
    .Z(io_out[32]));
 sky130_fd_sc_hd__ebufn_8 _2131_ (.A(net83),
    .TE_B(_0811_),
    .Z(io_out[33]));
 sky130_fd_sc_hd__ebufn_8 _2132_ (.A(net84),
    .TE_B(_0812_),
    .Z(io_out[34]));
 sky130_fd_sc_hd__ebufn_8 _2133_ (.A(net85),
    .TE_B(_0813_),
    .Z(io_out[35]));
 sky130_fd_sc_hd__ebufn_8 _2134_ (.A(net86),
    .TE_B(_0814_),
    .Z(io_out[36]));
 sky130_fd_sc_hd__ebufn_8 _2135_ (.A(net87),
    .TE_B(_0815_),
    .Z(io_out[37]));
 sky130_fd_sc_hd__ebufn_8 _2136_ (.A(net88),
    .TE_B(_0816_),
    .Z(io_oeb[0]));
 sky130_fd_sc_hd__ebufn_8 _2137_ (.A(net89),
    .TE_B(_0817_),
    .Z(io_oeb[1]));
 sky130_fd_sc_hd__ebufn_8 _2138_ (.A(net90),
    .TE_B(_0818_),
    .Z(io_oeb[2]));
 sky130_fd_sc_hd__ebufn_8 _2139_ (.A(net91),
    .TE_B(_0819_),
    .Z(io_oeb[3]));
 sky130_fd_sc_hd__ebufn_8 _2140_ (.A(net92),
    .TE_B(_0820_),
    .Z(io_oeb[4]));
 sky130_fd_sc_hd__ebufn_8 _2141_ (.A(net93),
    .TE_B(_0821_),
    .Z(io_oeb[5]));
 sky130_fd_sc_hd__ebufn_8 _2142_ (.A(net94),
    .TE_B(_0822_),
    .Z(io_oeb[6]));
 sky130_fd_sc_hd__ebufn_8 _2143_ (.A(net95),
    .TE_B(_0823_),
    .Z(io_oeb[7]));
 sky130_fd_sc_hd__ebufn_8 _2144_ (.A(net96),
    .TE_B(_0824_),
    .Z(io_oeb[8]));
 sky130_fd_sc_hd__ebufn_8 _2145_ (.A(net97),
    .TE_B(_0825_),
    .Z(io_oeb[9]));
 sky130_fd_sc_hd__ebufn_8 _2146_ (.A(net98),
    .TE_B(_0826_),
    .Z(io_oeb[10]));
 sky130_fd_sc_hd__ebufn_8 _2147_ (.A(net99),
    .TE_B(_0827_),
    .Z(io_oeb[11]));
 sky130_fd_sc_hd__ebufn_8 _2148_ (.A(net100),
    .TE_B(_0828_),
    .Z(io_oeb[12]));
 sky130_fd_sc_hd__ebufn_8 _2149_ (.A(net101),
    .TE_B(_0829_),
    .Z(io_oeb[13]));
 sky130_fd_sc_hd__ebufn_8 _2150_ (.A(net102),
    .TE_B(_0830_),
    .Z(io_oeb[14]));
 sky130_fd_sc_hd__ebufn_8 _2151_ (.A(net103),
    .TE_B(_0831_),
    .Z(io_oeb[15]));
 sky130_fd_sc_hd__ebufn_8 _2152_ (.A(net104),
    .TE_B(_0832_),
    .Z(io_oeb[16]));
 sky130_fd_sc_hd__ebufn_8 _2153_ (.A(net105),
    .TE_B(_0833_),
    .Z(io_oeb[17]));
 sky130_fd_sc_hd__ebufn_8 _2154_ (.A(net106),
    .TE_B(_0834_),
    .Z(io_oeb[18]));
 sky130_fd_sc_hd__ebufn_8 _2155_ (.A(net107),
    .TE_B(_0835_),
    .Z(io_oeb[19]));
 sky130_fd_sc_hd__ebufn_8 _2156_ (.A(net108),
    .TE_B(_0836_),
    .Z(io_oeb[20]));
 sky130_fd_sc_hd__ebufn_8 _2157_ (.A(net109),
    .TE_B(_0837_),
    .Z(io_oeb[21]));
 sky130_fd_sc_hd__ebufn_8 _2158_ (.A(net110),
    .TE_B(_0838_),
    .Z(io_oeb[22]));
 sky130_fd_sc_hd__ebufn_8 _2159_ (.A(net111),
    .TE_B(_0839_),
    .Z(io_oeb[23]));
 sky130_fd_sc_hd__ebufn_8 _2160_ (.A(net112),
    .TE_B(_0840_),
    .Z(io_oeb[24]));
 sky130_fd_sc_hd__ebufn_8 _2161_ (.A(net113),
    .TE_B(_0841_),
    .Z(io_oeb[25]));
 sky130_fd_sc_hd__ebufn_8 _2162_ (.A(net114),
    .TE_B(_0842_),
    .Z(io_oeb[26]));
 sky130_fd_sc_hd__ebufn_8 _2163_ (.A(net115),
    .TE_B(_0843_),
    .Z(io_oeb[27]));
 sky130_fd_sc_hd__ebufn_8 _2164_ (.A(net116),
    .TE_B(_0844_),
    .Z(io_oeb[28]));
 sky130_fd_sc_hd__ebufn_8 _2165_ (.A(net117),
    .TE_B(_0845_),
    .Z(io_oeb[29]));
 sky130_fd_sc_hd__ebufn_8 _2166_ (.A(net118),
    .TE_B(_0846_),
    .Z(io_oeb[30]));
 sky130_fd_sc_hd__ebufn_8 _2167_ (.A(net119),
    .TE_B(_0847_),
    .Z(io_oeb[31]));
 sky130_fd_sc_hd__ebufn_8 _2168_ (.A(net120),
    .TE_B(_0848_),
    .Z(io_oeb[32]));
 sky130_fd_sc_hd__ebufn_8 _2169_ (.A(net121),
    .TE_B(_0849_),
    .Z(io_oeb[33]));
 sky130_fd_sc_hd__ebufn_8 _2170_ (.A(net122),
    .TE_B(_0850_),
    .Z(io_oeb[34]));
 sky130_fd_sc_hd__ebufn_8 _2171_ (.A(net123),
    .TE_B(_0851_),
    .Z(io_oeb[35]));
 sky130_fd_sc_hd__ebufn_8 _2172_ (.A(net124),
    .TE_B(_0852_),
    .Z(io_oeb[36]));
 sky130_fd_sc_hd__ebufn_8 _2173_ (.A(net125),
    .TE_B(_0853_),
    .Z(io_oeb[37]));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(active),
    .X(net1));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(io_in[23]),
    .X(net2));
 sky130_fd_sc_hd__buf_4 input3 (.A(la1_data_in[0]),
    .X(net3));
 sky130_fd_sc_hd__buf_2 input4 (.A(la1_data_in[16]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(la1_data_in[17]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(la1_data_in[18]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(la1_data_in[19]),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input8 (.A(la1_data_in[1]),
    .X(net8));
 sky130_fd_sc_hd__buf_2 input9 (.A(la1_data_in[20]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 input10 (.A(la1_data_in[21]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(la1_data_in[22]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 input12 (.A(la1_data_in[23]),
    .X(net12));
 sky130_fd_sc_hd__buf_2 input13 (.A(la1_data_in[24]),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input14 (.A(la1_data_in[25]),
    .X(net14));
 sky130_fd_sc_hd__buf_2 input15 (.A(la1_data_in[26]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(la1_data_in[27]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(la1_data_in[28]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(la1_data_in[29]),
    .X(net18));
 sky130_fd_sc_hd__buf_2 input19 (.A(la1_data_in[2]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(la1_data_in[30]),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(la1_data_in[31]),
    .X(net21));
 sky130_fd_sc_hd__dlymetal6s2s_1 input22 (.A(la1_data_in[3]),
    .X(net22));
 sky130_fd_sc_hd__buf_2 input23 (.A(la1_data_in[4]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(la1_data_in[5]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(la1_data_in[6]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_4 fanout26 (.A(net28),
    .X(net26));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout27 (.A(net28),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 fanout28 (.A(\gps_channel0.ca_full_chip ),
    .X(net28));
 sky130_fd_sc_hd__conb_1 _2066__29 (.LO(net29));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_4_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_5_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_6_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_7_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_8_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_9_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_10_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_11_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_12_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_13_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_14_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_15_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net10));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_514 ();
endmodule

