magic
tech sky130B
magscale 1 2
timestamp 1671924824
<< viali >>
rect 6561 47141 6595 47175
rect 9137 47141 9171 47175
rect 17693 47141 17727 47175
rect 19625 47141 19659 47175
rect 24777 47141 24811 47175
rect 42809 47141 42843 47175
rect 5089 47073 5123 47107
rect 14749 47073 14783 47107
rect 38301 47073 38335 47107
rect 46765 47073 46799 47107
rect 2697 47005 2731 47039
rect 3433 47005 3467 47039
rect 5549 47005 5583 47039
rect 9321 47005 9355 47039
rect 12449 47005 12483 47039
rect 13737 47005 13771 47039
rect 14289 47005 14323 47039
rect 17509 47005 17543 47039
rect 19441 47005 19475 47039
rect 22569 47005 22603 47039
rect 24593 47005 24627 47039
rect 25329 47005 25363 47039
rect 29837 47005 29871 47039
rect 32321 47005 32355 47039
rect 33149 47005 33183 47039
rect 38945 47005 38979 47039
rect 40141 47005 40175 47039
rect 41521 47005 41555 47039
rect 42625 47005 42659 47039
rect 47225 47005 47259 47039
rect 48237 47005 48271 47039
rect 2329 46937 2363 46971
rect 4077 46937 4111 46971
rect 4445 46937 4479 46971
rect 14473 46937 14507 46971
rect 47041 46937 47075 46971
rect 47869 46937 47903 46971
rect 3341 46869 3375 46903
rect 32505 46869 32539 46903
rect 7205 46665 7239 46699
rect 3525 46597 3559 46631
rect 4169 46597 4203 46631
rect 3709 46529 3743 46563
rect 6009 46529 6043 46563
rect 7389 46529 7423 46563
rect 12081 46529 12115 46563
rect 22477 46529 22511 46563
rect 24777 46529 24811 46563
rect 33057 46529 33091 46563
rect 39773 46529 39807 46563
rect 42625 46529 42659 46563
rect 47777 46529 47811 46563
rect 2605 46461 2639 46495
rect 5825 46461 5859 46495
rect 12265 46461 12299 46495
rect 13001 46461 13035 46495
rect 14381 46461 14415 46495
rect 14565 46461 14599 46495
rect 14841 46461 14875 46495
rect 22661 46461 22695 46495
rect 23213 46461 23247 46495
rect 24961 46461 24995 46495
rect 25789 46461 25823 46495
rect 28733 46461 28767 46495
rect 29193 46461 29227 46495
rect 29377 46461 29411 46495
rect 29653 46461 29687 46495
rect 33241 46461 33275 46495
rect 33517 46461 33551 46495
rect 36277 46461 36311 46495
rect 37473 46461 37507 46495
rect 37657 46461 37691 46495
rect 37933 46461 37967 46495
rect 39957 46461 39991 46495
rect 40233 46461 40267 46495
rect 42809 46461 42843 46495
rect 43085 46461 43119 46495
rect 45385 46461 45419 46495
rect 45569 46461 45603 46495
rect 46397 46461 46431 46495
rect 6561 46325 6595 46359
rect 10517 46325 10551 46359
rect 16865 46325 16899 46359
rect 35449 46325 35483 46359
rect 47869 46325 47903 46359
rect 6285 46121 6319 46155
rect 12909 46121 12943 46155
rect 13645 46121 13679 46155
rect 14473 46121 14507 46155
rect 22661 46121 22695 46155
rect 29101 46121 29135 46155
rect 33241 46121 33275 46155
rect 38393 46121 38427 46155
rect 45937 46121 45971 46155
rect 4445 46053 4479 46087
rect 2789 45985 2823 46019
rect 3249 45985 3283 46019
rect 10517 45985 10551 46019
rect 11069 45985 11103 46019
rect 15485 45985 15519 46019
rect 16865 45985 16899 46019
rect 25145 45985 25179 46019
rect 29745 45985 29779 46019
rect 30389 45985 30423 46019
rect 35357 45985 35391 46019
rect 36093 45985 36127 46019
rect 40141 45985 40175 46019
rect 40601 45985 40635 46019
rect 45385 45985 45419 46019
rect 46489 45985 46523 46019
rect 46673 45985 46707 46019
rect 48329 45985 48363 46019
rect 3433 45917 3467 45951
rect 6377 45917 6411 45951
rect 7021 45917 7055 45951
rect 13001 45917 13035 45951
rect 13553 45917 13587 45951
rect 14381 45917 14415 45951
rect 22569 45917 22603 45951
rect 23857 45917 23891 45951
rect 24593 45917 24627 45951
rect 29009 45917 29043 45951
rect 33149 45917 33183 45951
rect 38301 45917 38335 45951
rect 38945 45917 38979 45951
rect 46029 45917 46063 45951
rect 5733 45849 5767 45883
rect 10701 45849 10735 45883
rect 16681 45849 16715 45883
rect 23949 45849 23983 45883
rect 24777 45849 24811 45883
rect 29929 45849 29963 45883
rect 35541 45849 35575 45883
rect 40325 45849 40359 45883
rect 6929 45781 6963 45815
rect 39037 45781 39071 45815
rect 10609 45577 10643 45611
rect 25237 45577 25271 45611
rect 3801 45509 3835 45543
rect 29929 45509 29963 45543
rect 35633 45509 35667 45543
rect 36277 45509 36311 45543
rect 39129 45509 39163 45543
rect 41613 45509 41647 45543
rect 47133 45509 47167 45543
rect 4997 45441 5031 45475
rect 6745 45441 6779 45475
rect 10517 45441 10551 45475
rect 14473 45441 14507 45475
rect 15117 45441 15151 45475
rect 15209 45441 15243 45475
rect 24685 45441 24719 45475
rect 25329 45441 25363 45475
rect 29837 45441 29871 45475
rect 35725 45441 35759 45475
rect 36185 45441 36219 45475
rect 38945 45441 38979 45475
rect 41521 45441 41555 45475
rect 45937 45441 45971 45475
rect 47225 45441 47259 45475
rect 2881 45373 2915 45407
rect 3985 45373 4019 45407
rect 5457 45373 5491 45407
rect 7389 45373 7423 45407
rect 40785 45373 40819 45407
rect 47961 45237 47995 45271
rect 5273 45033 5307 45067
rect 40417 45033 40451 45067
rect 6837 44897 6871 44931
rect 46857 44897 46891 44931
rect 48329 44897 48363 44931
rect 1961 44829 1995 44863
rect 2421 44829 2455 44863
rect 3985 44829 4019 44863
rect 6193 44829 6227 44863
rect 40509 44829 40543 44863
rect 3249 44761 3283 44795
rect 48145 44761 48179 44795
rect 4445 44489 4479 44523
rect 47869 44489 47903 44523
rect 2053 44353 2087 44387
rect 4537 44353 4571 44387
rect 4997 44353 5031 44387
rect 47225 44353 47259 44387
rect 47777 44353 47811 44387
rect 2237 44285 2271 44319
rect 3157 44285 3191 44319
rect 5825 44285 5859 44319
rect 6745 44149 6779 44183
rect 3065 43809 3099 43843
rect 4629 43809 4663 43843
rect 5733 43809 5767 43843
rect 7297 43809 7331 43843
rect 1961 43741 1995 43775
rect 3433 43741 3467 43775
rect 4997 43741 5031 43775
rect 7113 43673 7147 43707
rect 5917 43401 5951 43435
rect 5181 43333 5215 43367
rect 2053 43265 2087 43299
rect 4537 43265 4571 43299
rect 6009 43265 6043 43299
rect 47777 43265 47811 43299
rect 2237 43197 2271 43231
rect 2789 43197 2823 43231
rect 47041 43061 47075 43095
rect 47869 43061 47903 43095
rect 2421 42857 2455 42891
rect 3065 42721 3099 42755
rect 46489 42721 46523 42755
rect 48237 42721 48271 42755
rect 2513 42653 2547 42687
rect 3157 42653 3191 42687
rect 5181 42653 5215 42687
rect 5733 42585 5767 42619
rect 46673 42585 46707 42619
rect 5641 41973 5675 42007
rect 47777 41973 47811 42007
rect 7297 41633 7331 41667
rect 46489 41633 46523 41667
rect 48237 41633 48271 41667
rect 5457 41497 5491 41531
rect 7113 41497 7147 41531
rect 46673 41497 46707 41531
rect 6653 41225 6687 41259
rect 47133 41225 47167 41259
rect 6561 41089 6595 41123
rect 47225 41089 47259 41123
rect 47777 40885 47811 40919
rect 46489 40545 46523 40579
rect 15853 40477 15887 40511
rect 18337 40477 18371 40511
rect 23673 40477 23707 40511
rect 23857 40477 23891 40511
rect 16037 40409 16071 40443
rect 17693 40409 17727 40443
rect 46673 40409 46707 40443
rect 48329 40409 48363 40443
rect 18245 40341 18279 40375
rect 23765 40341 23799 40375
rect 16037 40137 16071 40171
rect 22293 40137 22327 40171
rect 13001 40069 13035 40103
rect 17785 40069 17819 40103
rect 22109 40069 22143 40103
rect 15945 40001 15979 40035
rect 22017 40001 22051 40035
rect 22385 40001 22419 40035
rect 23857 40001 23891 40035
rect 24777 40001 24811 40035
rect 47133 40001 47167 40035
rect 47225 40001 47259 40035
rect 14657 39933 14691 39967
rect 14841 39933 14875 39967
rect 17601 39933 17635 39967
rect 19257 39933 19291 39967
rect 22201 39933 22235 39967
rect 23949 39933 23983 39967
rect 24501 39933 24535 39967
rect 24685 39865 24719 39899
rect 23581 39797 23615 39831
rect 24593 39797 24627 39831
rect 47961 39797 47995 39831
rect 13185 39593 13219 39627
rect 24593 39593 24627 39627
rect 25513 39525 25547 39559
rect 21465 39457 21499 39491
rect 22017 39457 22051 39491
rect 23857 39457 23891 39491
rect 46857 39457 46891 39491
rect 48329 39457 48363 39491
rect 13093 39389 13127 39423
rect 21741 39389 21775 39423
rect 22385 39389 22419 39423
rect 22753 39389 22787 39423
rect 23673 39389 23707 39423
rect 23765 39389 23799 39423
rect 23949 39389 23983 39423
rect 24777 39389 24811 39423
rect 25421 39389 25455 39423
rect 25605 39389 25639 39423
rect 24961 39321 24995 39355
rect 48145 39321 48179 39355
rect 23489 39253 23523 39287
rect 47869 39049 47903 39083
rect 20913 38981 20947 39015
rect 24593 38981 24627 39015
rect 24685 38981 24719 39015
rect 1685 38913 1719 38947
rect 14749 38913 14783 38947
rect 14933 38913 14967 38947
rect 16037 38913 16071 38947
rect 16129 38913 16163 38947
rect 18337 38913 18371 38947
rect 20545 38913 20579 38947
rect 22017 38913 22051 38947
rect 22109 38913 22143 38947
rect 22293 38913 22327 38947
rect 23581 38913 23615 38947
rect 24409 38913 24443 38947
rect 24777 38913 24811 38947
rect 47777 38913 47811 38947
rect 15945 38845 15979 38879
rect 16221 38845 16255 38879
rect 18429 38845 18463 38879
rect 20637 38845 20671 38879
rect 20821 38845 20855 38879
rect 23489 38845 23523 38879
rect 23857 38845 23891 38879
rect 23949 38845 23983 38879
rect 1869 38777 1903 38811
rect 22477 38777 22511 38811
rect 15117 38709 15151 38743
rect 15761 38709 15795 38743
rect 17969 38709 18003 38743
rect 23305 38709 23339 38743
rect 24961 38709 24995 38743
rect 13553 38505 13587 38539
rect 16957 38505 16991 38539
rect 18889 38505 18923 38539
rect 22293 38505 22327 38539
rect 23305 38505 23339 38539
rect 25973 38505 26007 38539
rect 15117 38437 15151 38471
rect 6745 38301 6779 38335
rect 12173 38301 12207 38335
rect 14841 38301 14875 38335
rect 15577 38301 15611 38335
rect 17509 38301 17543 38335
rect 22477 38301 22511 38335
rect 23581 38301 23615 38335
rect 24593 38301 24627 38335
rect 24860 38301 24894 38335
rect 47685 38301 47719 38335
rect 12440 38233 12474 38267
rect 15117 38233 15151 38267
rect 15844 38233 15878 38267
rect 17776 38233 17810 38267
rect 22661 38233 22695 38267
rect 23305 38233 23339 38267
rect 6561 38165 6595 38199
rect 14933 38165 14967 38199
rect 23489 38165 23523 38199
rect 6009 37961 6043 37995
rect 12909 37961 12943 37995
rect 13645 37961 13679 37995
rect 14013 37961 14047 37995
rect 14841 37961 14875 37995
rect 15669 37961 15703 37995
rect 18705 37961 18739 37995
rect 24501 37961 24535 37995
rect 6806 37893 6840 37927
rect 15009 37893 15043 37927
rect 15209 37893 15243 37927
rect 16313 37893 16347 37927
rect 17601 37893 17635 37927
rect 18337 37893 18371 37927
rect 18429 37893 18463 37927
rect 4813 37825 4847 37859
rect 5825 37825 5859 37859
rect 6561 37825 6595 37859
rect 8493 37825 8527 37859
rect 13093 37825 13127 37859
rect 15853 37825 15887 37859
rect 15945 37825 15979 37859
rect 17509 37825 17543 37859
rect 17693 37825 17727 37859
rect 18153 37825 18187 37859
rect 18521 37825 18555 37859
rect 19809 37825 19843 37859
rect 20453 37825 20487 37859
rect 23121 37825 23155 37859
rect 23388 37825 23422 37859
rect 47777 37825 47811 37859
rect 14105 37757 14139 37791
rect 14289 37757 14323 37791
rect 16221 37757 16255 37791
rect 19901 37757 19935 37791
rect 4813 37621 4847 37655
rect 7941 37621 7975 37655
rect 8493 37621 8527 37655
rect 15025 37621 15059 37655
rect 19533 37621 19567 37655
rect 20545 37621 20579 37655
rect 20913 37621 20947 37655
rect 47869 37621 47903 37655
rect 6193 37417 6227 37451
rect 6929 37417 6963 37451
rect 7941 37417 7975 37451
rect 18245 37417 18279 37451
rect 20637 37417 20671 37451
rect 6653 37349 6687 37383
rect 15945 37349 15979 37383
rect 27905 37349 27939 37383
rect 1961 37281 1995 37315
rect 4813 37281 4847 37315
rect 13737 37281 13771 37315
rect 15393 37281 15427 37315
rect 18705 37281 18739 37315
rect 20085 37281 20119 37315
rect 28457 37281 28491 37315
rect 48145 37281 48179 37315
rect 4169 37213 4203 37247
rect 7113 37213 7147 37247
rect 7665 37213 7699 37247
rect 9321 37213 9355 37247
rect 12725 37213 12759 37247
rect 13369 37213 13403 37247
rect 13553 37213 13587 37247
rect 14657 37213 14691 37247
rect 14933 37213 14967 37247
rect 15577 37213 15611 37247
rect 18429 37213 18463 37247
rect 18613 37213 18647 37247
rect 19717 37213 19751 37247
rect 19809 37213 19843 37247
rect 20177 37213 20211 37247
rect 22017 37213 22051 37247
rect 27445 37213 27479 37247
rect 28089 37213 28123 37247
rect 28181 37213 28215 37247
rect 46489 37213 46523 37247
rect 48329 37213 48363 37247
rect 1685 37145 1719 37179
rect 5058 37145 5092 37179
rect 14473 37145 14507 37179
rect 14841 37145 14875 37179
rect 15761 37145 15795 37179
rect 21750 37145 21784 37179
rect 27200 37145 27234 37179
rect 28549 37145 28583 37179
rect 4353 37077 4387 37111
rect 8125 37077 8159 37111
rect 9137 37077 9171 37111
rect 12909 37077 12943 37111
rect 15669 37077 15703 37111
rect 19533 37077 19567 37111
rect 26065 37077 26099 37111
rect 15577 36873 15611 36907
rect 20913 36873 20947 36907
rect 22477 36873 22511 36907
rect 25513 36873 25547 36907
rect 8116 36805 8150 36839
rect 13176 36805 13210 36839
rect 15393 36805 15427 36839
rect 20637 36805 20671 36839
rect 22109 36805 22143 36839
rect 24777 36805 24811 36839
rect 4528 36737 4562 36771
rect 7849 36737 7883 36771
rect 12909 36737 12943 36771
rect 15301 36737 15335 36771
rect 15669 36737 15703 36771
rect 19533 36737 19567 36771
rect 20361 36737 20395 36771
rect 20545 36737 20579 36771
rect 20729 36737 20763 36771
rect 22017 36737 22051 36771
rect 22293 36737 22327 36771
rect 24685 36737 24719 36771
rect 24961 36737 24995 36771
rect 25421 36737 25455 36771
rect 25605 36737 25639 36771
rect 27721 36737 27755 36771
rect 27988 36737 28022 36771
rect 4261 36669 4295 36703
rect 15485 36669 15519 36703
rect 19441 36669 19475 36703
rect 19901 36669 19935 36703
rect 14289 36601 14323 36635
rect 5641 36533 5675 36567
rect 9229 36533 9263 36567
rect 24685 36533 24719 36567
rect 29101 36533 29135 36567
rect 47961 36533 47995 36567
rect 4353 36329 4387 36363
rect 5089 36329 5123 36363
rect 5457 36329 5491 36363
rect 6009 36329 6043 36363
rect 9229 36329 9263 36363
rect 17325 36329 17359 36363
rect 21373 36329 21407 36363
rect 23949 36329 23983 36363
rect 26525 36329 26559 36363
rect 26709 36329 26743 36363
rect 27997 36329 28031 36363
rect 9597 36193 9631 36227
rect 21741 36193 21775 36227
rect 46857 36193 46891 36227
rect 48329 36193 48363 36227
rect 4537 36125 4571 36159
rect 5549 36125 5583 36159
rect 6193 36125 6227 36159
rect 8125 36125 8159 36159
rect 9137 36125 9171 36159
rect 10241 36125 10275 36159
rect 17049 36125 17083 36159
rect 21557 36125 21591 36159
rect 23857 36125 23891 36159
rect 24041 36125 24075 36159
rect 24961 36125 24995 36159
rect 25145 36125 25179 36159
rect 25605 36125 25639 36159
rect 25789 36125 25823 36159
rect 27445 36125 27479 36159
rect 27721 36125 27755 36159
rect 27813 36125 27847 36159
rect 8401 36057 8435 36091
rect 24777 36057 24811 36091
rect 25697 36057 25731 36091
rect 26341 36057 26375 36091
rect 27629 36057 27663 36091
rect 48145 36057 48179 36091
rect 10057 35989 10091 36023
rect 26541 35989 26575 36023
rect 5641 35785 5675 35819
rect 14105 35785 14139 35819
rect 21373 35785 21407 35819
rect 24961 35785 24995 35819
rect 47869 35785 47903 35819
rect 9352 35717 9386 35751
rect 27169 35717 27203 35751
rect 5181 35649 5215 35683
rect 9597 35649 9631 35683
rect 14102 35649 14136 35683
rect 14565 35649 14599 35683
rect 18153 35649 18187 35683
rect 21281 35649 21315 35683
rect 22293 35649 22327 35683
rect 23305 35649 23339 35683
rect 24777 35649 24811 35683
rect 25053 35649 25087 35683
rect 25973 35649 26007 35683
rect 26157 35649 26191 35683
rect 26341 35649 26375 35683
rect 26433 35649 26467 35683
rect 27445 35649 27479 35683
rect 32321 35649 32355 35683
rect 32588 35649 32622 35683
rect 35265 35649 35299 35683
rect 35449 35649 35483 35683
rect 47777 35649 47811 35683
rect 18061 35581 18095 35615
rect 23213 35581 23247 35615
rect 27169 35581 27203 35615
rect 17785 35513 17819 35547
rect 23673 35513 23707 35547
rect 5457 35445 5491 35479
rect 8217 35445 8251 35479
rect 13921 35445 13955 35479
rect 14473 35445 14507 35479
rect 22201 35445 22235 35479
rect 24593 35445 24627 35479
rect 27353 35445 27387 35479
rect 33701 35445 33735 35479
rect 35357 35445 35391 35479
rect 5733 35241 5767 35275
rect 21005 35241 21039 35275
rect 22569 35241 22603 35275
rect 25053 35241 25087 35275
rect 25145 35241 25179 35275
rect 25789 35241 25823 35275
rect 26249 35241 26283 35275
rect 27353 35241 27387 35275
rect 33057 35241 33091 35275
rect 17049 35173 17083 35207
rect 24961 35173 24995 35207
rect 28365 35173 28399 35207
rect 8401 35105 8435 35139
rect 15669 35105 15703 35139
rect 17785 35105 17819 35139
rect 20821 35105 20855 35139
rect 26157 35105 26191 35139
rect 27629 35105 27663 35139
rect 28641 35105 28675 35139
rect 33517 35105 33551 35139
rect 36921 35105 36955 35139
rect 4353 35037 4387 35071
rect 8309 35037 8343 35071
rect 17693 35037 17727 35071
rect 17877 35037 17911 35071
rect 17969 35037 18003 35071
rect 20637 35037 20671 35071
rect 21005 35037 21039 35071
rect 23949 35037 23983 35071
rect 24869 35037 24903 35071
rect 25329 35037 25363 35071
rect 25973 35037 26007 35071
rect 26249 35037 26283 35071
rect 27721 35037 27755 35071
rect 28733 35037 28767 35071
rect 29837 35037 29871 35071
rect 31953 35037 31987 35071
rect 32137 35037 32171 35071
rect 32413 35037 32447 35071
rect 32597 35037 32631 35071
rect 33241 35037 33275 35071
rect 33425 35037 33459 35071
rect 35725 35037 35759 35071
rect 36185 35037 36219 35071
rect 36369 35037 36403 35071
rect 38761 35037 38795 35071
rect 38945 35037 38979 35071
rect 39221 35037 39255 35071
rect 4620 34969 4654 35003
rect 15936 34969 15970 35003
rect 21833 34969 21867 35003
rect 23682 34969 23716 35003
rect 24593 34969 24627 35003
rect 30082 34969 30116 35003
rect 35449 34969 35483 35003
rect 35633 34969 35667 35003
rect 37166 34969 37200 35003
rect 7941 34901 7975 34935
rect 17509 34901 17543 34935
rect 20729 34901 20763 34935
rect 21557 34901 21591 34935
rect 31217 34901 31251 34935
rect 35541 34901 35575 34935
rect 36277 34901 36311 34935
rect 38301 34901 38335 34935
rect 39405 34901 39439 34935
rect 1777 34697 1811 34731
rect 4445 34697 4479 34731
rect 5733 34697 5767 34731
rect 9045 34697 9079 34731
rect 16129 34697 16163 34731
rect 16865 34697 16899 34731
rect 20913 34697 20947 34731
rect 22385 34697 22419 34731
rect 23673 34697 23707 34731
rect 24869 34697 24903 34731
rect 27169 34697 27203 34731
rect 29377 34697 29411 34731
rect 33885 34697 33919 34731
rect 36001 34697 36035 34731
rect 36921 34697 36955 34731
rect 37565 34697 37599 34731
rect 23949 34629 23983 34663
rect 24041 34629 24075 34663
rect 24179 34629 24213 34663
rect 34529 34629 34563 34663
rect 35817 34629 35851 34663
rect 38568 34629 38602 34663
rect 1593 34561 1627 34595
rect 4629 34561 4663 34595
rect 5089 34561 5123 34595
rect 5273 34561 5307 34595
rect 5917 34561 5951 34595
rect 7389 34561 7423 34595
rect 8861 34561 8895 34595
rect 9689 34561 9723 34595
rect 14022 34561 14056 34595
rect 14289 34561 14323 34595
rect 14749 34561 14783 34595
rect 15025 34561 15059 34595
rect 16037 34561 16071 34595
rect 16313 34561 16347 34595
rect 17141 34561 17175 34595
rect 17417 34561 17451 34595
rect 18429 34561 18463 34595
rect 18521 34561 18555 34595
rect 18705 34561 18739 34595
rect 20729 34561 20763 34595
rect 22385 34561 22419 34595
rect 23857 34561 23891 34595
rect 24777 34561 24811 34595
rect 27353 34561 27387 34595
rect 27537 34561 27571 34595
rect 29561 34561 29595 34595
rect 30297 34561 30331 34595
rect 30481 34561 30515 34595
rect 30757 34561 30791 34595
rect 30941 34561 30975 34595
rect 33701 34561 33735 34595
rect 33885 34561 33919 34595
rect 34345 34561 34379 34595
rect 35633 34561 35667 34595
rect 36461 34561 36495 34595
rect 36737 34561 36771 34595
rect 37473 34561 37507 34595
rect 37657 34561 37691 34595
rect 7113 34493 7147 34527
rect 7297 34493 7331 34527
rect 17049 34493 17083 34527
rect 17509 34493 17543 34527
rect 22017 34493 22051 34527
rect 22569 34493 22603 34527
rect 24317 34493 24351 34527
rect 29837 34493 29871 34527
rect 36553 34493 36587 34527
rect 38301 34493 38335 34527
rect 16313 34425 16347 34459
rect 34713 34425 34747 34459
rect 5181 34357 5215 34391
rect 7205 34357 7239 34391
rect 9597 34357 9631 34391
rect 12909 34357 12943 34391
rect 18429 34357 18463 34391
rect 27353 34357 27387 34391
rect 29745 34357 29779 34391
rect 39681 34357 39715 34391
rect 14473 34153 14507 34187
rect 18337 34153 18371 34187
rect 19809 34153 19843 34187
rect 20821 34153 20855 34187
rect 21005 34153 21039 34187
rect 27261 34153 27295 34187
rect 27629 34153 27663 34187
rect 36369 34153 36403 34187
rect 37657 34153 37691 34187
rect 35449 34085 35483 34119
rect 9413 34017 9447 34051
rect 15393 34017 15427 34051
rect 19625 34017 19659 34051
rect 32413 34017 32447 34051
rect 36553 34017 36587 34051
rect 38761 34017 38795 34051
rect 39221 34017 39255 34051
rect 4169 33949 4203 33983
rect 4436 33949 4470 33983
rect 7021 33949 7055 33983
rect 7297 33949 7331 33983
rect 8033 33949 8067 33983
rect 9680 33949 9714 33983
rect 12081 33949 12115 33983
rect 13553 33949 13587 33983
rect 14289 33949 14323 33983
rect 14473 33949 14507 33983
rect 17417 33949 17451 33983
rect 17509 33949 17543 33983
rect 17739 33949 17773 33983
rect 17877 33949 17911 33983
rect 18521 33949 18555 33983
rect 18797 33949 18831 33983
rect 19441 33949 19475 33983
rect 19717 33949 19751 33983
rect 19901 33949 19935 33983
rect 26249 33949 26283 33983
rect 27169 33949 27203 33983
rect 27445 33949 27479 33983
rect 30113 33949 30147 33983
rect 30297 33949 30331 33983
rect 30389 33949 30423 33983
rect 35173 33949 35207 33983
rect 35357 33949 35391 33983
rect 35541 33949 35575 33983
rect 35633 33949 35667 33983
rect 36277 33949 36311 33983
rect 37841 33949 37875 33983
rect 38117 33949 38151 33983
rect 38301 33949 38335 33983
rect 38945 33949 38979 33983
rect 39129 33949 39163 33983
rect 7205 33881 7239 33915
rect 15660 33881 15694 33915
rect 17233 33881 17267 33915
rect 17601 33881 17635 33915
rect 21189 33881 21223 33915
rect 26065 33881 26099 33915
rect 32680 33881 32714 33915
rect 5549 33813 5583 33847
rect 6837 33813 6871 33847
rect 7849 33813 7883 33847
rect 10793 33813 10827 33847
rect 12265 33813 12299 33847
rect 13461 33813 13495 33847
rect 16773 33813 16807 33847
rect 18705 33813 18739 33847
rect 20177 33813 20211 33847
rect 20989 33813 21023 33847
rect 25881 33813 25915 33847
rect 29929 33813 29963 33847
rect 33793 33813 33827 33847
rect 35817 33813 35851 33847
rect 36553 33813 36587 33847
rect 4353 33609 4387 33643
rect 5457 33609 5491 33643
rect 6929 33609 6963 33643
rect 9689 33609 9723 33643
rect 19441 33609 19475 33643
rect 21189 33609 21223 33643
rect 28089 33609 28123 33643
rect 30573 33609 30607 33643
rect 32781 33609 32815 33643
rect 7634 33541 7668 33575
rect 10241 33541 10275 33575
rect 12826 33541 12860 33575
rect 17785 33541 17819 33575
rect 17969 33541 18003 33575
rect 25605 33541 25639 33575
rect 25697 33541 25731 33575
rect 27353 33541 27387 33575
rect 4537 33473 4571 33507
rect 4997 33473 5031 33507
rect 6745 33473 6779 33507
rect 7389 33473 7423 33507
rect 9229 33473 9263 33507
rect 10333 33473 10367 33507
rect 13093 33473 13127 33507
rect 17141 33473 17175 33507
rect 17325 33473 17359 33507
rect 18705 33473 18739 33507
rect 18797 33473 18831 33507
rect 18889 33473 18923 33507
rect 19625 33473 19659 33507
rect 19717 33473 19751 33507
rect 20177 33473 20211 33507
rect 20361 33473 20395 33507
rect 21097 33473 21131 33507
rect 21281 33473 21315 33507
rect 24685 33473 24719 33507
rect 25513 33473 25547 33507
rect 25815 33473 25849 33507
rect 25973 33473 26007 33507
rect 26433 33473 26467 33507
rect 26617 33473 26651 33507
rect 27169 33473 27203 33507
rect 27997 33473 28031 33507
rect 28181 33473 28215 33507
rect 29929 33473 29963 33507
rect 30113 33473 30147 33507
rect 30389 33473 30423 33507
rect 32965 33473 32999 33507
rect 35357 33473 35391 33507
rect 46949 33473 46983 33507
rect 19441 33405 19475 33439
rect 23857 33405 23891 33439
rect 35449 33405 35483 33439
rect 20269 33337 20303 33371
rect 26525 33337 26559 33371
rect 34989 33337 35023 33371
rect 5273 33269 5307 33303
rect 8769 33269 8803 33303
rect 9321 33269 9355 33303
rect 11713 33269 11747 33303
rect 17233 33269 17267 33303
rect 18153 33269 18187 33303
rect 25329 33269 25363 33303
rect 27537 33269 27571 33303
rect 47041 33269 47075 33303
rect 7389 33065 7423 33099
rect 8033 33065 8067 33099
rect 20269 33065 20303 33099
rect 26341 33065 26375 33099
rect 27445 33065 27479 33099
rect 31125 33065 31159 33099
rect 33057 33065 33091 33099
rect 40417 33065 40451 33099
rect 5273 32997 5307 33031
rect 7849 32997 7883 33031
rect 10333 32929 10367 32963
rect 12817 32929 12851 32963
rect 17601 32929 17635 32963
rect 20729 32929 20763 32963
rect 21097 32929 21131 32963
rect 22477 32929 22511 32963
rect 22661 32929 22695 32963
rect 24961 32929 24995 32963
rect 29745 32929 29779 32963
rect 31585 32929 31619 32963
rect 33701 32929 33735 32963
rect 46673 32929 46707 32963
rect 3985 32861 4019 32895
rect 6009 32861 6043 32895
rect 6276 32861 6310 32895
rect 8309 32861 8343 32895
rect 10149 32861 10183 32895
rect 12541 32861 12575 32895
rect 13737 32861 13771 32895
rect 20085 32861 20119 32895
rect 20269 32861 20303 32895
rect 20913 32861 20947 32895
rect 21741 32861 21775 32895
rect 21833 32861 21867 32895
rect 22385 32861 22419 32895
rect 23949 32861 23983 32895
rect 25228 32861 25262 32895
rect 27353 32861 27387 32895
rect 27537 32861 27571 32895
rect 30012 32861 30046 32895
rect 31769 32861 31803 32895
rect 33425 32861 33459 32895
rect 35357 32861 35391 32895
rect 35541 32861 35575 32895
rect 38945 32861 38979 32895
rect 39129 32861 39163 32895
rect 40233 32861 40267 32895
rect 40509 32861 40543 32895
rect 45753 32861 45787 32895
rect 46489 32861 46523 32895
rect 5457 32793 5491 32827
rect 12633 32793 12667 32827
rect 18429 32793 18463 32827
rect 48329 32793 48363 32827
rect 9781 32725 9815 32759
rect 10241 32725 10275 32759
rect 12173 32725 12207 32759
rect 13553 32725 13587 32759
rect 21557 32725 21591 32759
rect 22661 32725 22695 32759
rect 23949 32725 23983 32759
rect 31953 32725 31987 32759
rect 33517 32725 33551 32759
rect 35449 32725 35483 32759
rect 38945 32725 38979 32759
rect 40049 32725 40083 32759
rect 45661 32725 45695 32759
rect 1777 32521 1811 32555
rect 6653 32521 6687 32555
rect 10333 32521 10367 32555
rect 10793 32521 10827 32555
rect 12265 32521 12299 32555
rect 14565 32521 14599 32555
rect 15393 32521 15427 32555
rect 15485 32521 15519 32555
rect 18061 32521 18095 32555
rect 24685 32521 24719 32555
rect 26249 32521 26283 32555
rect 28549 32521 28583 32555
rect 33149 32521 33183 32555
rect 33609 32521 33643 32555
rect 34069 32521 34103 32555
rect 40509 32521 40543 32555
rect 9220 32453 9254 32487
rect 13452 32453 13486 32487
rect 33977 32453 34011 32487
rect 36369 32453 36403 32487
rect 45569 32453 45603 32487
rect 47225 32453 47259 32487
rect 1593 32385 1627 32419
rect 3801 32385 3835 32419
rect 6837 32385 6871 32419
rect 10977 32385 11011 32419
rect 13185 32385 13219 32419
rect 17969 32385 18003 32419
rect 18153 32385 18187 32419
rect 18981 32385 19015 32419
rect 20729 32385 20763 32419
rect 21465 32385 21499 32419
rect 22273 32385 22307 32419
rect 24777 32385 24811 32419
rect 25053 32385 25087 32419
rect 26157 32385 26191 32419
rect 26433 32385 26467 32419
rect 27169 32385 27203 32419
rect 27425 32385 27459 32419
rect 31401 32385 31435 32419
rect 32505 32385 32539 32419
rect 32689 32385 32723 32419
rect 33057 32385 33091 32419
rect 35173 32385 35207 32419
rect 35541 32385 35575 32419
rect 35725 32385 35759 32419
rect 36553 32385 36587 32419
rect 38025 32385 38059 32419
rect 38292 32385 38326 32419
rect 39865 32385 39899 32419
rect 40049 32385 40083 32419
rect 40325 32385 40359 32419
rect 44741 32385 44775 32419
rect 47777 32385 47811 32419
rect 3985 32317 4019 32351
rect 4261 32317 4295 32351
rect 8953 32317 8987 32351
rect 11805 32317 11839 32351
rect 15577 32317 15611 32351
rect 19073 32317 19107 32351
rect 20637 32317 20671 32351
rect 21189 32317 21223 32351
rect 22017 32317 22051 32351
rect 26617 32317 26651 32351
rect 31493 32317 31527 32351
rect 32321 32317 32355 32351
rect 34253 32317 34287 32351
rect 35357 32317 35391 32351
rect 35449 32317 35483 32351
rect 45385 32317 45419 32351
rect 12173 32249 12207 32283
rect 21373 32249 21407 32283
rect 31033 32249 31067 32283
rect 15025 32181 15059 32215
rect 19349 32181 19383 32215
rect 20361 32181 20395 32215
rect 20545 32181 20579 32215
rect 21281 32181 21315 32215
rect 23397 32181 23431 32215
rect 34989 32181 35023 32215
rect 36185 32181 36219 32215
rect 39405 32181 39439 32215
rect 44833 32181 44867 32215
rect 4537 31977 4571 32011
rect 9229 31977 9263 32011
rect 11069 31977 11103 32011
rect 14289 31977 14323 32011
rect 19441 31977 19475 32011
rect 21925 31977 21959 32011
rect 36737 31977 36771 32011
rect 38301 31977 38335 32011
rect 38945 31977 38979 32011
rect 41429 31977 41463 32011
rect 6193 31909 6227 31943
rect 14473 31909 14507 31943
rect 23857 31909 23891 31943
rect 31125 31909 31159 31943
rect 7021 31841 7055 31875
rect 10425 31841 10459 31875
rect 15209 31841 15243 31875
rect 17601 31841 17635 31875
rect 20821 31841 20855 31875
rect 22109 31841 22143 31875
rect 22477 31841 22511 31875
rect 22569 31841 22603 31875
rect 31769 31841 31803 31875
rect 31953 31841 31987 31875
rect 35357 31841 35391 31875
rect 37933 31841 37967 31875
rect 40049 31841 40083 31875
rect 46029 31841 46063 31875
rect 47685 31841 47719 31875
rect 4629 31773 4663 31807
rect 5917 31773 5951 31807
rect 7113 31773 7147 31807
rect 9229 31773 9263 31807
rect 10609 31773 10643 31807
rect 14749 31773 14783 31807
rect 22201 31773 22235 31807
rect 23673 31773 23707 31807
rect 24777 31773 24811 31807
rect 25053 31773 25087 31807
rect 25605 31773 25639 31807
rect 30849 31773 30883 31807
rect 30941 31773 30975 31807
rect 31125 31773 31159 31807
rect 31861 31773 31895 31807
rect 32045 31773 32079 31807
rect 35613 31773 35647 31807
rect 37565 31773 37599 31807
rect 37749 31773 37783 31807
rect 37841 31773 37875 31807
rect 38117 31773 38151 31807
rect 39313 31773 39347 31807
rect 40305 31773 40339 31807
rect 45845 31773 45879 31807
rect 10701 31705 10735 31739
rect 15476 31705 15510 31739
rect 17417 31705 17451 31739
rect 17509 31705 17543 31739
rect 20554 31705 20588 31739
rect 39129 31705 39163 31739
rect 6745 31637 6779 31671
rect 16589 31637 16623 31671
rect 17049 31637 17083 31671
rect 25697 31637 25731 31671
rect 31585 31637 31619 31671
rect 13093 31433 13127 31467
rect 13461 31433 13495 31467
rect 20177 31433 20211 31467
rect 24869 31433 24903 31467
rect 25789 31433 25823 31467
rect 35081 31433 35115 31467
rect 36001 31433 36035 31467
rect 44281 31433 44315 31467
rect 5917 31365 5951 31399
rect 6745 31365 6779 31399
rect 15485 31365 15519 31399
rect 16957 31365 16991 31399
rect 19901 31365 19935 31399
rect 35633 31365 35667 31399
rect 6009 31297 6043 31331
rect 6561 31297 6595 31331
rect 9045 31297 9079 31331
rect 10517 31297 10551 31331
rect 12633 31297 12667 31331
rect 18061 31297 18095 31331
rect 19533 31297 19567 31331
rect 19691 31297 19725 31331
rect 19809 31297 19843 31331
rect 19993 31297 20027 31331
rect 24685 31297 24719 31331
rect 24777 31297 24811 31331
rect 25145 31297 25179 31331
rect 25697 31297 25731 31331
rect 25881 31297 25915 31331
rect 28365 31297 28399 31331
rect 28632 31297 28666 31331
rect 30205 31297 30239 31331
rect 30389 31297 30423 31331
rect 31309 31297 31343 31331
rect 31493 31297 31527 31331
rect 33701 31297 33735 31331
rect 33968 31297 34002 31331
rect 35541 31297 35575 31331
rect 35817 31297 35851 31331
rect 37841 31297 37875 31331
rect 39037 31297 39071 31331
rect 39221 31297 39255 31331
rect 43157 31297 43191 31331
rect 44741 31297 44775 31331
rect 8217 31229 8251 31263
rect 13553 31229 13587 31263
rect 13645 31229 13679 31263
rect 17417 31229 17451 31263
rect 37473 31229 37507 31263
rect 37749 31229 37783 31263
rect 42901 31229 42935 31263
rect 15853 31161 15887 31195
rect 17325 31161 17359 31195
rect 9229 31093 9263 31127
rect 10333 31093 10367 31127
rect 12449 31093 12483 31127
rect 15945 31093 15979 31127
rect 17877 31093 17911 31127
rect 25053 31093 25087 31127
rect 25145 31093 25179 31127
rect 29745 31093 29779 31127
rect 30297 31093 30331 31127
rect 31493 31093 31527 31127
rect 39129 31093 39163 31127
rect 44925 31093 44959 31127
rect 13737 30889 13771 30923
rect 15669 30889 15703 30923
rect 28917 30889 28951 30923
rect 36461 30889 36495 30923
rect 42625 30889 42659 30923
rect 46581 30889 46615 30923
rect 6837 30753 6871 30787
rect 12357 30753 12391 30787
rect 30297 30753 30331 30787
rect 43729 30753 43763 30787
rect 45201 30753 45235 30787
rect 6101 30685 6135 30719
rect 8585 30685 8619 30719
rect 9597 30685 9631 30719
rect 9873 30685 9907 30719
rect 10517 30685 10551 30719
rect 10784 30685 10818 30719
rect 15853 30685 15887 30719
rect 17713 30685 17747 30719
rect 17969 30685 18003 30719
rect 25421 30685 25455 30719
rect 25569 30685 25603 30719
rect 25927 30685 25961 30719
rect 29101 30685 29135 30719
rect 37197 30685 37231 30719
rect 37289 30685 37323 30719
rect 37473 30685 37507 30719
rect 42441 30685 42475 30719
rect 44465 30685 44499 30719
rect 44649 30685 44683 30719
rect 45457 30685 45491 30719
rect 12624 30617 12658 30651
rect 25697 30617 25731 30651
rect 25789 30617 25823 30651
rect 36093 30617 36127 30651
rect 36277 30617 36311 30651
rect 43453 30617 43487 30651
rect 8401 30549 8435 30583
rect 11897 30549 11931 30583
rect 16589 30549 16623 30583
rect 26065 30549 26099 30583
rect 29745 30549 29779 30583
rect 30113 30549 30147 30583
rect 30205 30549 30239 30583
rect 43085 30549 43119 30583
rect 43545 30549 43579 30583
rect 44281 30549 44315 30583
rect 11713 30345 11747 30379
rect 12909 30345 12943 30379
rect 29929 30345 29963 30379
rect 40147 30345 40181 30379
rect 44189 30345 44223 30379
rect 9680 30277 9714 30311
rect 17693 30277 17727 30311
rect 40233 30277 40267 30311
rect 44341 30277 44375 30311
rect 44557 30277 44591 30311
rect 6929 30209 6963 30243
rect 9413 30209 9447 30243
rect 12081 30209 12115 30243
rect 13093 30209 13127 30243
rect 15577 30209 15611 30243
rect 22201 30209 22235 30243
rect 23029 30209 23063 30243
rect 23296 30209 23330 30243
rect 25789 30209 25823 30243
rect 27353 30209 27387 30243
rect 29561 30209 29595 30243
rect 32505 30209 32539 30243
rect 34345 30209 34379 30243
rect 34621 30209 34655 30243
rect 34805 30209 34839 30243
rect 35449 30209 35483 30243
rect 35725 30209 35759 30243
rect 35909 30209 35943 30243
rect 38485 30209 38519 30243
rect 38669 30209 38703 30243
rect 39589 30209 39623 30243
rect 40049 30209 40083 30243
rect 40325 30209 40359 30243
rect 40785 30209 40819 30243
rect 40969 30209 41003 30243
rect 43269 30209 43303 30243
rect 43361 30209 43395 30243
rect 43545 30209 43579 30243
rect 47777 30209 47811 30243
rect 6837 30141 6871 30175
rect 12173 30141 12207 30175
rect 12265 30141 12299 30175
rect 18429 30141 18463 30175
rect 22477 30141 22511 30175
rect 25053 30141 25087 30175
rect 27537 30141 27571 30175
rect 29653 30141 29687 30175
rect 32781 30141 32815 30175
rect 38393 30141 38427 30175
rect 39313 30141 39347 30175
rect 39497 30141 39531 30175
rect 10793 30073 10827 30107
rect 32689 30073 32723 30107
rect 40785 30073 40819 30107
rect 6561 30005 6595 30039
rect 15393 30005 15427 30039
rect 22017 30005 22051 30039
rect 22385 30005 22419 30039
rect 24409 30005 24443 30039
rect 27169 30005 27203 30039
rect 32321 30005 32355 30039
rect 34161 30005 34195 30039
rect 35265 30005 35299 30039
rect 38853 30005 38887 30039
rect 39405 30005 39439 30039
rect 43729 30005 43763 30039
rect 44373 30005 44407 30039
rect 47041 30005 47075 30039
rect 47869 30005 47903 30039
rect 44097 29801 44131 29835
rect 13093 29733 13127 29767
rect 17509 29733 17543 29767
rect 23305 29733 23339 29767
rect 27353 29733 27387 29767
rect 32873 29733 32907 29767
rect 33885 29733 33919 29767
rect 42901 29733 42935 29767
rect 6745 29665 6779 29699
rect 7205 29665 7239 29699
rect 10977 29665 11011 29699
rect 12449 29665 12483 29699
rect 18061 29665 18095 29699
rect 25145 29665 25179 29699
rect 25421 29665 25455 29699
rect 25973 29665 26007 29699
rect 35633 29665 35667 29699
rect 37933 29665 37967 29699
rect 40049 29665 40083 29699
rect 43085 29665 43119 29699
rect 43729 29665 43763 29699
rect 46489 29665 46523 29699
rect 46673 29665 46707 29699
rect 10885 29597 10919 29631
rect 14289 29597 14323 29631
rect 15025 29597 15059 29631
rect 19441 29597 19475 29631
rect 19625 29597 19659 29631
rect 19901 29597 19935 29631
rect 21281 29597 21315 29631
rect 23489 29597 23523 29631
rect 25237 29597 25271 29631
rect 25329 29597 25363 29631
rect 26240 29597 26274 29631
rect 29745 29597 29779 29631
rect 29929 29597 29963 29631
rect 30205 29597 30239 29631
rect 31493 29597 31527 29631
rect 34069 29597 34103 29631
rect 34253 29597 34287 29631
rect 34345 29597 34379 29631
rect 37657 29597 37691 29631
rect 37841 29597 37875 29631
rect 38025 29597 38059 29631
rect 38209 29597 38243 29631
rect 38669 29597 38703 29631
rect 38853 29597 38887 29631
rect 39129 29597 39163 29631
rect 42901 29597 42935 29631
rect 43269 29597 43303 29631
rect 43913 29597 43947 29631
rect 6929 29529 6963 29563
rect 12725 29529 12759 29563
rect 15292 29529 15326 29563
rect 17877 29529 17911 29563
rect 17969 29529 18003 29563
rect 21548 29529 21582 29563
rect 31760 29529 31794 29563
rect 34897 29529 34931 29563
rect 37473 29529 37507 29563
rect 40294 29529 40328 29563
rect 43177 29529 43211 29563
rect 48329 29529 48363 29563
rect 10517 29461 10551 29495
rect 12633 29461 12667 29495
rect 14473 29461 14507 29495
rect 16405 29461 16439 29495
rect 20085 29461 20119 29495
rect 22661 29461 22695 29495
rect 24961 29461 24995 29495
rect 30389 29461 30423 29495
rect 39037 29461 39071 29495
rect 41429 29461 41463 29495
rect 6837 29257 6871 29291
rect 15485 29257 15519 29291
rect 29837 29257 29871 29291
rect 8392 29189 8426 29223
rect 14482 29189 14516 29223
rect 19104 29189 19138 29223
rect 40141 29189 40175 29223
rect 40693 29189 40727 29223
rect 43637 29189 43671 29223
rect 5641 29121 5675 29155
rect 6745 29121 6779 29155
rect 15669 29121 15703 29155
rect 15853 29121 15887 29155
rect 19349 29121 19383 29155
rect 19809 29121 19843 29155
rect 20076 29121 20110 29155
rect 22017 29121 22051 29155
rect 22201 29121 22235 29155
rect 22477 29121 22511 29155
rect 22661 29121 22695 29155
rect 24317 29121 24351 29155
rect 25329 29121 25363 29155
rect 25421 29121 25455 29155
rect 25605 29121 25639 29155
rect 27537 29121 27571 29155
rect 28724 29121 28758 29155
rect 30297 29121 30331 29155
rect 30481 29121 30515 29155
rect 30757 29121 30791 29155
rect 32505 29121 32539 29155
rect 32781 29121 32815 29155
rect 32965 29121 32999 29155
rect 33517 29121 33551 29155
rect 33701 29121 33735 29155
rect 34345 29121 34379 29155
rect 34601 29121 34635 29155
rect 36369 29121 36403 29155
rect 36645 29121 36679 29155
rect 36829 29121 36863 29155
rect 38393 29121 38427 29155
rect 38485 29121 38519 29155
rect 38577 29121 38611 29155
rect 38761 29121 38795 29155
rect 40601 29121 40635 29155
rect 40785 29121 40819 29155
rect 43361 29121 43395 29155
rect 43729 29121 43763 29155
rect 47225 29121 47259 29155
rect 8125 29053 8159 29087
rect 14749 29053 14783 29087
rect 24409 29053 24443 29087
rect 27169 29053 27203 29087
rect 27445 29053 27479 29087
rect 28457 29053 28491 29087
rect 30665 29053 30699 29087
rect 33425 29053 33459 29087
rect 33885 29053 33919 29087
rect 43545 29053 43579 29087
rect 5549 28985 5583 29019
rect 13369 28985 13403 29019
rect 23949 28985 23983 29019
rect 25605 28985 25639 29019
rect 36185 28985 36219 29019
rect 38117 28985 38151 29019
rect 39865 28985 39899 29019
rect 43361 28985 43395 29019
rect 47961 28985 47995 29019
rect 9505 28917 9539 28951
rect 17969 28917 18003 28951
rect 21189 28917 21223 28951
rect 32321 28917 32355 28951
rect 35725 28917 35759 28951
rect 39681 28917 39715 28951
rect 46581 28917 46615 28951
rect 47133 28917 47167 28951
rect 8125 28713 8159 28747
rect 13369 28713 13403 28747
rect 16865 28713 16899 28747
rect 19441 28713 19475 28747
rect 19809 28713 19843 28747
rect 22569 28713 22603 28747
rect 23305 28713 23339 28747
rect 24685 28713 24719 28747
rect 31217 28713 31251 28747
rect 36461 28713 36495 28747
rect 38301 28713 38335 28747
rect 39313 28713 39347 28747
rect 12173 28645 12207 28679
rect 40325 28645 40359 28679
rect 5549 28577 5583 28611
rect 6929 28577 6963 28611
rect 7113 28577 7147 28611
rect 9597 28577 9631 28611
rect 9689 28577 9723 28611
rect 12265 28577 12299 28611
rect 14841 28577 14875 28611
rect 17325 28577 17359 28611
rect 17509 28577 17543 28611
rect 23765 28577 23799 28611
rect 23857 28577 23891 28611
rect 30113 28577 30147 28611
rect 32597 28577 32631 28611
rect 35081 28577 35115 28611
rect 42441 28577 42475 28611
rect 42533 28577 42567 28611
rect 46489 28577 46523 28611
rect 46673 28577 46707 28611
rect 48237 28577 48271 28611
rect 8125 28509 8159 28543
rect 12725 28509 12759 28543
rect 14749 28509 14783 28543
rect 17233 28509 17267 28543
rect 18245 28509 18279 28543
rect 18337 28509 18371 28543
rect 18613 28509 18647 28543
rect 19625 28509 19659 28543
rect 19901 28509 19935 28543
rect 20545 28509 20579 28543
rect 20821 28509 20855 28543
rect 21005 28509 21039 28543
rect 22385 28509 22419 28543
rect 22661 28509 22695 28543
rect 24593 28509 24627 28543
rect 24777 28509 24811 28543
rect 29929 28509 29963 28543
rect 30205 28509 30239 28543
rect 33057 28509 33091 28543
rect 33150 28509 33184 28543
rect 33522 28509 33556 28543
rect 37197 28509 37231 28543
rect 37381 28509 37415 28543
rect 38489 28509 38523 28543
rect 38577 28509 38611 28543
rect 38669 28509 38703 28543
rect 39221 28509 39255 28543
rect 39405 28509 39439 28543
rect 40049 28509 40083 28543
rect 40325 28509 40359 28543
rect 42349 28509 42383 28543
rect 42625 28509 42659 28543
rect 43637 28509 43671 28543
rect 43913 28509 43947 28543
rect 11805 28441 11839 28475
rect 13553 28441 13587 28475
rect 13737 28441 13771 28475
rect 18429 28441 18463 28475
rect 32330 28441 32364 28475
rect 33333 28441 33367 28475
rect 33425 28441 33459 28475
rect 35326 28441 35360 28475
rect 40141 28441 40175 28475
rect 9137 28373 9171 28407
rect 9505 28373 9539 28407
rect 12909 28373 12943 28407
rect 14289 28373 14323 28407
rect 14657 28373 14691 28407
rect 18061 28373 18095 28407
rect 20361 28373 20395 28407
rect 22201 28373 22235 28407
rect 23673 28373 23707 28407
rect 29745 28373 29779 28407
rect 33701 28373 33735 28407
rect 37565 28373 37599 28407
rect 42165 28373 42199 28407
rect 43729 28373 43763 28407
rect 44097 28373 44131 28407
rect 11069 28169 11103 28203
rect 18245 28169 18279 28203
rect 20085 28169 20119 28203
rect 23397 28169 23431 28203
rect 30205 28169 30239 28203
rect 34989 28169 35023 28203
rect 42809 28169 42843 28203
rect 43177 28169 43211 28203
rect 44005 28169 44039 28203
rect 12918 28101 12952 28135
rect 29092 28101 29126 28135
rect 38301 28101 38335 28135
rect 38485 28101 38519 28135
rect 40693 28101 40727 28135
rect 6745 28033 6779 28067
rect 9137 28033 9171 28067
rect 10701 28033 10735 28067
rect 13185 28033 13219 28067
rect 16865 28033 16899 28067
rect 17132 28033 17166 28067
rect 20269 28033 20303 28067
rect 20453 28033 20487 28067
rect 22284 28033 22318 28067
rect 25421 28033 25455 28067
rect 25697 28033 25731 28067
rect 27353 28033 27387 28067
rect 34805 28033 34839 28067
rect 39957 28033 39991 28067
rect 41889 28033 41923 28067
rect 43085 28033 43119 28067
rect 43453 28033 43487 28067
rect 43913 28033 43947 28067
rect 44649 28033 44683 28067
rect 44905 28033 44939 28067
rect 47777 28033 47811 28067
rect 6837 27965 6871 27999
rect 7113 27965 7147 27999
rect 10609 27965 10643 27999
rect 20545 27965 20579 27999
rect 22017 27965 22051 27999
rect 27629 27965 27663 27999
rect 28825 27965 28859 27999
rect 34529 27965 34563 27999
rect 41613 27965 41647 27999
rect 42993 27965 43027 27999
rect 43361 27965 43395 27999
rect 25605 27897 25639 27931
rect 27537 27897 27571 27931
rect 34621 27897 34655 27931
rect 8953 27829 8987 27863
rect 11805 27829 11839 27863
rect 25237 27829 25271 27863
rect 27169 27829 27203 27863
rect 46029 27829 46063 27863
rect 47869 27829 47903 27863
rect 12173 27625 12207 27659
rect 17417 27625 17451 27659
rect 22661 27625 22695 27659
rect 29745 27625 29779 27659
rect 38393 27625 38427 27659
rect 38577 27625 38611 27659
rect 44465 27625 44499 27659
rect 7205 27557 7239 27591
rect 8217 27557 8251 27591
rect 10609 27557 10643 27591
rect 26249 27557 26283 27591
rect 36461 27557 36495 27591
rect 40325 27557 40359 27591
rect 7941 27489 7975 27523
rect 10149 27489 10183 27523
rect 12725 27489 12759 27523
rect 14657 27489 14691 27523
rect 17693 27489 17727 27523
rect 17877 27489 17911 27523
rect 24869 27489 24903 27523
rect 33057 27489 33091 27523
rect 41521 27489 41555 27523
rect 46857 27489 46891 27523
rect 48145 27489 48179 27523
rect 48329 27489 48363 27523
rect 5365 27421 5399 27455
rect 5825 27421 5859 27455
rect 7849 27421 7883 27455
rect 10241 27421 10275 27455
rect 14473 27421 14507 27455
rect 14749 27421 14783 27455
rect 17601 27421 17635 27455
rect 17785 27421 17819 27455
rect 22845 27421 22879 27455
rect 23121 27421 23155 27455
rect 23305 27421 23339 27455
rect 26801 27421 26835 27455
rect 29929 27421 29963 27455
rect 30205 27421 30239 27455
rect 30389 27421 30423 27455
rect 32873 27421 32907 27455
rect 33149 27421 33183 27455
rect 36369 27421 36403 27455
rect 36553 27421 36587 27455
rect 38025 27421 38059 27455
rect 40049 27421 40083 27455
rect 41797 27421 41831 27455
rect 43913 27421 43947 27455
rect 44189 27421 44223 27455
rect 44281 27421 44315 27455
rect 5089 27353 5123 27387
rect 6092 27353 6126 27387
rect 12541 27353 12575 27387
rect 25136 27353 25170 27387
rect 27068 27353 27102 27387
rect 40325 27353 40359 27387
rect 44097 27353 44131 27387
rect 12633 27285 12667 27319
rect 14289 27285 14323 27319
rect 28181 27285 28215 27319
rect 32689 27285 32723 27319
rect 38393 27285 38427 27319
rect 40141 27285 40175 27319
rect 42901 27285 42935 27319
rect 6009 27081 6043 27115
rect 6745 27081 6779 27115
rect 7113 27081 7147 27115
rect 17877 27081 17911 27115
rect 21097 27081 21131 27115
rect 25329 27081 25363 27115
rect 27813 27081 27847 27115
rect 33701 27081 33735 27115
rect 37565 27081 37599 27115
rect 32588 27013 32622 27047
rect 36185 27013 36219 27047
rect 40141 27013 40175 27047
rect 5825 26945 5859 26979
rect 7205 26945 7239 26979
rect 8033 26945 8067 26979
rect 9036 26945 9070 26979
rect 14372 26945 14406 26979
rect 17049 26945 17083 26979
rect 18061 26945 18095 26979
rect 18245 26945 18279 26979
rect 25513 26945 25547 26979
rect 25789 26945 25823 26979
rect 25973 26945 26007 26979
rect 27169 26945 27203 26979
rect 27353 26945 27387 26979
rect 27629 26945 27663 26979
rect 35357 26945 35391 26979
rect 37473 26945 37507 26979
rect 37657 26945 37691 26979
rect 39313 26945 39347 26979
rect 40325 26945 40359 26979
rect 41429 26945 41463 26979
rect 41889 26945 41923 26979
rect 43913 26945 43947 26979
rect 44180 26945 44214 26979
rect 46857 26945 46891 26979
rect 47777 26945 47811 26979
rect 7389 26877 7423 26911
rect 8309 26877 8343 26911
rect 8769 26877 8803 26911
rect 14105 26877 14139 26911
rect 17141 26877 17175 26911
rect 17417 26877 17451 26911
rect 21189 26877 21223 26911
rect 21373 26877 21407 26911
rect 32321 26877 32355 26911
rect 36277 26877 36311 26911
rect 36461 26877 36495 26911
rect 39221 26877 39255 26911
rect 39681 26877 39715 26911
rect 42073 26877 42107 26911
rect 10149 26741 10183 26775
rect 15485 26741 15519 26775
rect 20729 26741 20763 26775
rect 35173 26741 35207 26775
rect 35817 26741 35851 26775
rect 40509 26741 40543 26775
rect 45293 26741 45327 26775
rect 46765 26741 46799 26775
rect 47869 26741 47903 26775
rect 9965 26537 9999 26571
rect 14565 26537 14599 26571
rect 18153 26537 18187 26571
rect 23765 26537 23799 26571
rect 26249 26537 26283 26571
rect 33425 26537 33459 26571
rect 36737 26537 36771 26571
rect 38945 26537 38979 26571
rect 44189 26537 44223 26571
rect 20453 26469 20487 26503
rect 37933 26469 37967 26503
rect 40049 26469 40083 26503
rect 9689 26401 9723 26435
rect 17233 26401 17267 26435
rect 17601 26401 17635 26435
rect 21097 26401 21131 26435
rect 24593 26401 24627 26435
rect 32045 26401 32079 26435
rect 37013 26401 37047 26435
rect 37749 26401 37783 26435
rect 38209 26401 38243 26435
rect 46489 26401 46523 26435
rect 46673 26401 46707 26435
rect 47961 26401 47995 26435
rect 9597 26333 9631 26367
rect 12265 26333 12299 26367
rect 14749 26333 14783 26367
rect 15025 26333 15059 26367
rect 15209 26333 15243 26367
rect 17141 26333 17175 26367
rect 18061 26333 18095 26367
rect 18245 26333 18279 26367
rect 19809 26333 19843 26367
rect 20821 26333 20855 26367
rect 23581 26333 23615 26367
rect 23857 26333 23891 26367
rect 24777 26333 24811 26367
rect 25053 26333 25087 26367
rect 25237 26333 25271 26367
rect 25973 26333 26007 26367
rect 34897 26333 34931 26367
rect 37105 26333 37139 26367
rect 39129 26333 39163 26367
rect 39313 26333 39347 26367
rect 39497 26333 39531 26367
rect 41429 26333 41463 26367
rect 44005 26333 44039 26367
rect 32312 26265 32346 26299
rect 35164 26265 35198 26299
rect 39221 26265 39255 26299
rect 41162 26265 41196 26299
rect 12081 26197 12115 26231
rect 16957 26197 16991 26231
rect 19993 26197 20027 26231
rect 20913 26197 20947 26231
rect 23397 26197 23431 26231
rect 36277 26197 36311 26231
rect 7941 25993 7975 26027
rect 21465 25993 21499 26027
rect 24317 25993 24351 26027
rect 33057 25993 33091 26027
rect 35449 25993 35483 26027
rect 35909 25993 35943 26027
rect 40233 25993 40267 26027
rect 43821 25993 43855 26027
rect 11980 25925 12014 25959
rect 18429 25925 18463 25959
rect 20330 25925 20364 25959
rect 23204 25925 23238 25959
rect 6828 25857 6862 25891
rect 17785 25857 17819 25891
rect 18613 25857 18647 25891
rect 18705 25857 18739 25891
rect 19165 25857 19199 25891
rect 22017 25857 22051 25891
rect 22201 25857 22235 25891
rect 22937 25857 22971 25891
rect 25329 25857 25363 25891
rect 26249 25857 26283 25891
rect 26433 25857 26467 25891
rect 30685 25857 30719 25891
rect 32413 25857 32447 25891
rect 32597 25857 32631 25891
rect 32873 25857 32907 25891
rect 33885 25857 33919 25891
rect 35817 25857 35851 25891
rect 38025 25857 38059 25891
rect 38117 25857 38151 25891
rect 38209 25857 38243 25891
rect 38853 25857 38887 25891
rect 39037 25857 39071 25891
rect 39129 25857 39163 25891
rect 39221 25857 39255 25891
rect 40049 25857 40083 25891
rect 40325 25857 40359 25891
rect 44189 25857 44223 25891
rect 6561 25789 6595 25823
rect 11713 25789 11747 25823
rect 20085 25789 20119 25823
rect 25605 25789 25639 25823
rect 30941 25789 30975 25823
rect 34621 25789 34655 25823
rect 36093 25789 36127 25823
rect 39865 25789 39899 25823
rect 44281 25789 44315 25823
rect 44465 25789 44499 25823
rect 46765 25789 46799 25823
rect 47041 25789 47075 25823
rect 47225 25789 47259 25823
rect 18429 25721 18463 25755
rect 19533 25721 19567 25755
rect 22017 25721 22051 25755
rect 39405 25721 39439 25755
rect 2329 25653 2363 25687
rect 13093 25653 13127 25687
rect 17877 25653 17911 25687
rect 19625 25653 19659 25687
rect 26433 25653 26467 25687
rect 29561 25653 29595 25687
rect 38393 25653 38427 25687
rect 47961 25653 47995 25687
rect 6469 25449 6503 25483
rect 7113 25449 7147 25483
rect 11437 25449 11471 25483
rect 18613 25449 18647 25483
rect 21557 25449 21591 25483
rect 24961 25449 24995 25483
rect 28457 25449 28491 25483
rect 31217 25449 31251 25483
rect 32229 25449 32263 25483
rect 43085 25449 43119 25483
rect 43913 25449 43947 25483
rect 44097 25449 44131 25483
rect 45201 25449 45235 25483
rect 45385 25449 45419 25483
rect 18521 25381 18555 25415
rect 21005 25381 21039 25415
rect 42073 25381 42107 25415
rect 3433 25313 3467 25347
rect 9597 25313 9631 25347
rect 9689 25313 9723 25347
rect 12817 25313 12851 25347
rect 17049 25313 17083 25347
rect 20545 25313 20579 25347
rect 23765 25313 23799 25347
rect 31677 25313 31711 25347
rect 33517 25313 33551 25347
rect 43269 25313 43303 25347
rect 46857 25313 46891 25347
rect 48145 25313 48179 25347
rect 48329 25313 48363 25347
rect 1593 25245 1627 25279
rect 6469 25245 6503 25279
rect 7297 25245 7331 25279
rect 8309 25245 8343 25279
rect 9505 25245 9539 25279
rect 12633 25245 12667 25279
rect 15025 25245 15059 25279
rect 15945 25245 15979 25279
rect 16221 25245 16255 25279
rect 16313 25245 16347 25279
rect 17141 25245 17175 25279
rect 18429 25245 18463 25279
rect 18705 25245 18739 25279
rect 18889 25245 18923 25279
rect 20637 25245 20671 25279
rect 21465 25245 21499 25279
rect 21649 25245 21683 25279
rect 23673 25245 23707 25279
rect 25789 25245 25823 25279
rect 26056 25245 26090 25279
rect 28641 25245 28675 25279
rect 30113 25245 30147 25279
rect 30297 25245 30331 25279
rect 30573 25245 30607 25279
rect 30757 25245 30791 25279
rect 31401 25245 31435 25279
rect 31585 25245 31619 25279
rect 32413 25245 32447 25279
rect 32597 25245 32631 25279
rect 32689 25245 32723 25279
rect 33701 25245 33735 25279
rect 33977 25245 34011 25279
rect 34161 25245 34195 25279
rect 40141 25245 40175 25279
rect 42349 25245 42383 25279
rect 43085 25245 43119 25279
rect 43453 25245 43487 25279
rect 3249 25177 3283 25211
rect 8585 25177 8619 25211
rect 11621 25177 11655 25211
rect 11805 25177 11839 25211
rect 16129 25177 16163 25211
rect 25145 25177 25179 25211
rect 25329 25177 25363 25211
rect 40877 25177 40911 25211
rect 42073 25177 42107 25211
rect 43361 25177 43395 25211
rect 44281 25177 44315 25211
rect 45569 25177 45603 25211
rect 9137 25109 9171 25143
rect 12265 25109 12299 25143
rect 12725 25109 12759 25143
rect 14841 25109 14875 25143
rect 16497 25109 16531 25143
rect 17509 25109 17543 25143
rect 18153 25109 18187 25143
rect 23305 25109 23339 25143
rect 27169 25109 27203 25143
rect 42257 25109 42291 25143
rect 44081 25109 44115 25143
rect 45359 25109 45393 25143
rect 9505 24905 9539 24939
rect 15761 24905 15795 24939
rect 17877 24905 17911 24939
rect 23397 24905 23431 24939
rect 27353 24905 27387 24939
rect 32597 24905 32631 24939
rect 41981 24905 42015 24939
rect 45661 24905 45695 24939
rect 10333 24837 10367 24871
rect 14648 24837 14682 24871
rect 25237 24837 25271 24871
rect 2605 24769 2639 24803
rect 7573 24769 7607 24803
rect 8392 24769 8426 24803
rect 10241 24769 10275 24803
rect 11713 24769 11747 24803
rect 11969 24769 12003 24803
rect 13553 24769 13587 24803
rect 13737 24769 13771 24803
rect 16865 24769 16899 24803
rect 17049 24769 17083 24803
rect 17693 24769 17727 24803
rect 17877 24769 17911 24803
rect 18337 24769 18371 24803
rect 18521 24769 18555 24803
rect 19717 24769 19751 24803
rect 22201 24769 22235 24803
rect 23673 24769 23707 24803
rect 25881 24769 25915 24803
rect 26249 24769 26283 24803
rect 27169 24769 27203 24803
rect 27445 24769 27479 24803
rect 30297 24769 30331 24803
rect 30757 24769 30791 24803
rect 30941 24769 30975 24803
rect 31217 24769 31251 24803
rect 31401 24769 31435 24803
rect 32321 24769 32355 24803
rect 32781 24769 32815 24803
rect 33609 24769 33643 24803
rect 33793 24769 33827 24803
rect 34069 24769 34103 24803
rect 39037 24769 39071 24803
rect 41797 24769 41831 24803
rect 42073 24769 42107 24803
rect 43176 24769 43210 24803
rect 44281 24769 44315 24803
rect 44548 24769 44582 24803
rect 46397 24769 46431 24803
rect 46489 24769 46523 24803
rect 47225 24769 47259 24803
rect 48237 24769 48271 24803
rect 2513 24701 2547 24735
rect 7665 24701 7699 24735
rect 8125 24701 8159 24735
rect 10057 24701 10091 24735
rect 14381 24701 14415 24735
rect 17233 24701 17267 24735
rect 19993 24701 20027 24735
rect 23121 24701 23155 24735
rect 23765 24701 23799 24735
rect 38761 24701 38795 24735
rect 41705 24701 41739 24735
rect 43085 24701 43119 24735
rect 43269 24701 43303 24735
rect 43361 24701 43395 24735
rect 27169 24633 27203 24667
rect 29009 24633 29043 24667
rect 48053 24633 48087 24667
rect 10701 24565 10735 24599
rect 13093 24565 13127 24599
rect 13921 24565 13955 24599
rect 18429 24565 18463 24599
rect 19533 24565 19567 24599
rect 19901 24565 19935 24599
rect 22109 24565 22143 24599
rect 34253 24565 34287 24599
rect 38853 24565 38887 24599
rect 39221 24565 39255 24599
rect 41613 24565 41647 24599
rect 43545 24565 43579 24599
rect 11805 24361 11839 24395
rect 13001 24361 13035 24395
rect 16773 24361 16807 24395
rect 19625 24361 19659 24395
rect 27169 24361 27203 24395
rect 38117 24361 38151 24395
rect 42717 24361 42751 24395
rect 43545 24361 43579 24395
rect 9137 24225 9171 24259
rect 12449 24225 12483 24259
rect 12541 24225 12575 24259
rect 16037 24225 16071 24259
rect 17785 24225 17819 24259
rect 17877 24225 17911 24259
rect 21833 24225 21867 24259
rect 22017 24225 22051 24259
rect 22845 24225 22879 24259
rect 26617 24225 26651 24259
rect 29009 24225 29043 24259
rect 32873 24225 32907 24259
rect 43177 24225 43211 24259
rect 44005 24225 44039 24259
rect 48145 24225 48179 24259
rect 8217 24157 8251 24191
rect 11161 24157 11195 24191
rect 11621 24157 11655 24191
rect 14565 24157 14599 24191
rect 14841 24157 14875 24191
rect 15025 24157 15059 24191
rect 15945 24157 15979 24191
rect 16681 24157 16715 24191
rect 16865 24157 16899 24191
rect 19809 24157 19843 24191
rect 20085 24157 20119 24191
rect 20269 24157 20303 24191
rect 25697 24157 25731 24191
rect 26801 24157 26835 24191
rect 28365 24157 28399 24191
rect 28549 24157 28583 24191
rect 28641 24157 28675 24191
rect 28733 24157 28767 24191
rect 30941 24157 30975 24191
rect 31585 24157 31619 24191
rect 36093 24157 36127 24191
rect 39497 24157 39531 24191
rect 41337 24157 41371 24191
rect 43361 24157 43395 24191
rect 44189 24157 44223 24191
rect 46489 24157 46523 24191
rect 6377 24089 6411 24123
rect 8033 24089 8067 24123
rect 9404 24089 9438 24123
rect 12633 24089 12667 24123
rect 15853 24089 15887 24123
rect 17693 24089 17727 24123
rect 30757 24089 30791 24123
rect 31125 24089 31159 24123
rect 31861 24089 31895 24123
rect 33140 24089 33174 24123
rect 36338 24089 36372 24123
rect 39230 24089 39264 24123
rect 41604 24089 41638 24123
rect 46673 24089 46707 24123
rect 10517 24021 10551 24055
rect 10977 24021 11011 24055
rect 14381 24021 14415 24055
rect 15485 24021 15519 24055
rect 17325 24021 17359 24055
rect 25881 24021 25915 24055
rect 26709 24021 26743 24055
rect 34253 24021 34287 24055
rect 37473 24021 37507 24055
rect 44373 24021 44407 24055
rect 6653 23817 6687 23851
rect 8861 23817 8895 23851
rect 9689 23817 9723 23851
rect 10149 23817 10183 23851
rect 15393 23817 15427 23851
rect 20637 23817 20671 23851
rect 22753 23817 22787 23851
rect 23581 23817 23615 23851
rect 24041 23817 24075 23851
rect 26433 23817 26467 23851
rect 27169 23817 27203 23851
rect 28549 23817 28583 23851
rect 36093 23817 36127 23851
rect 38853 23817 38887 23851
rect 44465 23817 44499 23851
rect 47869 23817 47903 23851
rect 26525 23749 26559 23783
rect 29684 23749 29718 23783
rect 6561 23681 6595 23715
rect 9045 23681 9079 23715
rect 10057 23681 10091 23715
rect 14280 23681 14314 23715
rect 19257 23681 19291 23715
rect 19513 23681 19547 23715
rect 22569 23681 22603 23715
rect 22753 23681 22787 23715
rect 23213 23681 23247 23715
rect 23397 23681 23431 23715
rect 24041 23681 24075 23715
rect 24225 23681 24259 23715
rect 27721 23681 27755 23715
rect 30389 23681 30423 23715
rect 31493 23681 31527 23715
rect 33333 23681 33367 23715
rect 33609 23681 33643 23715
rect 33793 23681 33827 23715
rect 34253 23681 34287 23715
rect 34520 23681 34554 23715
rect 36277 23681 36311 23715
rect 36645 23681 36679 23715
rect 36829 23681 36863 23715
rect 39037 23681 39071 23715
rect 39313 23681 39347 23715
rect 39497 23681 39531 23715
rect 40693 23681 40727 23715
rect 44281 23681 44315 23715
rect 47041 23681 47075 23715
rect 47777 23681 47811 23715
rect 10241 23613 10275 23647
rect 14013 23613 14047 23647
rect 27445 23613 27479 23647
rect 29929 23613 29963 23647
rect 36461 23613 36495 23647
rect 36553 23613 36587 23647
rect 30573 23545 30607 23579
rect 27353 23477 27387 23511
rect 31677 23477 31711 23511
rect 33149 23477 33183 23511
rect 35633 23477 35667 23511
rect 40417 23477 40451 23511
rect 14289 23273 14323 23307
rect 26341 23273 26375 23307
rect 31769 23273 31803 23307
rect 33057 23273 33091 23307
rect 34897 23273 34931 23307
rect 37657 23273 37691 23307
rect 42349 23273 42383 23307
rect 42625 23205 42659 23239
rect 12357 23137 12391 23171
rect 14749 23137 14783 23171
rect 22385 23137 22419 23171
rect 22477 23137 22511 23171
rect 24961 23137 24995 23171
rect 27997 23137 28031 23171
rect 33425 23137 33459 23171
rect 33517 23137 33551 23171
rect 35357 23137 35391 23171
rect 42717 23137 42751 23171
rect 12081 23069 12115 23103
rect 14473 23069 14507 23103
rect 14657 23069 14691 23103
rect 19901 23069 19935 23103
rect 24777 23069 24811 23103
rect 25053 23069 25087 23103
rect 27629 23069 27663 23103
rect 28457 23069 28491 23103
rect 28641 23069 28675 23103
rect 30297 23069 30331 23103
rect 30481 23069 30515 23103
rect 30757 23069 30791 23103
rect 33241 23069 33275 23103
rect 35081 23069 35115 23103
rect 35265 23069 35299 23103
rect 36553 23069 36587 23103
rect 36737 23069 36771 23103
rect 37565 23069 37599 23103
rect 37749 23069 37783 23103
rect 42533 23069 42567 23103
rect 42809 23069 42843 23103
rect 19625 23001 19659 23035
rect 26325 23001 26359 23035
rect 26525 23001 26559 23035
rect 27813 23001 27847 23035
rect 28825 23001 28859 23035
rect 31493 23001 31527 23035
rect 11713 22933 11747 22967
rect 12173 22933 12207 22967
rect 22569 22933 22603 22967
rect 22937 22933 22971 22967
rect 24593 22933 24627 22967
rect 26157 22933 26191 22967
rect 30941 22933 30975 22967
rect 36369 22933 36403 22967
rect 11161 22729 11195 22763
rect 11713 22729 11747 22763
rect 23397 22729 23431 22763
rect 27445 22729 27479 22763
rect 12826 22661 12860 22695
rect 20116 22661 20150 22695
rect 20821 22661 20855 22695
rect 24400 22661 24434 22695
rect 26525 22661 26559 22695
rect 28273 22661 28307 22695
rect 29253 22661 29287 22695
rect 29469 22661 29503 22695
rect 30205 22661 30239 22695
rect 33609 22661 33643 22695
rect 42994 22661 43028 22695
rect 43111 22661 43145 22695
rect 2605 22593 2639 22627
rect 10977 22593 11011 22627
rect 16313 22593 16347 22627
rect 16865 22593 16899 22627
rect 17049 22593 17083 22627
rect 21005 22593 21039 22627
rect 21281 22593 21315 22627
rect 22284 22593 22318 22627
rect 24133 22593 24167 22627
rect 26433 22593 26467 22627
rect 27445 22593 27479 22627
rect 28457 22593 28491 22627
rect 30573 22593 30607 22627
rect 31309 22593 31343 22627
rect 31493 22593 31527 22627
rect 31585 22593 31619 22627
rect 33793 22593 33827 22627
rect 36277 22593 36311 22627
rect 36461 22593 36495 22627
rect 37473 22593 37507 22627
rect 37657 22593 37691 22627
rect 38945 22593 38979 22627
rect 39201 22593 39235 22627
rect 41889 22593 41923 22627
rect 42809 22593 42843 22627
rect 42901 22593 42935 22627
rect 43729 22593 43763 22627
rect 43913 22593 43947 22627
rect 13093 22525 13127 22559
rect 15577 22525 15611 22559
rect 20361 22525 20395 22559
rect 22017 22525 22051 22559
rect 36369 22525 36403 22559
rect 41705 22525 41739 22559
rect 43269 22525 43303 22559
rect 42073 22457 42107 22491
rect 44097 22457 44131 22491
rect 2513 22389 2547 22423
rect 17049 22389 17083 22423
rect 18981 22389 19015 22423
rect 21189 22389 21223 22423
rect 25513 22389 25547 22423
rect 28641 22389 28675 22423
rect 29101 22389 29135 22423
rect 29285 22389 29319 22423
rect 31125 22389 31159 22423
rect 33977 22389 34011 22423
rect 37565 22389 37599 22423
rect 40325 22389 40359 22423
rect 42625 22389 42659 22423
rect 47961 22389 47995 22423
rect 14657 22185 14691 22219
rect 22569 22185 22603 22219
rect 23213 22185 23247 22219
rect 24593 22185 24627 22219
rect 26617 22185 26651 22219
rect 27905 22185 27939 22219
rect 32321 22185 32355 22219
rect 37841 22185 37875 22219
rect 39037 22185 39071 22219
rect 41337 22185 41371 22219
rect 44189 22185 44223 22219
rect 44281 22185 44315 22219
rect 11621 22117 11655 22151
rect 43453 22117 43487 22151
rect 3249 22049 3283 22083
rect 11437 22049 11471 22083
rect 11897 22049 11931 22083
rect 16129 22049 16163 22083
rect 20085 22049 20119 22083
rect 22017 22049 22051 22083
rect 23765 22049 23799 22083
rect 36369 22049 36403 22083
rect 36829 22049 36863 22083
rect 37381 22049 37415 22083
rect 43177 22049 43211 22083
rect 44097 22049 44131 22083
rect 46857 22049 46891 22083
rect 48329 22049 48363 22083
rect 3433 21981 3467 22015
rect 14473 21981 14507 22015
rect 14749 21981 14783 22015
rect 18153 21981 18187 22015
rect 18245 21981 18279 22015
rect 18337 21981 18371 22015
rect 18521 21981 18555 22015
rect 19441 21981 19475 22015
rect 19625 21981 19659 22015
rect 19901 21981 19935 22015
rect 22753 21981 22787 22015
rect 24777 21981 24811 22015
rect 25053 21981 25087 22015
rect 25237 21981 25271 22015
rect 26985 21981 27019 22015
rect 27537 21981 27571 22015
rect 27813 21981 27847 22015
rect 29009 21981 29043 22015
rect 29929 21981 29963 22015
rect 30113 21981 30147 22015
rect 30205 21981 30239 22015
rect 30941 21981 30975 22015
rect 31208 21981 31242 22015
rect 32781 21981 32815 22015
rect 35265 21981 35299 22015
rect 35449 21981 35483 22015
rect 36461 21981 36495 22015
rect 37473 21981 37507 22015
rect 38301 21981 38335 22015
rect 38485 21981 38519 22015
rect 39221 21981 39255 22015
rect 39497 21981 39531 22015
rect 40417 21981 40451 22015
rect 42450 21981 42484 22015
rect 42717 21981 42751 22015
rect 44373 21981 44407 22015
rect 1593 21913 1627 21947
rect 16396 21913 16430 21947
rect 21189 21913 21223 21947
rect 29193 21913 29227 21947
rect 33048 21913 33082 21947
rect 35357 21913 35391 21947
rect 38393 21913 38427 21947
rect 40785 21913 40819 21947
rect 48145 21913 48179 21947
rect 14289 21845 14323 21879
rect 17509 21845 17543 21879
rect 17969 21845 18003 21879
rect 23581 21845 23615 21879
rect 23673 21845 23707 21879
rect 26433 21845 26467 21879
rect 26617 21845 26651 21879
rect 28089 21845 28123 21879
rect 29745 21845 29779 21879
rect 34161 21845 34195 21879
rect 36185 21845 36219 21879
rect 39405 21845 39439 21879
rect 43637 21845 43671 21879
rect 22293 21641 22327 21675
rect 26525 21641 26559 21675
rect 33333 21641 33367 21675
rect 33885 21641 33919 21675
rect 37841 21641 37875 21675
rect 42625 21641 42659 21675
rect 45293 21641 45327 21675
rect 47869 21641 47903 21675
rect 13544 21573 13578 21607
rect 16313 21573 16347 21607
rect 23428 21573 23462 21607
rect 24133 21573 24167 21607
rect 25513 21573 25547 21607
rect 27445 21573 27479 21607
rect 27629 21573 27663 21607
rect 28733 21573 28767 21607
rect 31401 21573 31435 21607
rect 2329 21505 2363 21539
rect 13277 21505 13311 21539
rect 16129 21505 16163 21539
rect 17233 21505 17267 21539
rect 17325 21505 17359 21539
rect 17877 21505 17911 21539
rect 18245 21505 18279 21539
rect 23673 21505 23707 21539
rect 24317 21505 24351 21539
rect 24593 21505 24627 21539
rect 26341 21505 26375 21539
rect 29561 21505 29595 21539
rect 29828 21505 29862 21539
rect 31585 21505 31619 21539
rect 31769 21505 31803 21539
rect 32597 21505 32631 21539
rect 32781 21505 32815 21539
rect 32873 21505 32907 21539
rect 33149 21505 33183 21539
rect 33793 21505 33827 21539
rect 33977 21505 34011 21539
rect 35541 21505 35575 21539
rect 36369 21505 36403 21539
rect 36553 21505 36587 21539
rect 37657 21505 37691 21539
rect 37933 21505 37967 21539
rect 42993 21505 43027 21539
rect 44465 21505 44499 21539
rect 45109 21505 45143 21539
rect 46397 21505 46431 21539
rect 47777 21505 47811 21539
rect 15945 21437 15979 21471
rect 16865 21437 16899 21471
rect 17049 21437 17083 21471
rect 17141 21437 17175 21471
rect 18153 21437 18187 21471
rect 25237 21437 25271 21471
rect 32965 21437 32999 21471
rect 35633 21437 35667 21471
rect 42901 21437 42935 21471
rect 44373 21437 44407 21471
rect 14657 21369 14691 21403
rect 18061 21369 18095 21403
rect 27261 21369 27295 21403
rect 28917 21369 28951 21403
rect 30941 21369 30975 21403
rect 35173 21369 35207 21403
rect 44097 21369 44131 21403
rect 17969 21301 18003 21335
rect 24501 21301 24535 21335
rect 27445 21301 27479 21335
rect 36185 21301 36219 21335
rect 37473 21301 37507 21335
rect 42809 21301 42843 21335
rect 46489 21301 46523 21335
rect 47041 21301 47075 21335
rect 14289 21097 14323 21131
rect 19993 21097 20027 21131
rect 23581 21097 23615 21131
rect 25605 21097 25639 21131
rect 26341 21097 26375 21131
rect 27261 21097 27295 21131
rect 30021 21097 30055 21131
rect 35265 21097 35299 21131
rect 36553 21097 36587 21131
rect 36921 21097 36955 21131
rect 17325 21029 17359 21063
rect 28825 21029 28859 21063
rect 43269 20961 43303 20995
rect 46489 20961 46523 20995
rect 46673 20961 46707 20995
rect 48237 20961 48271 20995
rect 2145 20893 2179 20927
rect 14473 20893 14507 20927
rect 14749 20893 14783 20927
rect 14933 20893 14967 20927
rect 16129 20893 16163 20927
rect 16313 20893 16347 20927
rect 16773 20893 16807 20927
rect 16865 20893 16899 20927
rect 17049 20893 17083 20927
rect 17141 20893 17175 20927
rect 19809 20893 19843 20927
rect 20085 20893 20119 20927
rect 22937 20893 22971 20927
rect 23121 20893 23155 20927
rect 23397 20893 23431 20927
rect 26249 20893 26283 20927
rect 27077 20893 27111 20927
rect 27261 20893 27295 20927
rect 27905 20893 27939 20927
rect 28641 20893 28675 20927
rect 30205 20893 30239 20927
rect 30481 20893 30515 20927
rect 30665 20893 30699 20927
rect 35357 20893 35391 20927
rect 36553 20893 36587 20927
rect 36737 20893 36771 20927
rect 25329 20825 25363 20859
rect 43536 20825 43570 20859
rect 16313 20757 16347 20791
rect 19625 20757 19659 20791
rect 27445 20757 27479 20791
rect 28089 20757 28123 20791
rect 34897 20757 34931 20791
rect 44649 20757 44683 20791
rect 29745 20553 29779 20587
rect 33885 20553 33919 20587
rect 43729 20553 43763 20587
rect 15209 20485 15243 20519
rect 17877 20485 17911 20519
rect 34589 20485 34623 20519
rect 34805 20485 34839 20519
rect 2053 20417 2087 20451
rect 12541 20417 12575 20451
rect 12725 20417 12759 20451
rect 14105 20417 14139 20451
rect 15117 20417 15151 20451
rect 15301 20417 15335 20451
rect 15945 20417 15979 20451
rect 16037 20417 16071 20451
rect 16313 20417 16347 20451
rect 17049 20417 17083 20451
rect 17233 20417 17267 20451
rect 17325 20417 17359 20451
rect 18061 20417 18095 20451
rect 18153 20417 18187 20451
rect 19257 20417 19291 20451
rect 19513 20417 19547 20451
rect 22017 20417 22051 20451
rect 27813 20417 27847 20451
rect 29561 20417 29595 20451
rect 33701 20417 33735 20451
rect 33977 20417 34011 20451
rect 35633 20417 35667 20451
rect 36001 20417 36035 20451
rect 39396 20417 39430 20451
rect 41797 20417 41831 20451
rect 44005 20417 44039 20451
rect 44281 20417 44315 20451
rect 46213 20417 46247 20451
rect 2237 20349 2271 20383
rect 2789 20349 2823 20383
rect 12817 20349 12851 20383
rect 16865 20349 16899 20383
rect 17142 20349 17176 20383
rect 39129 20349 39163 20383
rect 41061 20349 41095 20383
rect 41521 20349 41555 20383
rect 43913 20349 43947 20383
rect 44373 20349 44407 20383
rect 27997 20281 28031 20315
rect 40509 20281 40543 20315
rect 12357 20213 12391 20247
rect 14289 20213 14323 20247
rect 15761 20213 15795 20247
rect 16221 20213 16255 20247
rect 17877 20213 17911 20247
rect 20637 20213 20671 20247
rect 22201 20213 22235 20247
rect 33701 20213 33735 20247
rect 34437 20213 34471 20247
rect 34621 20213 34655 20247
rect 36001 20213 36035 20247
rect 36185 20213 36219 20247
rect 46305 20213 46339 20247
rect 46857 20213 46891 20247
rect 2421 20009 2455 20043
rect 15669 20009 15703 20043
rect 17877 20009 17911 20043
rect 19717 20009 19751 20043
rect 29101 20009 29135 20043
rect 35449 20009 35483 20043
rect 44097 20009 44131 20043
rect 33793 19941 33827 19975
rect 39497 19941 39531 19975
rect 29745 19873 29779 19907
rect 31677 19873 31711 19907
rect 33609 19873 33643 19907
rect 40233 19873 40267 19907
rect 41153 19873 41187 19907
rect 41521 19873 41555 19907
rect 44281 19873 44315 19907
rect 44557 19873 44591 19907
rect 46489 19873 46523 19907
rect 46673 19873 46707 19907
rect 48237 19873 48271 19907
rect 2513 19805 2547 19839
rect 11897 19805 11931 19839
rect 14289 19805 14323 19839
rect 16313 19805 16347 19839
rect 17693 19805 17727 19839
rect 17877 19805 17911 19839
rect 19901 19805 19935 19839
rect 20177 19805 20211 19839
rect 20361 19805 20395 19839
rect 21833 19805 21867 19839
rect 22017 19805 22051 19839
rect 22293 19805 22327 19839
rect 25697 19805 25731 19839
rect 25881 19805 25915 19839
rect 26157 19805 26191 19839
rect 28917 19805 28951 19839
rect 29193 19805 29227 19839
rect 29929 19805 29963 19839
rect 30205 19805 30239 19839
rect 30389 19805 30423 19839
rect 33885 19805 33919 19839
rect 35357 19805 35391 19839
rect 35541 19805 35575 19839
rect 39221 19805 39255 19839
rect 39313 19805 39347 19839
rect 39497 19805 39531 19839
rect 40325 19805 40359 19839
rect 40601 19805 40635 19839
rect 40693 19805 40727 19839
rect 41337 19805 41371 19839
rect 41429 19805 41463 19839
rect 41613 19805 41647 19839
rect 44373 19805 44407 19839
rect 44465 19805 44499 19839
rect 12164 19737 12198 19771
rect 14556 19737 14590 19771
rect 17141 19737 17175 19771
rect 31944 19737 31978 19771
rect 13277 19669 13311 19703
rect 22477 19669 22511 19703
rect 26341 19669 26375 19703
rect 28733 19669 28767 19703
rect 33057 19669 33091 19703
rect 33885 19669 33919 19703
rect 40049 19669 40083 19703
rect 12817 19465 12851 19499
rect 14657 19465 14691 19499
rect 15025 19465 15059 19499
rect 16221 19465 16255 19499
rect 25237 19465 25271 19499
rect 27169 19465 27203 19499
rect 29837 19465 29871 19499
rect 32321 19465 32355 19499
rect 34529 19465 34563 19499
rect 39129 19465 39163 19499
rect 44195 19465 44229 19499
rect 15117 19397 15151 19431
rect 16865 19397 16899 19431
rect 20637 19397 20671 19431
rect 21465 19397 21499 19431
rect 26372 19397 26406 19431
rect 28724 19397 28758 19431
rect 32597 19397 32631 19431
rect 32689 19397 32723 19431
rect 39865 19397 39899 19431
rect 44097 19397 44131 19431
rect 44925 19397 44959 19431
rect 13001 19329 13035 19363
rect 13277 19329 13311 19363
rect 13461 19329 13495 19363
rect 16037 19329 16071 19363
rect 17095 19329 17129 19363
rect 17233 19329 17267 19363
rect 17325 19329 17359 19363
rect 17509 19329 17543 19363
rect 19349 19329 19383 19363
rect 19533 19329 19567 19363
rect 22201 19329 22235 19363
rect 22385 19329 22419 19363
rect 23664 19329 23698 19363
rect 26617 19329 26651 19363
rect 27353 19329 27387 19363
rect 27537 19329 27571 19363
rect 28457 19329 28491 19363
rect 30665 19329 30699 19363
rect 30849 19329 30883 19363
rect 32459 19329 32493 19363
rect 32872 19329 32906 19363
rect 32965 19329 32999 19363
rect 33609 19329 33643 19363
rect 34437 19329 34471 19363
rect 34713 19329 34747 19363
rect 38016 19329 38050 19363
rect 39589 19329 39623 19363
rect 39773 19329 39807 19363
rect 39957 19329 39991 19363
rect 40095 19329 40129 19363
rect 40969 19329 41003 19363
rect 41797 19329 41831 19363
rect 43453 19329 43487 19363
rect 43637 19329 43671 19363
rect 44281 19329 44315 19363
rect 44373 19329 44407 19363
rect 44833 19329 44867 19363
rect 45017 19329 45051 19363
rect 47225 19329 47259 19363
rect 15209 19261 15243 19295
rect 15853 19261 15887 19295
rect 19257 19261 19291 19295
rect 22477 19261 22511 19295
rect 23397 19261 23431 19295
rect 27629 19261 27663 19295
rect 30941 19261 30975 19295
rect 33701 19261 33735 19295
rect 37749 19261 37783 19295
rect 40233 19261 40267 19295
rect 40693 19261 40727 19295
rect 41981 19261 42015 19295
rect 19717 19125 19751 19159
rect 22017 19125 22051 19159
rect 24777 19125 24811 19159
rect 30481 19125 30515 19159
rect 33977 19125 34011 19159
rect 34897 19125 34931 19159
rect 40785 19125 40819 19159
rect 41153 19125 41187 19159
rect 41613 19125 41647 19159
rect 43637 19125 43671 19159
rect 47133 19125 47167 19159
rect 47777 19125 47811 19159
rect 25237 18921 25271 18955
rect 31585 18921 31619 18955
rect 39405 18921 39439 18955
rect 40785 18921 40819 18955
rect 41245 18921 41279 18955
rect 42165 18921 42199 18955
rect 28641 18853 28675 18887
rect 35541 18853 35575 18887
rect 41613 18853 41647 18887
rect 22845 18785 22879 18819
rect 27813 18785 27847 18819
rect 35081 18785 35115 18819
rect 45845 18785 45879 18819
rect 46489 18785 46523 18819
rect 46673 18785 46707 18819
rect 48237 18785 48271 18819
rect 2053 18717 2087 18751
rect 15485 18717 15519 18751
rect 15669 18717 15703 18751
rect 17049 18717 17083 18751
rect 17325 18717 17359 18751
rect 19441 18717 19475 18751
rect 19708 18717 19742 18751
rect 22578 18717 22612 18751
rect 24593 18717 24627 18751
rect 24686 18717 24720 18751
rect 25099 18717 25133 18751
rect 28457 18717 28491 18751
rect 28733 18717 28767 18751
rect 30205 18717 30239 18751
rect 32781 18717 32815 18751
rect 35173 18717 35207 18751
rect 36369 18717 36403 18751
rect 36553 18717 36587 18751
rect 38393 18717 38427 18751
rect 39313 18717 39347 18751
rect 39497 18717 39531 18751
rect 40417 18717 40451 18751
rect 41245 18717 41279 18751
rect 41429 18717 41463 18751
rect 42073 18717 42107 18751
rect 42257 18717 42291 18751
rect 43545 18717 43579 18751
rect 43729 18717 43763 18751
rect 44189 18717 44223 18751
rect 45385 18717 45419 18751
rect 45477 18717 45511 18751
rect 15577 18649 15611 18683
rect 17233 18649 17267 18683
rect 23857 18649 23891 18683
rect 24041 18649 24075 18683
rect 24869 18649 24903 18683
rect 24961 18649 24995 18683
rect 27568 18649 27602 18683
rect 28273 18649 28307 18683
rect 30472 18649 30506 18683
rect 32045 18649 32079 18683
rect 37657 18649 37691 18683
rect 40601 18649 40635 18683
rect 44373 18649 44407 18683
rect 44557 18649 44591 18683
rect 45569 18649 45603 18683
rect 45707 18649 45741 18683
rect 16865 18581 16899 18615
rect 20821 18581 20855 18615
rect 21465 18581 21499 18615
rect 23673 18581 23707 18615
rect 26433 18581 26467 18615
rect 36553 18581 36587 18615
rect 43637 18581 43671 18615
rect 45201 18581 45235 18615
rect 19993 18377 20027 18411
rect 23949 18377 23983 18411
rect 27813 18377 27847 18411
rect 30941 18377 30975 18411
rect 36921 18377 36955 18411
rect 40417 18377 40451 18411
rect 43729 18377 43763 18411
rect 46029 18377 46063 18411
rect 18245 18309 18279 18343
rect 23581 18309 23615 18343
rect 23781 18309 23815 18343
rect 34897 18309 34931 18343
rect 35725 18309 35759 18343
rect 36553 18309 36587 18343
rect 36645 18309 36679 18343
rect 40049 18309 40083 18343
rect 40233 18309 40267 18343
rect 44097 18309 44131 18343
rect 44916 18309 44950 18343
rect 2053 18241 2087 18275
rect 12357 18241 12391 18275
rect 13093 18241 13127 18275
rect 13277 18241 13311 18275
rect 13553 18241 13587 18275
rect 13737 18241 13771 18275
rect 16129 18241 16163 18275
rect 16313 18241 16347 18275
rect 17969 18241 18003 18275
rect 18153 18241 18187 18275
rect 18337 18241 18371 18275
rect 20177 18241 20211 18275
rect 20453 18241 20487 18275
rect 20637 18241 20671 18275
rect 24409 18241 24443 18275
rect 24593 18241 24627 18275
rect 27169 18241 27203 18275
rect 27353 18241 27387 18275
rect 27629 18241 27663 18275
rect 30297 18241 30331 18275
rect 30481 18241 30515 18275
rect 30757 18241 30791 18275
rect 33793 18241 33827 18275
rect 33977 18241 34011 18275
rect 34529 18241 34563 18275
rect 34621 18241 34655 18275
rect 34713 18241 34747 18275
rect 36369 18241 36403 18275
rect 36737 18241 36771 18275
rect 38586 18241 38620 18275
rect 38853 18241 38887 18275
rect 41153 18241 41187 18275
rect 43913 18241 43947 18275
rect 44189 18241 44223 18275
rect 2237 18173 2271 18207
rect 2789 18173 2823 18207
rect 12173 18173 12207 18207
rect 12633 18173 12667 18207
rect 44649 18173 44683 18207
rect 35357 18105 35391 18139
rect 37473 18105 37507 18139
rect 12541 18037 12575 18071
rect 16221 18037 16255 18071
rect 18521 18037 18555 18071
rect 23765 18037 23799 18071
rect 24501 18037 24535 18071
rect 33977 18037 34011 18071
rect 35725 18037 35759 18071
rect 35909 18037 35943 18071
rect 41337 18037 41371 18071
rect 47961 18037 47995 18071
rect 2329 17833 2363 17867
rect 11437 17833 11471 17867
rect 13645 17833 13679 17867
rect 15485 17833 15519 17867
rect 16221 17833 16255 17867
rect 17141 17833 17175 17867
rect 19533 17833 19567 17867
rect 23305 17833 23339 17867
rect 28825 17833 28859 17867
rect 31861 17833 31895 17867
rect 35265 17833 35299 17867
rect 36645 17833 36679 17867
rect 40049 17833 40083 17867
rect 43913 17833 43947 17867
rect 45385 17833 45419 17867
rect 36277 17765 36311 17799
rect 43821 17765 43855 17799
rect 11345 17697 11379 17731
rect 18521 17697 18555 17731
rect 23029 17697 23063 17731
rect 28733 17697 28767 17731
rect 31401 17697 31435 17731
rect 33241 17697 33275 17731
rect 44005 17697 44039 17731
rect 46857 17697 46891 17731
rect 48329 17697 48363 17731
rect 2421 17629 2455 17663
rect 11621 17629 11655 17663
rect 12265 17629 12299 17663
rect 14473 17629 14507 17663
rect 14749 17629 14783 17663
rect 14933 17629 14967 17663
rect 15393 17629 15427 17663
rect 15577 17629 15611 17663
rect 16405 17629 16439 17663
rect 16681 17629 16715 17663
rect 19441 17629 19475 17663
rect 19717 17629 19751 17663
rect 20361 17629 20395 17663
rect 22937 17629 22971 17663
rect 23765 17629 23799 17663
rect 23949 17629 23983 17663
rect 29009 17629 29043 17663
rect 29745 17629 29779 17663
rect 29929 17629 29963 17663
rect 30205 17629 30239 17663
rect 30389 17629 30423 17663
rect 31125 17629 31159 17663
rect 31309 17629 31343 17663
rect 34897 17629 34931 17663
rect 35081 17629 35115 17663
rect 36185 17629 36219 17663
rect 36461 17629 36495 17663
rect 40233 17629 40267 17663
rect 40509 17629 40543 17663
rect 41337 17629 41371 17663
rect 43729 17629 43763 17663
rect 44121 17629 44155 17663
rect 45201 17629 45235 17663
rect 45477 17629 45511 17663
rect 12532 17561 12566 17595
rect 14289 17561 14323 17595
rect 18276 17561 18310 17595
rect 19901 17561 19935 17595
rect 20606 17561 20640 17595
rect 23857 17561 23891 17595
rect 30941 17561 30975 17595
rect 32974 17561 33008 17595
rect 40969 17561 41003 17595
rect 41245 17561 41279 17595
rect 45293 17561 45327 17595
rect 48145 17561 48179 17595
rect 11805 17493 11839 17527
rect 16589 17493 16623 17527
rect 21741 17493 21775 17527
rect 29193 17493 29227 17527
rect 40417 17493 40451 17527
rect 41153 17493 41187 17527
rect 41521 17493 41555 17527
rect 43453 17493 43487 17527
rect 13277 17289 13311 17323
rect 15117 17289 15151 17323
rect 16957 17289 16991 17323
rect 18153 17289 18187 17323
rect 18521 17289 18555 17323
rect 20821 17289 20855 17323
rect 30113 17289 30147 17323
rect 32689 17289 32723 17323
rect 34989 17289 35023 17323
rect 44281 17289 44315 17323
rect 47869 17289 47903 17323
rect 14933 17221 14967 17255
rect 15945 17221 15979 17255
rect 16129 17221 16163 17255
rect 29000 17221 29034 17255
rect 32781 17221 32815 17255
rect 11897 17153 11931 17187
rect 12153 17153 12187 17187
rect 14749 17153 14783 17187
rect 16865 17153 16899 17187
rect 18061 17153 18095 17187
rect 18337 17153 18371 17187
rect 21005 17153 21039 17187
rect 21281 17153 21315 17187
rect 21465 17153 21499 17187
rect 23121 17153 23155 17187
rect 28733 17153 28767 17187
rect 34897 17153 34931 17187
rect 35081 17153 35115 17187
rect 41061 17153 41095 17187
rect 41337 17153 41371 17187
rect 42625 17153 42659 17187
rect 43085 17153 43119 17187
rect 44465 17153 44499 17187
rect 44557 17153 44591 17187
rect 47777 17153 47811 17187
rect 2053 17085 2087 17119
rect 2237 17085 2271 17119
rect 2881 17085 2915 17119
rect 17233 17085 17267 17119
rect 23397 17085 23431 17119
rect 42901 17085 42935 17119
rect 44281 17085 44315 17119
rect 17141 17017 17175 17051
rect 41245 17017 41279 17051
rect 42993 17017 43027 17051
rect 16313 16949 16347 16983
rect 17325 16949 17359 16983
rect 17601 16949 17635 16983
rect 23213 16949 23247 16983
rect 23305 16949 23339 16983
rect 40877 16949 40911 16983
rect 42763 16949 42797 16983
rect 2145 16745 2179 16779
rect 16037 16745 16071 16779
rect 23121 16745 23155 16779
rect 30389 16745 30423 16779
rect 43453 16745 43487 16779
rect 45293 16745 45327 16779
rect 16865 16677 16899 16711
rect 16497 16609 16531 16643
rect 20821 16609 20855 16643
rect 37565 16609 37599 16643
rect 38117 16609 38151 16643
rect 40693 16609 40727 16643
rect 42993 16609 43027 16643
rect 46121 16609 46155 16643
rect 2881 16541 2915 16575
rect 2973 16541 3007 16575
rect 14749 16541 14783 16575
rect 14933 16541 14967 16575
rect 15669 16541 15703 16575
rect 16681 16541 16715 16575
rect 21465 16541 21499 16575
rect 21649 16541 21683 16575
rect 21833 16541 21867 16575
rect 23489 16541 23523 16575
rect 25237 16541 25271 16575
rect 25421 16541 25455 16575
rect 25605 16541 25639 16575
rect 29745 16541 29779 16575
rect 29929 16541 29963 16575
rect 30205 16541 30239 16575
rect 36093 16541 36127 16575
rect 36277 16541 36311 16575
rect 40233 16541 40267 16575
rect 40325 16541 40359 16575
rect 41889 16541 41923 16575
rect 42073 16541 42107 16575
rect 42165 16541 42199 16575
rect 42257 16541 42291 16575
rect 43085 16541 43119 16575
rect 43269 16541 43303 16575
rect 45201 16541 45235 16575
rect 45385 16541 45419 16575
rect 15853 16473 15887 16507
rect 20554 16473 20588 16507
rect 21557 16473 21591 16507
rect 23305 16473 23339 16507
rect 25329 16473 25363 16507
rect 36737 16473 36771 16507
rect 38384 16473 38418 16507
rect 40601 16473 40635 16507
rect 46388 16473 46422 16507
rect 14841 16405 14875 16439
rect 19441 16405 19475 16439
rect 21281 16405 21315 16439
rect 25053 16405 25087 16439
rect 36277 16405 36311 16439
rect 39497 16405 39531 16439
rect 40049 16405 40083 16439
rect 42533 16405 42567 16439
rect 47501 16405 47535 16439
rect 20269 16201 20303 16235
rect 20637 16201 20671 16235
rect 24501 16201 24535 16235
rect 37565 16201 37599 16235
rect 41337 16201 41371 16235
rect 45661 16201 45695 16235
rect 46673 16201 46707 16235
rect 30941 16133 30975 16167
rect 31769 16133 31803 16167
rect 46305 16133 46339 16167
rect 14565 16065 14599 16099
rect 14657 16065 14691 16099
rect 14841 16065 14875 16099
rect 15945 16065 15979 16099
rect 16129 16065 16163 16099
rect 16865 16065 16899 16099
rect 17049 16065 17083 16099
rect 20453 16065 20487 16099
rect 20729 16065 20763 16099
rect 22937 16065 22971 16099
rect 23213 16065 23247 16099
rect 23305 16065 23339 16099
rect 23489 16065 23523 16099
rect 24133 16065 24167 16099
rect 24961 16065 24995 16099
rect 25053 16065 25087 16099
rect 25237 16065 25271 16099
rect 26341 16065 26375 16099
rect 27169 16065 27203 16099
rect 27353 16065 27387 16099
rect 27629 16065 27663 16099
rect 27813 16065 27847 16099
rect 28365 16065 28399 16099
rect 28632 16065 28666 16099
rect 32321 16065 32355 16099
rect 32577 16065 32611 16099
rect 34161 16065 34195 16099
rect 34417 16065 34451 16099
rect 36001 16065 36035 16099
rect 36185 16065 36219 16099
rect 37473 16065 37507 16099
rect 37749 16065 37783 16099
rect 40049 16065 40083 16099
rect 41153 16065 41187 16099
rect 44281 16065 44315 16099
rect 45293 16065 45327 16099
rect 46121 16065 46155 16099
rect 46397 16065 46431 16099
rect 46489 16065 46523 16099
rect 15853 15997 15887 16031
rect 23121 15997 23155 16031
rect 24041 15997 24075 16031
rect 26525 15997 26559 16031
rect 26617 15997 26651 16031
rect 39957 15997 39991 16031
rect 40877 15997 40911 16031
rect 44373 15997 44407 16031
rect 45385 15997 45419 16031
rect 15025 15929 15059 15963
rect 16313 15929 16347 15963
rect 37749 15929 37783 15963
rect 16957 15861 16991 15895
rect 22753 15861 22787 15895
rect 25421 15861 25455 15895
rect 26157 15861 26191 15895
rect 29745 15861 29779 15895
rect 33701 15861 33735 15895
rect 35541 15861 35575 15895
rect 36369 15861 36403 15895
rect 40417 15861 40451 15895
rect 40969 15861 41003 15895
rect 44649 15861 44683 15895
rect 14657 15657 14691 15691
rect 21465 15657 21499 15691
rect 23305 15657 23339 15691
rect 23673 15657 23707 15691
rect 24593 15657 24627 15691
rect 27445 15657 27479 15691
rect 28733 15657 28767 15691
rect 29101 15657 29135 15691
rect 31309 15657 31343 15691
rect 33609 15657 33643 15691
rect 35633 15657 35667 15691
rect 44005 15657 44039 15691
rect 44189 15657 44223 15691
rect 45477 15657 45511 15691
rect 40325 15589 40359 15623
rect 13645 15521 13679 15555
rect 15025 15521 15059 15555
rect 15761 15521 15795 15555
rect 18337 15521 18371 15555
rect 21005 15521 21039 15555
rect 29193 15521 29227 15555
rect 34069 15521 34103 15555
rect 36369 15521 36403 15555
rect 36461 15521 36495 15555
rect 37565 15521 37599 15555
rect 37841 15521 37875 15555
rect 43545 15521 43579 15555
rect 4721 15453 4755 15487
rect 13553 15453 13587 15487
rect 13737 15453 13771 15487
rect 14565 15453 14599 15487
rect 15669 15453 15703 15487
rect 18061 15453 18095 15487
rect 18245 15453 18279 15487
rect 20453 15453 20487 15487
rect 20821 15453 20855 15487
rect 21465 15453 21499 15487
rect 21649 15453 21683 15487
rect 23765 15453 23799 15487
rect 24593 15453 24627 15487
rect 24777 15453 24811 15487
rect 25237 15453 25271 15487
rect 25421 15453 25455 15487
rect 26065 15453 26099 15487
rect 28917 15453 28951 15487
rect 30389 15453 30423 15487
rect 30665 15453 30699 15487
rect 30849 15453 30883 15487
rect 31493 15453 31527 15487
rect 31677 15453 31711 15487
rect 31769 15453 31803 15487
rect 32413 15453 32447 15487
rect 33793 15453 33827 15487
rect 33977 15453 34011 15487
rect 34161 15453 34195 15487
rect 34345 15453 34379 15487
rect 35541 15453 35575 15487
rect 35725 15453 35759 15487
rect 37473 15453 37507 15487
rect 38301 15453 38335 15487
rect 38485 15453 38519 15487
rect 40049 15453 40083 15487
rect 40325 15453 40359 15487
rect 42533 15453 42567 15487
rect 42717 15453 42751 15487
rect 43269 15453 43303 15487
rect 43361 15453 43395 15487
rect 45201 15453 45235 15487
rect 45293 15453 45327 15487
rect 47685 15453 47719 15487
rect 25329 15385 25363 15419
rect 26310 15385 26344 15419
rect 30205 15385 30239 15419
rect 32229 15385 32263 15419
rect 38393 15385 38427 15419
rect 42349 15385 42383 15419
rect 44173 15385 44207 15419
rect 44373 15385 44407 15419
rect 45477 15385 45511 15419
rect 16037 15317 16071 15351
rect 17877 15317 17911 15351
rect 20821 15317 20855 15351
rect 32597 15317 32631 15351
rect 36185 15317 36219 15351
rect 36829 15317 36863 15351
rect 40141 15317 40175 15351
rect 43545 15317 43579 15351
rect 14289 15113 14323 15147
rect 19993 15113 20027 15147
rect 20745 15113 20779 15147
rect 20913 15113 20947 15147
rect 30113 15113 30147 15147
rect 31217 15113 31251 15147
rect 37841 15113 37875 15147
rect 4169 15045 4203 15079
rect 17776 15045 17810 15079
rect 20545 15045 20579 15079
rect 24308 15045 24342 15079
rect 6009 14977 6043 15011
rect 14197 14977 14231 15011
rect 14381 14977 14415 15011
rect 17509 14977 17543 15011
rect 19901 14977 19935 15011
rect 20085 14977 20119 15011
rect 26157 14977 26191 15011
rect 26341 14977 26375 15011
rect 28733 14977 28767 15011
rect 29000 14977 29034 15011
rect 30573 14977 30607 15011
rect 30757 14977 30791 15011
rect 31033 14977 31067 15011
rect 32321 14977 32355 15011
rect 32588 14977 32622 15011
rect 35449 14977 35483 15011
rect 36645 14977 36679 15011
rect 36829 14977 36863 15011
rect 37473 14977 37507 15011
rect 40325 14977 40359 15011
rect 41521 14977 41555 15011
rect 42901 14977 42935 15011
rect 44005 14977 44039 15011
rect 44833 14977 44867 15011
rect 45017 14977 45051 15011
rect 47777 14977 47811 15011
rect 5825 14909 5859 14943
rect 24041 14909 24075 14943
rect 26433 14909 26467 14943
rect 35541 14909 35575 14943
rect 36737 14909 36771 14943
rect 37565 14909 37599 14943
rect 40417 14909 40451 14943
rect 41429 14909 41463 14943
rect 42993 14909 43027 14943
rect 43269 14909 43303 14943
rect 43913 14909 43947 14943
rect 44281 14909 44315 14943
rect 44373 14909 44407 14943
rect 25421 14841 25455 14875
rect 33701 14841 33735 14875
rect 41153 14841 41187 14875
rect 45201 14841 45235 14875
rect 2329 14773 2363 14807
rect 18889 14773 18923 14807
rect 20729 14773 20763 14807
rect 25973 14773 26007 14807
rect 35173 14773 35207 14807
rect 37473 14773 37507 14807
rect 40601 14773 40635 14807
rect 43729 14773 43763 14807
rect 47869 14773 47903 14807
rect 5089 14569 5123 14603
rect 18153 14569 18187 14603
rect 20177 14569 20211 14603
rect 21281 14569 21315 14603
rect 31309 14569 31343 14603
rect 32597 14569 32631 14603
rect 33977 14569 34011 14603
rect 35081 14569 35115 14603
rect 35449 14569 35483 14603
rect 41613 14569 41647 14603
rect 44649 14569 44683 14603
rect 30941 14501 30975 14535
rect 36461 14501 36495 14535
rect 3433 14433 3467 14467
rect 14841 14433 14875 14467
rect 15025 14433 15059 14467
rect 16589 14433 16623 14467
rect 16773 14433 16807 14467
rect 30389 14433 30423 14467
rect 32965 14433 32999 14467
rect 36645 14433 36679 14467
rect 46857 14433 46891 14467
rect 48145 14433 48179 14467
rect 48329 14433 48363 14467
rect 1593 14365 1627 14399
rect 5181 14365 5215 14399
rect 13737 14365 13771 14399
rect 18337 14365 18371 14399
rect 18613 14365 18647 14399
rect 18797 14365 18831 14399
rect 19993 14365 20027 14399
rect 21097 14365 21131 14399
rect 21373 14365 21407 14399
rect 26626 14365 26660 14399
rect 26893 14365 26927 14399
rect 29745 14365 29779 14399
rect 29929 14365 29963 14399
rect 30205 14365 30239 14399
rect 30849 14365 30883 14399
rect 31125 14365 31159 14399
rect 32781 14365 32815 14399
rect 33057 14365 33091 14399
rect 33149 14365 33183 14399
rect 33333 14365 33367 14399
rect 33793 14365 33827 14399
rect 33977 14365 34011 14399
rect 34989 14365 35023 14399
rect 36369 14365 36403 14399
rect 40233 14365 40267 14399
rect 43269 14365 43303 14399
rect 3249 14297 3283 14331
rect 14749 14297 14783 14331
rect 19809 14297 19843 14331
rect 40500 14297 40534 14331
rect 43536 14297 43570 14331
rect 13553 14229 13587 14263
rect 14381 14229 14415 14263
rect 16129 14229 16163 14263
rect 16497 14229 16531 14263
rect 20913 14229 20947 14263
rect 25513 14229 25547 14263
rect 36645 14229 36679 14263
rect 2421 14025 2455 14059
rect 14565 14025 14599 14059
rect 19533 14025 19567 14059
rect 25789 14025 25823 14059
rect 33241 14025 33275 14059
rect 40509 14025 40543 14059
rect 34161 13957 34195 13991
rect 35909 13957 35943 13991
rect 40877 13957 40911 13991
rect 2513 13889 2547 13923
rect 13185 13889 13219 13923
rect 13452 13889 13486 13923
rect 19441 13889 19475 13923
rect 19625 13889 19659 13923
rect 20352 13889 20386 13923
rect 23397 13889 23431 13923
rect 23581 13889 23615 13923
rect 25973 13889 26007 13923
rect 26249 13889 26283 13923
rect 26433 13889 26467 13923
rect 30021 13889 30055 13923
rect 30205 13889 30239 13923
rect 33057 13889 33091 13923
rect 33241 13889 33275 13923
rect 33793 13889 33827 13923
rect 40693 13889 40727 13923
rect 40785 13889 40819 13923
rect 41061 13889 41095 13923
rect 20085 13821 20119 13855
rect 23673 13821 23707 13855
rect 29929 13821 29963 13855
rect 47961 13821 47995 13855
rect 36185 13753 36219 13787
rect 21465 13685 21499 13719
rect 23213 13685 23247 13719
rect 30389 13685 30423 13719
rect 36369 13685 36403 13719
rect 21005 13481 21039 13515
rect 27353 13481 27387 13515
rect 28549 13481 28583 13515
rect 32689 13481 32723 13515
rect 36277 13481 36311 13515
rect 20177 13413 20211 13447
rect 22661 13345 22695 13379
rect 31309 13345 31343 13379
rect 33517 13345 33551 13379
rect 36369 13345 36403 13379
rect 37657 13345 37691 13379
rect 37749 13345 37783 13379
rect 46857 13345 46891 13379
rect 48329 13345 48363 13379
rect 16221 13277 16255 13311
rect 18245 13277 18279 13311
rect 18521 13277 18555 13311
rect 18705 13277 18739 13311
rect 19901 13277 19935 13311
rect 19993 13277 20027 13311
rect 20177 13277 20211 13311
rect 21189 13277 21223 13311
rect 21465 13277 21499 13311
rect 21649 13277 21683 13311
rect 22928 13277 22962 13311
rect 26065 13277 26099 13311
rect 26249 13277 26283 13311
rect 26525 13277 26559 13311
rect 27169 13277 27203 13311
rect 28365 13277 28399 13311
rect 28641 13277 28675 13311
rect 29929 13277 29963 13311
rect 30113 13277 30147 13311
rect 30389 13277 30423 13311
rect 30573 13277 30607 13311
rect 33333 13277 33367 13311
rect 33609 13277 33643 13311
rect 36001 13277 36035 13311
rect 37565 13277 37599 13311
rect 37841 13277 37875 13311
rect 16488 13209 16522 13243
rect 31576 13209 31610 13243
rect 33149 13209 33183 13243
rect 36461 13209 36495 13243
rect 48145 13209 48179 13243
rect 17601 13141 17635 13175
rect 18061 13141 18095 13175
rect 24041 13141 24075 13175
rect 26709 13141 26743 13175
rect 28181 13141 28215 13175
rect 36093 13141 36127 13175
rect 37381 13141 37415 13175
rect 17049 12937 17083 12971
rect 20453 12937 20487 12971
rect 23305 12937 23339 12971
rect 25237 12937 25271 12971
rect 33609 12937 33643 12971
rect 35541 12937 35575 12971
rect 36737 12937 36771 12971
rect 47869 12937 47903 12971
rect 30288 12869 30322 12903
rect 33425 12869 33459 12903
rect 38770 12869 38804 12903
rect 17233 12801 17267 12835
rect 23489 12801 23523 12835
rect 23765 12801 23799 12835
rect 23949 12801 23983 12835
rect 26350 12801 26384 12835
rect 26617 12801 26651 12835
rect 27721 12801 27755 12835
rect 27988 12801 28022 12835
rect 30021 12801 30055 12835
rect 33241 12801 33275 12835
rect 34897 12801 34931 12835
rect 35081 12801 35115 12835
rect 35725 12801 35759 12835
rect 35909 12801 35943 12835
rect 36369 12801 36403 12835
rect 39037 12801 39071 12835
rect 46397 12801 46431 12835
rect 47777 12801 47811 12835
rect 17509 12733 17543 12767
rect 20545 12733 20579 12767
rect 20637 12733 20671 12767
rect 36461 12733 36495 12767
rect 17417 12665 17451 12699
rect 20085 12597 20119 12631
rect 29101 12597 29135 12631
rect 31401 12597 31435 12631
rect 35081 12597 35115 12631
rect 35909 12597 35943 12631
rect 36369 12597 36403 12631
rect 37657 12597 37691 12631
rect 46489 12597 46523 12631
rect 47041 12597 47075 12631
rect 26157 12393 26191 12427
rect 26525 12393 26559 12427
rect 28457 12393 28491 12427
rect 30205 12393 30239 12427
rect 34989 12393 35023 12427
rect 38025 12393 38059 12427
rect 20269 12325 20303 12359
rect 17417 12257 17451 12291
rect 19993 12257 20027 12291
rect 23581 12257 23615 12291
rect 26617 12257 26651 12291
rect 33977 12257 34011 12291
rect 35909 12257 35943 12291
rect 36185 12257 36219 12291
rect 46489 12257 46523 12291
rect 46673 12257 46707 12291
rect 48237 12257 48271 12291
rect 2421 12189 2455 12223
rect 17233 12189 17267 12223
rect 18061 12189 18095 12223
rect 18245 12189 18279 12223
rect 18705 12189 18739 12223
rect 18889 12189 18923 12223
rect 19901 12189 19935 12223
rect 23397 12189 23431 12223
rect 25421 12189 25455 12223
rect 26341 12189 26375 12223
rect 28641 12189 28675 12223
rect 28917 12189 28951 12223
rect 29101 12189 29135 12223
rect 30389 12189 30423 12223
rect 30665 12189 30699 12223
rect 30849 12189 30883 12223
rect 34897 12189 34931 12223
rect 35173 12189 35207 12223
rect 35265 12189 35299 12223
rect 36093 12189 36127 12223
rect 36277 12189 36311 12223
rect 36369 12189 36403 12223
rect 37473 12189 37507 12223
rect 37657 12189 37691 12223
rect 37841 12189 37875 12223
rect 23489 12121 23523 12155
rect 33793 12121 33827 12155
rect 37749 12121 37783 12155
rect 2329 12053 2363 12087
rect 16865 12053 16899 12087
rect 17325 12053 17359 12087
rect 18245 12053 18279 12087
rect 18797 12053 18831 12087
rect 23029 12053 23063 12087
rect 25605 12053 25639 12087
rect 33425 12053 33459 12087
rect 33885 12053 33919 12087
rect 35449 12053 35483 12087
rect 19993 11849 20027 11883
rect 21281 11849 21315 11883
rect 22293 11849 22327 11883
rect 22385 11849 22419 11883
rect 25329 11849 25363 11883
rect 28733 11849 28767 11883
rect 34897 11849 34931 11883
rect 36461 11849 36495 11883
rect 37565 11849 37599 11883
rect 2237 11781 2271 11815
rect 18981 11781 19015 11815
rect 20177 11781 20211 11815
rect 22017 11781 22051 11815
rect 35357 11781 35391 11815
rect 17049 11713 17083 11747
rect 19901 11713 19935 11747
rect 21189 11713 21223 11747
rect 21465 11713 21499 11747
rect 22201 11713 22235 11747
rect 22569 11713 22603 11747
rect 28549 11713 28583 11747
rect 30665 11713 30699 11747
rect 30849 11713 30883 11747
rect 31125 11713 31159 11747
rect 31309 11713 31343 11747
rect 32505 11713 32539 11747
rect 32689 11713 32723 11747
rect 33517 11713 33551 11747
rect 34713 11713 34747 11747
rect 35541 11713 35575 11747
rect 35633 11713 35667 11747
rect 36093 11713 36127 11747
rect 36277 11713 36311 11747
rect 37473 11713 37507 11747
rect 37657 11713 37691 11747
rect 2053 11645 2087 11679
rect 2789 11645 2823 11679
rect 19441 11645 19475 11679
rect 25421 11645 25455 11679
rect 25513 11645 25547 11679
rect 32781 11645 32815 11679
rect 34529 11645 34563 11679
rect 19257 11577 19291 11611
rect 20177 11577 20211 11611
rect 35357 11577 35391 11611
rect 16865 11509 16899 11543
rect 21465 11509 21499 11543
rect 24961 11509 24995 11543
rect 32321 11509 32355 11543
rect 33333 11509 33367 11543
rect 36093 11509 36127 11543
rect 2053 11305 2087 11339
rect 17325 11305 17359 11339
rect 22937 11305 22971 11339
rect 26525 11305 26559 11339
rect 33057 11305 33091 11339
rect 35081 11305 35115 11339
rect 35633 11305 35667 11339
rect 37105 11305 37139 11339
rect 18153 11237 18187 11271
rect 22477 11169 22511 11203
rect 25145 11169 25179 11203
rect 26433 11169 26467 11203
rect 15945 11101 15979 11135
rect 17969 11101 18003 11135
rect 18245 11101 18279 11135
rect 19717 11101 19751 11135
rect 22569 11101 22603 11135
rect 24961 11101 24995 11135
rect 26709 11101 26743 11135
rect 28549 11101 28583 11135
rect 28733 11101 28767 11135
rect 29009 11101 29043 11135
rect 29745 11101 29779 11135
rect 31677 11101 31711 11135
rect 31944 11101 31978 11135
rect 34897 11101 34931 11135
rect 35081 11101 35115 11135
rect 35541 11101 35575 11135
rect 35725 11101 35759 11135
rect 36369 11101 36403 11135
rect 36553 11101 36587 11135
rect 37013 11101 37047 11135
rect 37197 11101 37231 11135
rect 16212 11033 16246 11067
rect 26893 11033 26927 11067
rect 29990 11033 30024 11067
rect 36185 11033 36219 11067
rect 17785 10965 17819 10999
rect 19533 10965 19567 10999
rect 24593 10965 24627 10999
rect 25053 10965 25087 10999
rect 29193 10965 29227 10999
rect 31125 10965 31159 10999
rect 22661 10761 22695 10795
rect 24593 10761 24627 10795
rect 29561 10761 29595 10795
rect 34529 10761 34563 10795
rect 17592 10693 17626 10727
rect 19432 10693 19466 10727
rect 22293 10693 22327 10727
rect 23949 10693 23983 10727
rect 2973 10625 3007 10659
rect 17325 10625 17359 10659
rect 19165 10625 19199 10659
rect 21281 10625 21315 10659
rect 21465 10625 21499 10659
rect 22017 10625 22051 10659
rect 22110 10625 22144 10659
rect 22385 10625 22419 10659
rect 22523 10625 22557 10659
rect 23397 10625 23431 10659
rect 23857 10625 23891 10659
rect 24041 10625 24075 10659
rect 25706 10625 25740 10659
rect 25973 10625 26007 10659
rect 28282 10625 28316 10659
rect 28549 10625 28583 10659
rect 29745 10625 29779 10659
rect 30021 10625 30055 10659
rect 33149 10625 33183 10659
rect 33416 10625 33450 10659
rect 23121 10557 23155 10591
rect 29929 10557 29963 10591
rect 23305 10489 23339 10523
rect 2329 10421 2363 10455
rect 2881 10421 2915 10455
rect 18705 10421 18739 10455
rect 20545 10421 20579 10455
rect 21373 10421 21407 10455
rect 23213 10421 23247 10455
rect 27169 10421 27203 10455
rect 18245 10217 18279 10251
rect 19901 10217 19935 10251
rect 21649 10217 21683 10251
rect 21833 10217 21867 10251
rect 26249 10217 26283 10251
rect 23857 10149 23891 10183
rect 24869 10149 24903 10183
rect 1593 10081 1627 10115
rect 3249 10081 3283 10115
rect 3433 10081 3467 10115
rect 20545 10081 20579 10115
rect 23397 10081 23431 10115
rect 18429 10013 18463 10047
rect 18705 10013 18739 10047
rect 18889 10013 18923 10047
rect 20361 10013 20395 10047
rect 22845 10013 22879 10047
rect 23489 10013 23523 10047
rect 24685 10013 24719 10047
rect 26433 10013 26467 10047
rect 26709 10013 26743 10047
rect 26893 10013 26927 10047
rect 20269 9945 20303 9979
rect 21465 9945 21499 9979
rect 22661 9945 22695 9979
rect 21675 9877 21709 9911
rect 22477 9877 22511 9911
rect 22201 9673 22235 9707
rect 23857 9673 23891 9707
rect 21097 9605 21131 9639
rect 21281 9605 21315 9639
rect 21465 9537 21499 9571
rect 22017 9537 22051 9571
rect 22201 9537 22235 9571
rect 23029 9537 23063 9571
rect 23213 9537 23247 9571
rect 23673 9537 23707 9571
rect 23857 9537 23891 9571
rect 2053 9469 2087 9503
rect 2237 9469 2271 9503
rect 2973 9469 3007 9503
rect 23121 9469 23155 9503
rect 2145 9129 2179 9163
rect 2881 9129 2915 9163
rect 47961 9129 47995 9163
rect 2973 8925 3007 8959
rect 48237 8857 48271 8891
rect 48329 8449 48363 8483
rect 48053 8381 48087 8415
rect 3433 7837 3467 7871
rect 1593 7769 1627 7803
rect 3249 7769 3283 7803
rect 2881 7497 2915 7531
rect 2329 7361 2363 7395
rect 2789 7361 2823 7395
rect 3433 7157 3467 7191
rect 43269 7157 43303 7191
rect 1593 6817 1627 6851
rect 3433 6817 3467 6851
rect 32321 6817 32355 6851
rect 42809 6817 42843 6851
rect 44649 6817 44683 6851
rect 31401 6749 31435 6783
rect 31861 6749 31895 6783
rect 46213 6749 46247 6783
rect 47041 6749 47075 6783
rect 47685 6749 47719 6783
rect 48145 6749 48179 6783
rect 3249 6681 3283 6715
rect 32045 6681 32079 6715
rect 42993 6681 43027 6715
rect 46949 6613 46983 6647
rect 47593 6613 47627 6647
rect 2421 6409 2455 6443
rect 32413 6409 32447 6443
rect 43085 6409 43119 6443
rect 2513 6273 2547 6307
rect 32505 6273 32539 6307
rect 42993 6273 43027 6307
rect 46397 6273 46431 6307
rect 47225 6273 47259 6307
rect 47777 6273 47811 6307
rect 1869 6069 1903 6103
rect 3157 6069 3191 6103
rect 46489 6069 46523 6103
rect 47133 6069 47167 6103
rect 47869 6069 47903 6103
rect 3433 5729 3467 5763
rect 46121 5729 46155 5763
rect 46305 5729 46339 5763
rect 47133 5729 47167 5763
rect 4169 5661 4203 5695
rect 45661 5661 45695 5695
rect 1593 5593 1627 5627
rect 3249 5593 3283 5627
rect 4077 5593 4111 5627
rect 45569 5525 45603 5559
rect 47041 5253 47075 5287
rect 4629 5185 4663 5219
rect 2789 5117 2823 5151
rect 3801 5117 3835 5151
rect 3985 5117 4019 5151
rect 46765 5117 46799 5151
rect 47225 5117 47259 5151
rect 4537 4981 4571 5015
rect 44741 4981 44775 5015
rect 47961 4981 47995 5015
rect 2513 4777 2547 4811
rect 3065 4777 3099 4811
rect 1777 4709 1811 4743
rect 46857 4641 46891 4675
rect 48145 4641 48179 4675
rect 48329 4641 48363 4675
rect 1593 4573 1627 4607
rect 2973 4573 3007 4607
rect 4169 4573 4203 4607
rect 4629 4573 4663 4607
rect 5457 4573 5491 4607
rect 39037 4573 39071 4607
rect 43085 4573 43119 4607
rect 43913 4573 43947 4607
rect 44557 4573 44591 4607
rect 45201 4573 45235 4607
rect 46029 4573 46063 4607
rect 4077 4437 4111 4471
rect 5365 4437 5399 4471
rect 43177 4437 43211 4471
rect 45293 4437 45327 4471
rect 1685 4165 1719 4199
rect 44281 4165 44315 4199
rect 4077 4097 4111 4131
rect 5825 4097 5859 4131
rect 6653 4097 6687 4131
rect 7573 4097 7607 4131
rect 10517 4097 10551 4131
rect 12541 4097 12575 4131
rect 13185 4097 13219 4131
rect 18613 4097 18647 4131
rect 26157 4097 26191 4131
rect 27169 4097 27203 4131
rect 38393 4097 38427 4131
rect 39037 4097 39071 4131
rect 41521 4097 41555 4131
rect 46765 4097 46799 4131
rect 47777 4097 47811 4131
rect 39221 4029 39255 4063
rect 40509 4029 40543 4063
rect 44005 4029 44039 4063
rect 44465 4029 44499 4063
rect 45753 4029 45787 4063
rect 46581 4029 46615 4063
rect 1961 3961 1995 3995
rect 18705 3961 18739 3995
rect 3065 3893 3099 3927
rect 4169 3893 4203 3927
rect 4997 3893 5031 3927
rect 5917 3893 5951 3927
rect 6745 3893 6779 3927
rect 7665 3893 7699 3927
rect 10609 3893 10643 3927
rect 12449 3893 12483 3927
rect 13277 3893 13311 3927
rect 20085 3893 20119 3927
rect 25329 3893 25363 3927
rect 26065 3893 26099 3927
rect 27261 3893 27295 3927
rect 38485 3893 38519 3927
rect 41429 3893 41463 3927
rect 38209 3621 38243 3655
rect 44189 3621 44223 3655
rect 3249 3553 3283 3587
rect 3433 3553 3467 3587
rect 6101 3553 6135 3587
rect 6469 3553 6503 3587
rect 10701 3553 10735 3587
rect 10977 3553 11011 3587
rect 25973 3553 26007 3587
rect 26433 3553 26467 3587
rect 40785 3553 40819 3587
rect 41245 3553 41279 3587
rect 45201 3553 45235 3587
rect 45385 3553 45419 3587
rect 45661 3553 45695 3587
rect 1593 3485 1627 3519
rect 4169 3485 4203 3519
rect 4813 3485 4847 3519
rect 5457 3485 5491 3519
rect 5917 3485 5951 3519
rect 8217 3485 8251 3519
rect 10517 3485 10551 3519
rect 13185 3485 13219 3519
rect 16957 3485 16991 3519
rect 17601 3485 17635 3519
rect 18889 3485 18923 3519
rect 19441 3485 19475 3519
rect 20085 3485 20119 3519
rect 25329 3485 25363 3519
rect 25789 3485 25823 3519
rect 28089 3485 28123 3519
rect 38117 3485 38151 3519
rect 38761 3485 38795 3519
rect 40601 3485 40635 3519
rect 43085 3485 43119 3519
rect 48329 3485 48363 3519
rect 20361 3417 20395 3451
rect 44005 3417 44039 3451
rect 4721 3349 4755 3383
rect 17509 3349 17543 3383
rect 19533 3349 19567 3383
rect 42993 3349 43027 3383
rect 48145 3349 48179 3383
rect 47869 3145 47903 3179
rect 3525 3077 3559 3111
rect 4353 3077 4387 3111
rect 7665 3077 7699 3111
rect 13369 3077 13403 3111
rect 17049 3077 17083 3111
rect 19809 3077 19843 3111
rect 27353 3077 27387 3111
rect 38945 3077 38979 3111
rect 42809 3077 42843 3111
rect 45109 3077 45143 3111
rect 3709 3009 3743 3043
rect 7481 3009 7515 3043
rect 10517 3009 10551 3043
rect 11713 3009 11747 3043
rect 13185 3009 13219 3043
rect 16865 3009 16899 3043
rect 24777 3009 24811 3043
rect 27169 3009 27203 3043
rect 38761 3009 38795 3043
rect 41061 3009 41095 3043
rect 44925 3009 44959 3043
rect 47777 3009 47811 3043
rect 3249 2941 3283 2975
rect 4169 2941 4203 2975
rect 5181 2941 5215 2975
rect 7941 2941 7975 2975
rect 13645 2941 13679 2975
rect 17417 2941 17451 2975
rect 19625 2941 19659 2975
rect 20637 2941 20671 2975
rect 24961 2941 24995 2975
rect 25789 2941 25823 2975
rect 27721 2941 27755 2975
rect 39313 2941 39347 2975
rect 41889 2941 41923 2975
rect 42625 2941 42659 2975
rect 43085 2941 43119 2975
rect 46765 2941 46799 2975
rect 11897 2873 11931 2907
rect 6653 2805 6687 2839
rect 12449 2805 12483 2839
rect 14473 2601 14507 2635
rect 25421 2601 25455 2635
rect 29929 2601 29963 2635
rect 1593 2465 1627 2499
rect 3433 2465 3467 2499
rect 4077 2465 4111 2499
rect 4537 2465 4571 2499
rect 6653 2465 6687 2499
rect 6837 2465 6871 2499
rect 7113 2465 7147 2499
rect 11897 2465 11931 2499
rect 12909 2465 12943 2499
rect 19441 2465 19475 2499
rect 19901 2465 19935 2499
rect 44097 2465 44131 2499
rect 44649 2465 44683 2499
rect 46765 2465 46799 2499
rect 14289 2397 14323 2431
rect 25513 2397 25547 2431
rect 47225 2397 47259 2431
rect 47777 2397 47811 2431
rect 3249 2329 3283 2363
rect 4261 2329 4295 2363
rect 12081 2329 12115 2363
rect 19625 2329 19659 2363
rect 29837 2329 29871 2363
rect 38945 2329 38979 2363
rect 44465 2329 44499 2363
rect 47041 2329 47075 2363
rect 38853 2261 38887 2295
<< metal1 >>
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 7190 47240 7196 47252
rect 2700 47212 7196 47240
rect 2700 47045 2728 47212
rect 7190 47200 7196 47212
rect 7248 47200 7254 47252
rect 4798 47132 4804 47184
rect 4856 47172 4862 47184
rect 6549 47175 6607 47181
rect 6549 47172 6561 47175
rect 4856 47144 6561 47172
rect 4856 47132 4862 47144
rect 6549 47141 6561 47144
rect 6595 47141 6607 47175
rect 6549 47135 6607 47141
rect 8294 47132 8300 47184
rect 8352 47172 8358 47184
rect 9125 47175 9183 47181
rect 9125 47172 9137 47175
rect 8352 47144 9137 47172
rect 8352 47132 8358 47144
rect 9125 47141 9137 47144
rect 9171 47141 9183 47175
rect 9125 47135 9183 47141
rect 17402 47132 17408 47184
rect 17460 47172 17466 47184
rect 17681 47175 17739 47181
rect 17681 47172 17693 47175
rect 17460 47144 17693 47172
rect 17460 47132 17466 47144
rect 17681 47141 17693 47144
rect 17727 47141 17739 47175
rect 17681 47135 17739 47141
rect 19613 47175 19671 47181
rect 19613 47141 19625 47175
rect 19659 47172 19671 47175
rect 20438 47172 20444 47184
rect 19659 47144 20444 47172
rect 19659 47141 19671 47144
rect 19613 47135 19671 47141
rect 20438 47132 20444 47144
rect 20496 47132 20502 47184
rect 24670 47132 24676 47184
rect 24728 47172 24734 47184
rect 24765 47175 24823 47181
rect 24765 47172 24777 47175
rect 24728 47144 24777 47172
rect 24728 47132 24734 47144
rect 24765 47141 24777 47144
rect 24811 47141 24823 47175
rect 24765 47135 24823 47141
rect 42797 47175 42855 47181
rect 42797 47141 42809 47175
rect 42843 47172 42855 47175
rect 43622 47172 43628 47184
rect 42843 47144 43628 47172
rect 42843 47141 42855 47144
rect 42797 47135 42855 47141
rect 43622 47132 43628 47144
rect 43680 47132 43686 47184
rect 4982 47104 4988 47116
rect 3436 47076 4988 47104
rect 3436 47045 3464 47076
rect 4982 47064 4988 47076
rect 5040 47064 5046 47116
rect 5077 47107 5135 47113
rect 5077 47073 5089 47107
rect 5123 47104 5135 47107
rect 5994 47104 6000 47116
rect 5123 47076 6000 47104
rect 5123 47073 5135 47076
rect 5077 47067 5135 47073
rect 5994 47064 6000 47076
rect 6052 47064 6058 47116
rect 14182 47064 14188 47116
rect 14240 47104 14246 47116
rect 14737 47107 14795 47113
rect 14737 47104 14749 47107
rect 14240 47076 14749 47104
rect 14240 47064 14246 47076
rect 14737 47073 14749 47076
rect 14783 47073 14795 47107
rect 14737 47067 14795 47073
rect 38289 47107 38347 47113
rect 38289 47073 38301 47107
rect 38335 47104 38347 47107
rect 39758 47104 39764 47116
rect 38335 47076 39764 47104
rect 38335 47073 38347 47076
rect 38289 47067 38347 47073
rect 39758 47064 39764 47076
rect 39816 47064 39822 47116
rect 46750 47104 46756 47116
rect 46711 47076 46756 47104
rect 46750 47064 46756 47076
rect 46808 47064 46814 47116
rect 2685 47039 2743 47045
rect 2685 47005 2697 47039
rect 2731 47005 2743 47039
rect 2685 46999 2743 47005
rect 3421 47039 3479 47045
rect 3421 47005 3433 47039
rect 3467 47005 3479 47039
rect 3421 46999 3479 47005
rect 4522 46996 4528 47048
rect 4580 47036 4586 47048
rect 5537 47039 5595 47045
rect 5537 47036 5549 47039
rect 4580 47008 5549 47036
rect 4580 46996 4586 47008
rect 5537 47005 5549 47008
rect 5583 47005 5595 47039
rect 5537 46999 5595 47005
rect 9030 46996 9036 47048
rect 9088 47036 9094 47048
rect 9309 47039 9367 47045
rect 9309 47036 9321 47039
rect 9088 47008 9321 47036
rect 9088 46996 9094 47008
rect 9309 47005 9321 47008
rect 9355 47005 9367 47039
rect 12434 47036 12440 47048
rect 12395 47008 12440 47036
rect 9309 46999 9367 47005
rect 12434 46996 12440 47008
rect 12492 46996 12498 47048
rect 13725 47039 13783 47045
rect 13725 47005 13737 47039
rect 13771 47036 13783 47039
rect 14277 47039 14335 47045
rect 14277 47036 14289 47039
rect 13771 47008 14289 47036
rect 13771 47005 13783 47008
rect 13725 46999 13783 47005
rect 14277 47005 14289 47008
rect 14323 47005 14335 47039
rect 17494 47036 17500 47048
rect 17455 47008 17500 47036
rect 14277 46999 14335 47005
rect 17494 46996 17500 47008
rect 17552 46996 17558 47048
rect 19334 46996 19340 47048
rect 19392 47036 19398 47048
rect 19429 47039 19487 47045
rect 19429 47036 19441 47039
rect 19392 47008 19441 47036
rect 19392 46996 19398 47008
rect 19429 47005 19441 47008
rect 19475 47005 19487 47039
rect 19429 46999 19487 47005
rect 22462 46996 22468 47048
rect 22520 47036 22526 47048
rect 22557 47039 22615 47045
rect 22557 47036 22569 47039
rect 22520 47008 22569 47036
rect 22520 46996 22526 47008
rect 22557 47005 22569 47008
rect 22603 47005 22615 47039
rect 22557 46999 22615 47005
rect 23842 46996 23848 47048
rect 23900 47036 23906 47048
rect 24581 47039 24639 47045
rect 24581 47036 24593 47039
rect 23900 47008 24593 47036
rect 23900 46996 23906 47008
rect 24581 47005 24593 47008
rect 24627 47005 24639 47039
rect 25314 47036 25320 47048
rect 25275 47008 25320 47036
rect 24581 46999 24639 47005
rect 25314 46996 25320 47008
rect 25372 46996 25378 47048
rect 29730 46996 29736 47048
rect 29788 47036 29794 47048
rect 29825 47039 29883 47045
rect 29825 47036 29837 47039
rect 29788 47008 29837 47036
rect 29788 46996 29794 47008
rect 29825 47005 29837 47008
rect 29871 47005 29883 47039
rect 29825 46999 29883 47005
rect 31754 46996 31760 47048
rect 31812 47036 31818 47048
rect 32309 47039 32367 47045
rect 32309 47036 32321 47039
rect 31812 47008 32321 47036
rect 31812 46996 31818 47008
rect 32309 47005 32321 47008
rect 32355 47005 32367 47039
rect 33134 47036 33140 47048
rect 33095 47008 33140 47036
rect 32309 46999 32367 47005
rect 33134 46996 33140 47008
rect 33192 46996 33198 47048
rect 38930 47036 38936 47048
rect 38891 47008 38936 47036
rect 38930 46996 38936 47008
rect 38988 46996 38994 47048
rect 40126 47036 40132 47048
rect 40087 47008 40132 47036
rect 40126 46996 40132 47008
rect 40184 46996 40190 47048
rect 41506 47036 41512 47048
rect 41467 47008 41512 47036
rect 41506 46996 41512 47008
rect 41564 46996 41570 47048
rect 42518 46996 42524 47048
rect 42576 47036 42582 47048
rect 42613 47039 42671 47045
rect 42613 47036 42625 47039
rect 42576 47008 42625 47036
rect 42576 46996 42582 47008
rect 42613 47005 42625 47008
rect 42659 47005 42671 47039
rect 42613 46999 42671 47005
rect 47210 46996 47216 47048
rect 47268 47036 47274 47048
rect 48225 47039 48283 47045
rect 47268 47008 47313 47036
rect 47268 46996 47274 47008
rect 48225 47005 48237 47039
rect 48271 47036 48283 47039
rect 48958 47036 48964 47048
rect 48271 47008 48964 47036
rect 48271 47005 48283 47008
rect 48225 46999 48283 47005
rect 48958 46996 48964 47008
rect 49016 46996 49022 47048
rect 2314 46968 2320 46980
rect 2275 46940 2320 46968
rect 2314 46928 2320 46940
rect 2372 46928 2378 46980
rect 4065 46971 4123 46977
rect 4065 46968 4077 46971
rect 2746 46940 4077 46968
rect 1302 46860 1308 46912
rect 1360 46900 1366 46912
rect 2746 46900 2774 46940
rect 4065 46937 4077 46940
rect 4111 46937 4123 46971
rect 4065 46931 4123 46937
rect 4433 46971 4491 46977
rect 4433 46937 4445 46971
rect 4479 46968 4491 46971
rect 4706 46968 4712 46980
rect 4479 46940 4712 46968
rect 4479 46937 4491 46940
rect 4433 46931 4491 46937
rect 4706 46928 4712 46940
rect 4764 46928 4770 46980
rect 13814 46928 13820 46980
rect 13872 46968 13878 46980
rect 14461 46971 14519 46977
rect 14461 46968 14473 46971
rect 13872 46940 14473 46968
rect 13872 46928 13878 46940
rect 14461 46937 14473 46940
rect 14507 46937 14519 46971
rect 47026 46968 47032 46980
rect 46987 46940 47032 46968
rect 14461 46931 14519 46937
rect 47026 46928 47032 46940
rect 47084 46928 47090 46980
rect 47762 46928 47768 46980
rect 47820 46968 47826 46980
rect 47857 46971 47915 46977
rect 47857 46968 47869 46971
rect 47820 46940 47869 46968
rect 47820 46928 47826 46940
rect 47857 46937 47869 46940
rect 47903 46937 47915 46971
rect 47857 46931 47915 46937
rect 1360 46872 2774 46900
rect 3329 46903 3387 46909
rect 1360 46860 1366 46872
rect 3329 46869 3341 46903
rect 3375 46900 3387 46903
rect 3510 46900 3516 46912
rect 3375 46872 3516 46900
rect 3375 46869 3387 46872
rect 3329 46863 3387 46869
rect 3510 46860 3516 46872
rect 3568 46860 3574 46912
rect 32490 46900 32496 46912
rect 32451 46872 32496 46900
rect 32490 46860 32496 46872
rect 32548 46860 32554 46912
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 1946 46656 1952 46708
rect 2004 46696 2010 46708
rect 7190 46696 7196 46708
rect 2004 46668 4200 46696
rect 7151 46668 7196 46696
rect 2004 46656 2010 46668
rect 3510 46628 3516 46640
rect 3471 46600 3516 46628
rect 3510 46588 3516 46600
rect 3568 46588 3574 46640
rect 4172 46637 4200 46668
rect 7190 46656 7196 46668
rect 7248 46656 7254 46708
rect 33134 46656 33140 46708
rect 33192 46656 33198 46708
rect 4157 46631 4215 46637
rect 4157 46597 4169 46631
rect 4203 46597 4215 46631
rect 4157 46591 4215 46597
rect 4614 46588 4620 46640
rect 4672 46628 4678 46640
rect 12434 46628 12440 46640
rect 4672 46600 8432 46628
rect 4672 46588 4678 46600
rect 3697 46563 3755 46569
rect 3697 46529 3709 46563
rect 3743 46560 3755 46563
rect 4522 46560 4528 46572
rect 3743 46532 4528 46560
rect 3743 46529 3755 46532
rect 3697 46523 3755 46529
rect 4522 46520 4528 46532
rect 4580 46520 4586 46572
rect 5994 46520 6000 46572
rect 6052 46560 6058 46572
rect 7377 46563 7435 46569
rect 6052 46532 6097 46560
rect 6052 46520 6058 46532
rect 7377 46529 7389 46563
rect 7423 46529 7435 46563
rect 7377 46523 7435 46529
rect 2590 46492 2596 46504
rect 2551 46464 2596 46492
rect 2590 46452 2596 46464
rect 2648 46452 2654 46504
rect 5810 46492 5816 46504
rect 5771 46464 5816 46492
rect 5810 46452 5816 46464
rect 5868 46452 5874 46504
rect 4062 46384 4068 46436
rect 4120 46424 4126 46436
rect 7392 46424 7420 46523
rect 4120 46396 7420 46424
rect 8404 46424 8432 46600
rect 12084 46600 12440 46628
rect 12084 46569 12112 46600
rect 12434 46588 12440 46600
rect 12492 46588 12498 46640
rect 25314 46628 25320 46640
rect 24780 46600 25320 46628
rect 12069 46563 12127 46569
rect 12069 46529 12081 46563
rect 12115 46529 12127 46563
rect 22462 46560 22468 46572
rect 22423 46532 22468 46560
rect 12069 46523 12127 46529
rect 22462 46520 22468 46532
rect 22520 46520 22526 46572
rect 24780 46569 24808 46600
rect 25314 46588 25320 46600
rect 25372 46588 25378 46640
rect 33152 46628 33180 46656
rect 33060 46600 33180 46628
rect 33060 46569 33088 46600
rect 24765 46563 24823 46569
rect 24765 46529 24777 46563
rect 24811 46529 24823 46563
rect 24765 46523 24823 46529
rect 33045 46563 33103 46569
rect 33045 46529 33057 46563
rect 33091 46529 33103 46563
rect 39758 46560 39764 46572
rect 39719 46532 39764 46560
rect 33045 46523 33103 46529
rect 39758 46520 39764 46532
rect 39816 46520 39822 46572
rect 41506 46520 41512 46572
rect 41564 46560 41570 46572
rect 42613 46563 42671 46569
rect 42613 46560 42625 46563
rect 41564 46532 42625 46560
rect 41564 46520 41570 46532
rect 42613 46529 42625 46532
rect 42659 46529 42671 46563
rect 42613 46523 42671 46529
rect 47394 46520 47400 46572
rect 47452 46560 47458 46572
rect 47765 46563 47823 46569
rect 47765 46560 47777 46563
rect 47452 46532 47777 46560
rect 47452 46520 47458 46532
rect 47765 46529 47777 46532
rect 47811 46529 47823 46563
rect 47765 46523 47823 46529
rect 12253 46495 12311 46501
rect 12253 46461 12265 46495
rect 12299 46492 12311 46495
rect 12894 46492 12900 46504
rect 12299 46464 12900 46492
rect 12299 46461 12311 46464
rect 12253 46455 12311 46461
rect 12894 46452 12900 46464
rect 12952 46452 12958 46504
rect 12986 46452 12992 46504
rect 13044 46492 13050 46504
rect 14366 46492 14372 46504
rect 13044 46464 13089 46492
rect 14327 46464 14372 46492
rect 13044 46452 13050 46464
rect 14366 46452 14372 46464
rect 14424 46452 14430 46504
rect 14550 46492 14556 46504
rect 14511 46464 14556 46492
rect 14550 46452 14556 46464
rect 14608 46452 14614 46504
rect 14826 46492 14832 46504
rect 14787 46464 14832 46492
rect 14826 46452 14832 46464
rect 14884 46452 14890 46504
rect 22646 46492 22652 46504
rect 22607 46464 22652 46492
rect 22646 46452 22652 46464
rect 22704 46452 22710 46504
rect 23198 46492 23204 46504
rect 23159 46464 23204 46492
rect 23198 46452 23204 46464
rect 23256 46452 23262 46504
rect 24946 46492 24952 46504
rect 24907 46464 24952 46492
rect 24946 46452 24952 46464
rect 25004 46452 25010 46504
rect 25774 46492 25780 46504
rect 25735 46464 25780 46492
rect 25774 46452 25780 46464
rect 25832 46452 25838 46504
rect 28721 46495 28779 46501
rect 28721 46461 28733 46495
rect 28767 46492 28779 46495
rect 29181 46495 29239 46501
rect 29181 46492 29193 46495
rect 28767 46464 29193 46492
rect 28767 46461 28779 46464
rect 28721 46455 28779 46461
rect 29181 46461 29193 46464
rect 29227 46461 29239 46495
rect 29362 46492 29368 46504
rect 29323 46464 29368 46492
rect 29181 46455 29239 46461
rect 29362 46452 29368 46464
rect 29420 46452 29426 46504
rect 29638 46492 29644 46504
rect 29599 46464 29644 46492
rect 29638 46452 29644 46464
rect 29696 46452 29702 46504
rect 33226 46492 33232 46504
rect 33187 46464 33232 46492
rect 33226 46452 33232 46464
rect 33284 46452 33290 46504
rect 33502 46492 33508 46504
rect 33463 46464 33508 46492
rect 33502 46452 33508 46464
rect 33560 46452 33566 46504
rect 36265 46495 36323 46501
rect 36265 46461 36277 46495
rect 36311 46492 36323 46495
rect 37461 46495 37519 46501
rect 37461 46492 37473 46495
rect 36311 46464 37473 46492
rect 36311 46461 36323 46464
rect 36265 46455 36323 46461
rect 37461 46461 37473 46464
rect 37507 46461 37519 46495
rect 37642 46492 37648 46504
rect 37603 46464 37648 46492
rect 37461 46455 37519 46461
rect 37642 46452 37648 46464
rect 37700 46452 37706 46504
rect 37921 46495 37979 46501
rect 37921 46461 37933 46495
rect 37967 46461 37979 46495
rect 39942 46492 39948 46504
rect 39903 46464 39948 46492
rect 37921 46455 37979 46461
rect 8404 46396 13032 46424
rect 4120 46384 4126 46396
rect 13004 46368 13032 46396
rect 36722 46384 36728 46436
rect 36780 46424 36786 46436
rect 37936 46424 37964 46455
rect 39942 46452 39948 46464
rect 40000 46452 40006 46504
rect 40221 46495 40279 46501
rect 40221 46461 40233 46495
rect 40267 46461 40279 46495
rect 42794 46492 42800 46504
rect 42755 46464 42800 46492
rect 40221 46455 40279 46461
rect 36780 46396 37964 46424
rect 36780 46384 36786 46396
rect 38654 46384 38660 46436
rect 38712 46424 38718 46436
rect 40236 46424 40264 46455
rect 42794 46452 42800 46464
rect 42852 46452 42858 46504
rect 43073 46495 43131 46501
rect 43073 46461 43085 46495
rect 43119 46461 43131 46495
rect 43073 46455 43131 46461
rect 45373 46495 45431 46501
rect 45373 46461 45385 46495
rect 45419 46461 45431 46495
rect 45373 46455 45431 46461
rect 45557 46495 45615 46501
rect 45557 46461 45569 46495
rect 45603 46492 45615 46495
rect 45922 46492 45928 46504
rect 45603 46464 45928 46492
rect 45603 46461 45615 46464
rect 45557 46455 45615 46461
rect 38712 46396 40264 46424
rect 38712 46384 38718 46396
rect 41874 46384 41880 46436
rect 41932 46424 41938 46436
rect 43088 46424 43116 46455
rect 41932 46396 43116 46424
rect 45388 46424 45416 46455
rect 45922 46452 45928 46464
rect 45980 46452 45986 46504
rect 46382 46492 46388 46504
rect 46343 46464 46388 46492
rect 46382 46452 46388 46464
rect 46440 46452 46446 46504
rect 45830 46424 45836 46436
rect 45388 46396 45836 46424
rect 41932 46384 41938 46396
rect 45830 46384 45836 46396
rect 45888 46384 45894 46436
rect 4890 46316 4896 46368
rect 4948 46356 4954 46368
rect 6549 46359 6607 46365
rect 6549 46356 6561 46359
rect 4948 46328 6561 46356
rect 4948 46316 4954 46328
rect 6549 46325 6561 46328
rect 6595 46325 6607 46359
rect 10502 46356 10508 46368
rect 10463 46328 10508 46356
rect 6549 46319 6607 46325
rect 10502 46316 10508 46328
rect 10560 46316 10566 46368
rect 12986 46316 12992 46368
rect 13044 46316 13050 46368
rect 16850 46356 16856 46368
rect 16811 46328 16856 46356
rect 16850 46316 16856 46328
rect 16908 46316 16914 46368
rect 19242 46316 19248 46368
rect 19300 46356 19306 46368
rect 27062 46356 27068 46368
rect 19300 46328 27068 46356
rect 19300 46316 19306 46328
rect 27062 46316 27068 46328
rect 27120 46316 27126 46368
rect 35342 46316 35348 46368
rect 35400 46356 35406 46368
rect 35437 46359 35495 46365
rect 35437 46356 35449 46359
rect 35400 46328 35449 46356
rect 35400 46316 35406 46328
rect 35437 46325 35449 46328
rect 35483 46325 35495 46359
rect 35437 46319 35495 46325
rect 46658 46316 46664 46368
rect 46716 46356 46722 46368
rect 47857 46359 47915 46365
rect 47857 46356 47869 46359
rect 46716 46328 47869 46356
rect 46716 46316 46722 46328
rect 47857 46325 47869 46328
rect 47903 46325 47915 46359
rect 47857 46319 47915 46325
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 5810 46112 5816 46164
rect 5868 46152 5874 46164
rect 6273 46155 6331 46161
rect 6273 46152 6285 46155
rect 5868 46124 6285 46152
rect 5868 46112 5874 46124
rect 6273 46121 6285 46124
rect 6319 46121 6331 46155
rect 12894 46152 12900 46164
rect 12855 46124 12900 46152
rect 6273 46115 6331 46121
rect 12894 46112 12900 46124
rect 12952 46112 12958 46164
rect 13633 46155 13691 46161
rect 13633 46121 13645 46155
rect 13679 46152 13691 46155
rect 13814 46152 13820 46164
rect 13679 46124 13820 46152
rect 13679 46121 13691 46124
rect 13633 46115 13691 46121
rect 13814 46112 13820 46124
rect 13872 46112 13878 46164
rect 14461 46155 14519 46161
rect 14461 46121 14473 46155
rect 14507 46152 14519 46155
rect 14550 46152 14556 46164
rect 14507 46124 14556 46152
rect 14507 46121 14519 46124
rect 14461 46115 14519 46121
rect 14550 46112 14556 46124
rect 14608 46112 14614 46164
rect 22646 46152 22652 46164
rect 22607 46124 22652 46152
rect 22646 46112 22652 46124
rect 22704 46112 22710 46164
rect 29089 46155 29147 46161
rect 29089 46121 29101 46155
rect 29135 46152 29147 46155
rect 29362 46152 29368 46164
rect 29135 46124 29368 46152
rect 29135 46121 29147 46124
rect 29089 46115 29147 46121
rect 29362 46112 29368 46124
rect 29420 46112 29426 46164
rect 33226 46152 33232 46164
rect 33187 46124 33232 46152
rect 33226 46112 33232 46124
rect 33284 46112 33290 46164
rect 38381 46155 38439 46161
rect 38381 46121 38393 46155
rect 38427 46152 38439 46155
rect 39942 46152 39948 46164
rect 38427 46124 39948 46152
rect 38427 46121 38439 46124
rect 38381 46115 38439 46121
rect 39942 46112 39948 46124
rect 40000 46112 40006 46164
rect 45922 46152 45928 46164
rect 45883 46124 45928 46152
rect 45922 46112 45928 46124
rect 45980 46112 45986 46164
rect 4433 46087 4491 46093
rect 4433 46053 4445 46087
rect 4479 46084 4491 46087
rect 5074 46084 5080 46096
rect 4479 46056 5080 46084
rect 4479 46053 4491 46056
rect 4433 46047 4491 46053
rect 5074 46044 5080 46056
rect 5132 46084 5138 46096
rect 25222 46084 25228 46096
rect 5132 46056 7052 46084
rect 5132 46044 5138 46056
rect 2774 45976 2780 46028
rect 2832 46016 2838 46028
rect 3237 46019 3295 46025
rect 2832 45988 2877 46016
rect 2832 45976 2838 45988
rect 3237 45985 3249 46019
rect 3283 46016 3295 46019
rect 4614 46016 4620 46028
rect 3283 45988 4620 46016
rect 3283 45985 3295 45988
rect 3237 45979 3295 45985
rect 4614 45976 4620 45988
rect 4672 45976 4678 46028
rect 7024 45960 7052 46056
rect 23860 46056 25228 46084
rect 10502 46016 10508 46028
rect 10463 45988 10508 46016
rect 10502 45976 10508 45988
rect 10560 45976 10566 46028
rect 10962 45976 10968 46028
rect 11020 46016 11026 46028
rect 11057 46019 11115 46025
rect 11057 46016 11069 46019
rect 11020 45988 11069 46016
rect 11020 45976 11026 45988
rect 11057 45985 11069 45988
rect 11103 45985 11115 46019
rect 15470 46016 15476 46028
rect 15431 45988 15476 46016
rect 11057 45979 11115 45985
rect 15470 45976 15476 45988
rect 15528 45976 15534 46028
rect 16850 46016 16856 46028
rect 16811 45988 16856 46016
rect 16850 45976 16856 45988
rect 16908 45976 16914 46028
rect 23860 46016 23888 46056
rect 25222 46044 25228 46056
rect 25280 46044 25286 46096
rect 33152 46056 39988 46084
rect 25130 46016 25136 46028
rect 21928 45988 23888 46016
rect 25091 45988 25136 46016
rect 3421 45951 3479 45957
rect 3421 45917 3433 45951
rect 3467 45948 3479 45951
rect 4798 45948 4804 45960
rect 3467 45920 4804 45948
rect 3467 45917 3479 45920
rect 3421 45911 3479 45917
rect 4798 45908 4804 45920
rect 4856 45908 4862 45960
rect 6362 45948 6368 45960
rect 6275 45920 6368 45948
rect 6362 45908 6368 45920
rect 6420 45948 6426 45960
rect 7006 45948 7012 45960
rect 6420 45920 6868 45948
rect 6967 45920 7012 45948
rect 6420 45908 6426 45920
rect 5534 45840 5540 45892
rect 5592 45880 5598 45892
rect 5721 45883 5779 45889
rect 5721 45880 5733 45883
rect 5592 45852 5733 45880
rect 5592 45840 5598 45852
rect 5721 45849 5733 45852
rect 5767 45849 5779 45883
rect 6840 45880 6868 45920
rect 7006 45908 7012 45920
rect 7064 45908 7070 45960
rect 12989 45951 13047 45957
rect 12989 45917 13001 45951
rect 13035 45948 13047 45951
rect 13262 45948 13268 45960
rect 13035 45920 13268 45948
rect 13035 45917 13047 45920
rect 12989 45911 13047 45917
rect 13262 45908 13268 45920
rect 13320 45948 13326 45960
rect 13541 45951 13599 45957
rect 13541 45948 13553 45951
rect 13320 45920 13553 45948
rect 13320 45908 13326 45920
rect 13541 45917 13553 45920
rect 13587 45917 13599 45951
rect 14369 45951 14427 45957
rect 14369 45948 14381 45951
rect 13541 45911 13599 45917
rect 13648 45920 14381 45948
rect 10686 45880 10692 45892
rect 6840 45852 7052 45880
rect 10647 45852 10692 45880
rect 5721 45843 5779 45849
rect 6914 45812 6920 45824
rect 6875 45784 6920 45812
rect 6914 45772 6920 45784
rect 6972 45772 6978 45824
rect 7024 45812 7052 45852
rect 10686 45840 10692 45852
rect 10744 45840 10750 45892
rect 13648 45812 13676 45920
rect 14369 45917 14381 45920
rect 14415 45917 14427 45951
rect 14369 45911 14427 45917
rect 7024 45784 13676 45812
rect 14384 45812 14412 45911
rect 16666 45880 16672 45892
rect 16627 45852 16672 45880
rect 16666 45840 16672 45852
rect 16724 45840 16730 45892
rect 21928 45812 21956 45988
rect 23860 45957 23888 45988
rect 25130 45976 25136 45988
rect 25188 45976 25194 46028
rect 29730 46016 29736 46028
rect 29691 45988 29736 46016
rect 29730 45976 29736 45988
rect 29788 45976 29794 46028
rect 30282 45976 30288 46028
rect 30340 46016 30346 46028
rect 30377 46019 30435 46025
rect 30377 46016 30389 46019
rect 30340 45988 30389 46016
rect 30340 45976 30346 45988
rect 30377 45985 30389 45988
rect 30423 45985 30435 46019
rect 30377 45979 30435 45985
rect 33152 45960 33180 46056
rect 35342 46016 35348 46028
rect 35303 45988 35348 46016
rect 35342 45976 35348 45988
rect 35400 45976 35406 46028
rect 36078 46016 36084 46028
rect 36039 45988 36084 46016
rect 36078 45976 36084 45988
rect 36136 45976 36142 46028
rect 22557 45951 22615 45957
rect 22557 45917 22569 45951
rect 22603 45917 22615 45951
rect 22557 45911 22615 45917
rect 23845 45951 23903 45957
rect 23845 45917 23857 45951
rect 23891 45917 23903 45951
rect 24578 45948 24584 45960
rect 24539 45920 24584 45948
rect 23845 45911 23903 45917
rect 22572 45824 22600 45911
rect 24578 45908 24584 45920
rect 24636 45908 24642 45960
rect 28994 45948 29000 45960
rect 28955 45920 29000 45948
rect 28994 45908 29000 45920
rect 29052 45908 29058 45960
rect 33134 45948 33140 45960
rect 33047 45920 33140 45948
rect 33134 45908 33140 45920
rect 33192 45908 33198 45960
rect 38286 45948 38292 45960
rect 38247 45920 38292 45948
rect 38286 45908 38292 45920
rect 38344 45908 38350 45960
rect 38378 45908 38384 45960
rect 38436 45948 38442 45960
rect 38933 45951 38991 45957
rect 38933 45948 38945 45951
rect 38436 45920 38945 45948
rect 38436 45908 38442 45920
rect 38933 45917 38945 45920
rect 38979 45917 38991 45951
rect 38933 45911 38991 45917
rect 23937 45883 23995 45889
rect 23937 45849 23949 45883
rect 23983 45880 23995 45883
rect 24765 45883 24823 45889
rect 24765 45880 24777 45883
rect 23983 45852 24777 45880
rect 23983 45849 23995 45852
rect 23937 45843 23995 45849
rect 24765 45849 24777 45852
rect 24811 45849 24823 45883
rect 29914 45880 29920 45892
rect 29875 45852 29920 45880
rect 24765 45843 24823 45849
rect 29914 45840 29920 45852
rect 29972 45840 29978 45892
rect 35529 45883 35587 45889
rect 35529 45849 35541 45883
rect 35575 45880 35587 45883
rect 35618 45880 35624 45892
rect 35575 45852 35624 45880
rect 35575 45849 35587 45852
rect 35529 45843 35587 45849
rect 35618 45840 35624 45852
rect 35676 45840 35682 45892
rect 14384 45784 21956 45812
rect 22554 45772 22560 45824
rect 22612 45812 22618 45824
rect 25314 45812 25320 45824
rect 22612 45784 25320 45812
rect 22612 45772 22618 45784
rect 25314 45772 25320 45784
rect 25372 45772 25378 45824
rect 39025 45815 39083 45821
rect 39025 45781 39037 45815
rect 39071 45812 39083 45815
rect 39114 45812 39120 45824
rect 39071 45784 39120 45812
rect 39071 45781 39083 45784
rect 39025 45775 39083 45781
rect 39114 45772 39120 45784
rect 39172 45772 39178 45824
rect 39960 45812 39988 46056
rect 40126 46016 40132 46028
rect 40087 45988 40132 46016
rect 40126 45976 40132 45988
rect 40184 45976 40190 46028
rect 40586 46016 40592 46028
rect 40547 45988 40592 46016
rect 40586 45976 40592 45988
rect 40644 45976 40650 46028
rect 45373 46019 45431 46025
rect 45373 45985 45385 46019
rect 45419 46016 45431 46019
rect 46477 46019 46535 46025
rect 46477 46016 46489 46019
rect 45419 45988 46489 46016
rect 45419 45985 45431 45988
rect 45373 45979 45431 45985
rect 46477 45985 46489 45988
rect 46523 45985 46535 46019
rect 46658 46016 46664 46028
rect 46619 45988 46664 46016
rect 46477 45979 46535 45985
rect 46658 45976 46664 45988
rect 46716 45976 46722 46028
rect 48314 46016 48320 46028
rect 48275 45988 48320 46016
rect 48314 45976 48320 45988
rect 48372 45976 48378 46028
rect 46014 45948 46020 45960
rect 45975 45920 46020 45948
rect 46014 45908 46020 45920
rect 46072 45908 46078 45960
rect 40310 45880 40316 45892
rect 40271 45852 40316 45880
rect 40310 45840 40316 45852
rect 40368 45840 40374 45892
rect 47394 45812 47400 45824
rect 39960 45784 47400 45812
rect 47394 45772 47400 45784
rect 47452 45772 47458 45824
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 10597 45611 10655 45617
rect 10597 45577 10609 45611
rect 10643 45608 10655 45611
rect 10686 45608 10692 45620
rect 10643 45580 10692 45608
rect 10643 45577 10655 45580
rect 10597 45571 10655 45577
rect 10686 45568 10692 45580
rect 10744 45568 10750 45620
rect 24946 45568 24952 45620
rect 25004 45608 25010 45620
rect 25225 45611 25283 45617
rect 25225 45608 25237 45611
rect 25004 45580 25237 45608
rect 25004 45568 25010 45580
rect 25225 45577 25237 45580
rect 25271 45577 25283 45611
rect 25225 45571 25283 45577
rect 25314 45568 25320 45620
rect 25372 45608 25378 45620
rect 38378 45608 38384 45620
rect 25372 45580 38384 45608
rect 25372 45568 25378 45580
rect 38378 45568 38384 45580
rect 38436 45568 38442 45620
rect 3789 45543 3847 45549
rect 3789 45509 3801 45543
rect 3835 45540 3847 45543
rect 6914 45540 6920 45552
rect 3835 45512 6920 45540
rect 3835 45509 3847 45512
rect 3789 45503 3847 45509
rect 6914 45500 6920 45512
rect 6972 45500 6978 45552
rect 7006 45500 7012 45552
rect 7064 45540 7070 45552
rect 29914 45540 29920 45552
rect 7064 45512 26234 45540
rect 29875 45512 29920 45540
rect 7064 45500 7070 45512
rect 4985 45475 5043 45481
rect 4985 45441 4997 45475
rect 5031 45472 5043 45475
rect 5534 45472 5540 45484
rect 5031 45444 5540 45472
rect 5031 45441 5043 45444
rect 4985 45435 5043 45441
rect 5534 45432 5540 45444
rect 5592 45432 5598 45484
rect 6730 45472 6736 45484
rect 6691 45444 6736 45472
rect 6730 45432 6736 45444
rect 6788 45432 6794 45484
rect 10505 45475 10563 45481
rect 10505 45472 10517 45475
rect 9646 45444 10517 45472
rect 2866 45404 2872 45416
rect 2827 45376 2872 45404
rect 2866 45364 2872 45376
rect 2924 45364 2930 45416
rect 3973 45407 4031 45413
rect 3973 45373 3985 45407
rect 4019 45404 4031 45407
rect 4890 45404 4896 45416
rect 4019 45376 4896 45404
rect 4019 45373 4031 45376
rect 3973 45367 4031 45373
rect 4890 45364 4896 45376
rect 4948 45364 4954 45416
rect 5350 45364 5356 45416
rect 5408 45404 5414 45416
rect 5445 45407 5503 45413
rect 5445 45404 5457 45407
rect 5408 45376 5457 45404
rect 5408 45364 5414 45376
rect 5445 45373 5457 45376
rect 5491 45404 5503 45407
rect 6362 45404 6368 45416
rect 5491 45376 6368 45404
rect 5491 45373 5503 45376
rect 5445 45367 5503 45373
rect 6362 45364 6368 45376
rect 6420 45364 6426 45416
rect 7374 45404 7380 45416
rect 7335 45376 7380 45404
rect 7374 45364 7380 45376
rect 7432 45364 7438 45416
rect 9646 45336 9674 45444
rect 10505 45441 10517 45444
rect 10551 45472 10563 45475
rect 10551 45444 12480 45472
rect 10551 45441 10563 45444
rect 10505 45435 10563 45441
rect 5460 45308 9674 45336
rect 12452 45336 12480 45444
rect 14366 45432 14372 45484
rect 14424 45472 14430 45484
rect 14461 45475 14519 45481
rect 14461 45472 14473 45475
rect 14424 45444 14473 45472
rect 14424 45432 14430 45444
rect 14461 45441 14473 45444
rect 14507 45441 14519 45475
rect 15102 45472 15108 45484
rect 15063 45444 15108 45472
rect 14461 45435 14519 45441
rect 15102 45432 15108 45444
rect 15160 45432 15166 45484
rect 15197 45475 15255 45481
rect 15197 45441 15209 45475
rect 15243 45472 15255 45475
rect 16666 45472 16672 45484
rect 15243 45444 16672 45472
rect 15243 45441 15255 45444
rect 15197 45435 15255 45441
rect 16666 45432 16672 45444
rect 16724 45432 16730 45484
rect 24578 45432 24584 45484
rect 24636 45472 24642 45484
rect 24673 45475 24731 45481
rect 24673 45472 24685 45475
rect 24636 45444 24685 45472
rect 24636 45432 24642 45444
rect 24673 45441 24685 45444
rect 24719 45441 24731 45475
rect 24673 45435 24731 45441
rect 25222 45432 25228 45484
rect 25280 45472 25286 45484
rect 25317 45475 25375 45481
rect 25317 45472 25329 45475
rect 25280 45444 25329 45472
rect 25280 45432 25286 45444
rect 25317 45441 25329 45444
rect 25363 45441 25375 45475
rect 26206 45472 26234 45512
rect 29914 45500 29920 45512
rect 29972 45500 29978 45552
rect 35618 45540 35624 45552
rect 35579 45512 35624 45540
rect 35618 45500 35624 45512
rect 35676 45500 35682 45552
rect 36265 45543 36323 45549
rect 36265 45509 36277 45543
rect 36311 45540 36323 45543
rect 37642 45540 37648 45552
rect 36311 45512 37648 45540
rect 36311 45509 36323 45512
rect 36265 45503 36323 45509
rect 37642 45500 37648 45512
rect 37700 45500 37706 45552
rect 39114 45540 39120 45552
rect 39075 45512 39120 45540
rect 39114 45500 39120 45512
rect 39172 45500 39178 45552
rect 41601 45543 41659 45549
rect 41601 45509 41613 45543
rect 41647 45540 41659 45543
rect 42794 45540 42800 45552
rect 41647 45512 42800 45540
rect 41647 45509 41659 45512
rect 41601 45503 41659 45509
rect 42794 45500 42800 45512
rect 42852 45500 42858 45552
rect 46934 45540 46940 45552
rect 45526 45512 46940 45540
rect 29822 45472 29828 45484
rect 26206 45444 29828 45472
rect 25317 45435 25375 45441
rect 29822 45432 29828 45444
rect 29880 45432 29886 45484
rect 35713 45475 35771 45481
rect 35713 45441 35725 45475
rect 35759 45441 35771 45475
rect 35713 45435 35771 45441
rect 36173 45475 36231 45481
rect 36173 45441 36185 45475
rect 36219 45472 36231 45475
rect 37274 45472 37280 45484
rect 36219 45444 37280 45472
rect 36219 45441 36231 45444
rect 36173 45435 36231 45441
rect 12526 45364 12532 45416
rect 12584 45404 12590 45416
rect 22554 45404 22560 45416
rect 12584 45376 22560 45404
rect 12584 45364 12590 45376
rect 22554 45364 22560 45376
rect 22612 45364 22618 45416
rect 28994 45336 29000 45348
rect 12452 45308 29000 45336
rect 5460 45280 5488 45308
rect 28994 45296 29000 45308
rect 29052 45296 29058 45348
rect 35728 45280 35756 45435
rect 37274 45432 37280 45444
rect 37332 45472 37338 45484
rect 38286 45472 38292 45484
rect 37332 45444 38292 45472
rect 37332 45432 37338 45444
rect 38286 45432 38292 45444
rect 38344 45432 38350 45484
rect 38930 45472 38936 45484
rect 38891 45444 38936 45472
rect 38930 45432 38936 45444
rect 38988 45432 38994 45484
rect 41509 45475 41567 45481
rect 41509 45472 41521 45475
rect 40696 45444 41521 45472
rect 40126 45364 40132 45416
rect 40184 45404 40190 45416
rect 40696 45404 40724 45444
rect 41509 45441 41521 45444
rect 41555 45472 41567 45475
rect 45526 45472 45554 45512
rect 46934 45500 46940 45512
rect 46992 45500 46998 45552
rect 47026 45500 47032 45552
rect 47084 45540 47090 45552
rect 47121 45543 47179 45549
rect 47121 45540 47133 45543
rect 47084 45512 47133 45540
rect 47084 45500 47090 45512
rect 47121 45509 47133 45512
rect 47167 45509 47179 45543
rect 47121 45503 47179 45509
rect 41555 45444 45554 45472
rect 41555 45441 41567 45444
rect 41509 45435 41567 45441
rect 45830 45432 45836 45484
rect 45888 45472 45894 45484
rect 45925 45475 45983 45481
rect 45925 45472 45937 45475
rect 45888 45444 45937 45472
rect 45888 45432 45894 45444
rect 45925 45441 45937 45444
rect 45971 45441 45983 45475
rect 45925 45435 45983 45441
rect 47213 45475 47271 45481
rect 47213 45441 47225 45475
rect 47259 45472 47271 45475
rect 47394 45472 47400 45484
rect 47259 45444 47400 45472
rect 47259 45441 47271 45444
rect 47213 45435 47271 45441
rect 47394 45432 47400 45444
rect 47452 45432 47458 45484
rect 40184 45376 40724 45404
rect 40773 45407 40831 45413
rect 40184 45364 40190 45376
rect 40773 45373 40785 45407
rect 40819 45404 40831 45407
rect 46290 45404 46296 45416
rect 40819 45376 46296 45404
rect 40819 45373 40831 45376
rect 40773 45367 40831 45373
rect 46290 45364 46296 45376
rect 46348 45364 46354 45416
rect 5442 45228 5448 45280
rect 5500 45228 5506 45280
rect 6730 45228 6736 45280
rect 6788 45268 6794 45280
rect 12526 45268 12532 45280
rect 6788 45240 12532 45268
rect 6788 45228 6794 45240
rect 12526 45228 12532 45240
rect 12584 45228 12590 45280
rect 25222 45228 25228 45280
rect 25280 45268 25286 45280
rect 35710 45268 35716 45280
rect 25280 45240 35716 45268
rect 25280 45228 25286 45240
rect 35710 45228 35716 45240
rect 35768 45228 35774 45280
rect 47949 45271 48007 45277
rect 47949 45237 47961 45271
rect 47995 45268 48007 45271
rect 48314 45268 48320 45280
rect 47995 45240 48320 45268
rect 47995 45237 48007 45240
rect 47949 45231 48007 45237
rect 48314 45228 48320 45240
rect 48372 45228 48378 45280
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 4982 45024 4988 45076
rect 5040 45064 5046 45076
rect 5261 45067 5319 45073
rect 5261 45064 5273 45067
rect 5040 45036 5273 45064
rect 5040 45024 5046 45036
rect 5261 45033 5273 45036
rect 5307 45064 5319 45067
rect 5442 45064 5448 45076
rect 5307 45036 5448 45064
rect 5307 45033 5319 45036
rect 5261 45027 5319 45033
rect 5442 45024 5448 45036
rect 5500 45024 5506 45076
rect 15102 45024 15108 45076
rect 15160 45064 15166 45076
rect 40126 45064 40132 45076
rect 15160 45036 40132 45064
rect 15160 45024 15166 45036
rect 40126 45024 40132 45036
rect 40184 45024 40190 45076
rect 40310 45024 40316 45076
rect 40368 45064 40374 45076
rect 40405 45067 40463 45073
rect 40405 45064 40417 45067
rect 40368 45036 40417 45064
rect 40368 45024 40374 45036
rect 40405 45033 40417 45036
rect 40451 45033 40463 45067
rect 40405 45027 40463 45033
rect 7374 44956 7380 45008
rect 7432 44996 7438 45008
rect 7432 44968 26234 44996
rect 7432 44956 7438 44968
rect 6822 44928 6828 44940
rect 6783 44900 6828 44928
rect 6822 44888 6828 44900
rect 6880 44888 6886 44940
rect 1949 44863 2007 44869
rect 1949 44829 1961 44863
rect 1995 44860 2007 44863
rect 2038 44860 2044 44872
rect 1995 44832 2044 44860
rect 1995 44829 2007 44832
rect 1949 44823 2007 44829
rect 2038 44820 2044 44832
rect 2096 44820 2102 44872
rect 2314 44820 2320 44872
rect 2372 44860 2378 44872
rect 2409 44863 2467 44869
rect 2409 44860 2421 44863
rect 2372 44832 2421 44860
rect 2372 44820 2378 44832
rect 2409 44829 2421 44832
rect 2455 44860 2467 44863
rect 3973 44863 4031 44869
rect 3973 44860 3985 44863
rect 2455 44832 3985 44860
rect 2455 44829 2467 44832
rect 2409 44823 2467 44829
rect 3973 44829 3985 44832
rect 4019 44860 4031 44863
rect 5534 44860 5540 44872
rect 4019 44832 5540 44860
rect 4019 44829 4031 44832
rect 3973 44823 4031 44829
rect 5534 44820 5540 44832
rect 5592 44860 5598 44872
rect 6181 44863 6239 44869
rect 6181 44860 6193 44863
rect 5592 44832 6193 44860
rect 5592 44820 5598 44832
rect 6181 44829 6193 44832
rect 6227 44829 6239 44863
rect 26206 44860 26234 44968
rect 46842 44928 46848 44940
rect 46803 44900 46848 44928
rect 46842 44888 46848 44900
rect 46900 44888 46906 44940
rect 48314 44928 48320 44940
rect 48275 44900 48320 44928
rect 48314 44888 48320 44900
rect 48372 44888 48378 44940
rect 40497 44863 40555 44869
rect 40497 44860 40509 44863
rect 26206 44832 40509 44860
rect 6181 44823 6239 44829
rect 40497 44829 40509 44832
rect 40543 44860 40555 44863
rect 46014 44860 46020 44872
rect 40543 44832 46020 44860
rect 40543 44829 40555 44832
rect 40497 44823 40555 44829
rect 46014 44820 46020 44832
rect 46072 44860 46078 44872
rect 46382 44860 46388 44872
rect 46072 44832 46388 44860
rect 46072 44820 46078 44832
rect 46382 44820 46388 44832
rect 46440 44820 46446 44872
rect 3234 44792 3240 44804
rect 3195 44764 3240 44792
rect 3234 44752 3240 44764
rect 3292 44752 3298 44804
rect 47854 44752 47860 44804
rect 47912 44792 47918 44804
rect 48133 44795 48191 44801
rect 48133 44792 48145 44795
rect 47912 44764 48145 44792
rect 47912 44752 47918 44764
rect 48133 44761 48145 44764
rect 48179 44761 48191 44795
rect 48133 44755 48191 44761
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 4433 44523 4491 44529
rect 4433 44489 4445 44523
rect 4479 44520 4491 44523
rect 4614 44520 4620 44532
rect 4479 44492 4620 44520
rect 4479 44489 4491 44492
rect 4433 44483 4491 44489
rect 4614 44480 4620 44492
rect 4672 44480 4678 44532
rect 4724 44492 5672 44520
rect 3234 44412 3240 44464
rect 3292 44452 3298 44464
rect 4724 44452 4752 44492
rect 5534 44452 5540 44464
rect 3292 44424 4752 44452
rect 5000 44424 5540 44452
rect 3292 44412 3298 44424
rect 5000 44396 5028 44424
rect 5534 44412 5540 44424
rect 5592 44412 5598 44464
rect 5644 44452 5672 44492
rect 6822 44480 6828 44532
rect 6880 44520 6886 44532
rect 15102 44520 15108 44532
rect 6880 44492 15108 44520
rect 6880 44480 6886 44492
rect 15102 44480 15108 44492
rect 15160 44480 15166 44532
rect 47854 44520 47860 44532
rect 47815 44492 47860 44520
rect 47854 44480 47860 44492
rect 47912 44480 47918 44532
rect 13262 44452 13268 44464
rect 5644 44424 13268 44452
rect 13262 44412 13268 44424
rect 13320 44412 13326 44464
rect 46934 44412 46940 44464
rect 46992 44452 46998 44464
rect 46992 44424 47808 44452
rect 46992 44412 46998 44424
rect 2038 44384 2044 44396
rect 1999 44356 2044 44384
rect 2038 44344 2044 44356
rect 2096 44344 2102 44396
rect 4525 44387 4583 44393
rect 4525 44353 4537 44387
rect 4571 44353 4583 44387
rect 4982 44384 4988 44396
rect 4895 44356 4988 44384
rect 4525 44347 4583 44353
rect 2225 44319 2283 44325
rect 2225 44285 2237 44319
rect 2271 44316 2283 44319
rect 3050 44316 3056 44328
rect 2271 44288 3056 44316
rect 2271 44285 2283 44288
rect 2225 44279 2283 44285
rect 3050 44276 3056 44288
rect 3108 44276 3114 44328
rect 3142 44276 3148 44328
rect 3200 44316 3206 44328
rect 4540 44316 4568 44347
rect 4982 44344 4988 44356
rect 5040 44344 5046 44396
rect 5166 44384 5172 44396
rect 5092 44356 5172 44384
rect 5092 44316 5120 44356
rect 5166 44344 5172 44356
rect 5224 44384 5230 44396
rect 37274 44384 37280 44396
rect 5224 44356 37280 44384
rect 5224 44344 5230 44356
rect 37274 44344 37280 44356
rect 37332 44344 37338 44396
rect 47210 44384 47216 44396
rect 47171 44356 47216 44384
rect 47210 44344 47216 44356
rect 47268 44344 47274 44396
rect 47780 44393 47808 44424
rect 47765 44387 47823 44393
rect 47765 44353 47777 44387
rect 47811 44353 47823 44387
rect 47765 44347 47823 44353
rect 5810 44316 5816 44328
rect 3200 44288 3245 44316
rect 4540 44288 5120 44316
rect 5723 44288 5816 44316
rect 3200 44276 3206 44288
rect 5810 44276 5816 44288
rect 5868 44316 5874 44328
rect 33134 44316 33140 44328
rect 5868 44288 33140 44316
rect 5868 44276 5874 44288
rect 33134 44276 33140 44288
rect 33192 44276 33198 44328
rect 4614 44208 4620 44260
rect 4672 44248 4678 44260
rect 5074 44248 5080 44260
rect 4672 44220 5080 44248
rect 4672 44208 4678 44220
rect 5074 44208 5080 44220
rect 5132 44208 5138 44260
rect 6733 44183 6791 44189
rect 6733 44149 6745 44183
rect 6779 44180 6791 44183
rect 7282 44180 7288 44192
rect 6779 44152 7288 44180
rect 6779 44149 6791 44152
rect 6733 44143 6791 44149
rect 7282 44140 7288 44152
rect 7340 44140 7346 44192
rect 28994 44140 29000 44192
rect 29052 44180 29058 44192
rect 29638 44180 29644 44192
rect 29052 44152 29644 44180
rect 29052 44140 29058 44152
rect 29638 44140 29644 44152
rect 29696 44140 29702 44192
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 3053 43843 3111 43849
rect 3053 43809 3065 43843
rect 3099 43840 3111 43843
rect 3510 43840 3516 43852
rect 3099 43812 3516 43840
rect 3099 43809 3111 43812
rect 3053 43803 3111 43809
rect 3510 43800 3516 43812
rect 3568 43800 3574 43852
rect 4617 43843 4675 43849
rect 4617 43809 4629 43843
rect 4663 43840 4675 43843
rect 5258 43840 5264 43852
rect 4663 43812 5264 43840
rect 4663 43809 4675 43812
rect 4617 43803 4675 43809
rect 5258 43800 5264 43812
rect 5316 43800 5322 43852
rect 5718 43840 5724 43852
rect 5679 43812 5724 43840
rect 5718 43800 5724 43812
rect 5776 43800 5782 43852
rect 7282 43840 7288 43852
rect 7243 43812 7288 43840
rect 7282 43800 7288 43812
rect 7340 43800 7346 43852
rect 1949 43775 2007 43781
rect 1949 43741 1961 43775
rect 1995 43772 2007 43775
rect 2038 43772 2044 43784
rect 1995 43744 2044 43772
rect 1995 43741 2007 43744
rect 1949 43735 2007 43741
rect 2038 43732 2044 43744
rect 2096 43732 2102 43784
rect 3421 43775 3479 43781
rect 3421 43741 3433 43775
rect 3467 43772 3479 43775
rect 4982 43772 4988 43784
rect 3467 43744 4988 43772
rect 3467 43741 3479 43744
rect 3421 43735 3479 43741
rect 4982 43732 4988 43744
rect 5040 43732 5046 43784
rect 5902 43664 5908 43716
rect 5960 43704 5966 43716
rect 7101 43707 7159 43713
rect 7101 43704 7113 43707
rect 5960 43676 7113 43704
rect 5960 43664 5966 43676
rect 7101 43673 7113 43676
rect 7147 43673 7159 43707
rect 7101 43667 7159 43673
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 5902 43432 5908 43444
rect 5863 43404 5908 43432
rect 5902 43392 5908 43404
rect 5960 43392 5966 43444
rect 5166 43364 5172 43376
rect 5127 43336 5172 43364
rect 5166 43324 5172 43336
rect 5224 43324 5230 43376
rect 6730 43364 6736 43376
rect 5736 43336 6736 43364
rect 2038 43296 2044 43308
rect 1999 43268 2044 43296
rect 2038 43256 2044 43268
rect 2096 43256 2102 43308
rect 3510 43256 3516 43308
rect 3568 43296 3574 43308
rect 4525 43299 4583 43305
rect 4525 43296 4537 43299
rect 3568 43268 4537 43296
rect 3568 43256 3574 43268
rect 4525 43265 4537 43268
rect 4571 43296 4583 43299
rect 5736 43296 5764 43336
rect 6730 43324 6736 43336
rect 6788 43324 6794 43376
rect 5994 43296 6000 43308
rect 4571 43268 5764 43296
rect 5955 43268 6000 43296
rect 4571 43265 4583 43268
rect 4525 43259 4583 43265
rect 5994 43256 6000 43268
rect 6052 43256 6058 43308
rect 29822 43256 29828 43308
rect 29880 43296 29886 43308
rect 47670 43296 47676 43308
rect 29880 43268 47676 43296
rect 29880 43256 29886 43268
rect 47670 43256 47676 43268
rect 47728 43296 47734 43308
rect 47765 43299 47823 43305
rect 47765 43296 47777 43299
rect 47728 43268 47777 43296
rect 47728 43256 47734 43268
rect 47765 43265 47777 43268
rect 47811 43265 47823 43299
rect 47765 43259 47823 43265
rect 2222 43228 2228 43240
rect 2183 43200 2228 43228
rect 2222 43188 2228 43200
rect 2280 43188 2286 43240
rect 2774 43188 2780 43240
rect 2832 43228 2838 43240
rect 2832 43200 2877 43228
rect 2832 43188 2838 43200
rect 47026 43092 47032 43104
rect 46987 43064 47032 43092
rect 47026 43052 47032 43064
rect 47084 43052 47090 43104
rect 47854 43092 47860 43104
rect 47815 43064 47860 43092
rect 47854 43052 47860 43064
rect 47912 43052 47918 43104
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 2222 42848 2228 42900
rect 2280 42888 2286 42900
rect 2409 42891 2467 42897
rect 2409 42888 2421 42891
rect 2280 42860 2421 42888
rect 2280 42848 2286 42860
rect 2409 42857 2421 42860
rect 2455 42857 2467 42891
rect 2409 42851 2467 42857
rect 3510 42820 3516 42832
rect 2746 42792 3516 42820
rect 2498 42684 2504 42696
rect 2459 42656 2504 42684
rect 2498 42644 2504 42656
rect 2556 42684 2562 42696
rect 2746 42684 2774 42792
rect 3510 42780 3516 42792
rect 3568 42780 3574 42832
rect 3050 42752 3056 42764
rect 3011 42724 3056 42752
rect 3050 42712 3056 42724
rect 3108 42712 3114 42764
rect 5258 42752 5264 42764
rect 3160 42724 5264 42752
rect 3160 42693 3188 42724
rect 5258 42712 5264 42724
rect 5316 42712 5322 42764
rect 46477 42755 46535 42761
rect 46477 42721 46489 42755
rect 46523 42752 46535 42755
rect 47026 42752 47032 42764
rect 46523 42724 47032 42752
rect 46523 42721 46535 42724
rect 46477 42715 46535 42721
rect 47026 42712 47032 42724
rect 47084 42712 47090 42764
rect 48222 42752 48228 42764
rect 48183 42724 48228 42752
rect 48222 42712 48228 42724
rect 48280 42712 48286 42764
rect 2556 42656 2774 42684
rect 3145 42687 3203 42693
rect 2556 42644 2562 42656
rect 3145 42653 3157 42687
rect 3191 42653 3203 42687
rect 3145 42647 3203 42653
rect 4982 42644 4988 42696
rect 5040 42684 5046 42696
rect 5169 42687 5227 42693
rect 5169 42684 5181 42687
rect 5040 42656 5181 42684
rect 5040 42644 5046 42656
rect 5169 42653 5181 42656
rect 5215 42653 5227 42687
rect 5169 42647 5227 42653
rect 5626 42576 5632 42628
rect 5684 42616 5690 42628
rect 5721 42619 5779 42625
rect 5721 42616 5733 42619
rect 5684 42588 5733 42616
rect 5684 42576 5690 42588
rect 5721 42585 5733 42588
rect 5767 42616 5779 42619
rect 5994 42616 6000 42628
rect 5767 42588 6000 42616
rect 5767 42585 5779 42588
rect 5721 42579 5779 42585
rect 5994 42576 6000 42588
rect 6052 42616 6058 42628
rect 13078 42616 13084 42628
rect 6052 42588 13084 42616
rect 6052 42576 6058 42588
rect 13078 42576 13084 42588
rect 13136 42576 13142 42628
rect 46661 42619 46719 42625
rect 46661 42585 46673 42619
rect 46707 42616 46719 42619
rect 47854 42616 47860 42628
rect 46707 42588 47860 42616
rect 46707 42585 46719 42588
rect 46661 42579 46719 42585
rect 47854 42576 47860 42588
rect 47912 42576 47918 42628
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 5629 42007 5687 42013
rect 5629 41973 5641 42007
rect 5675 42004 5687 42007
rect 7282 42004 7288 42016
rect 5675 41976 7288 42004
rect 5675 41973 5687 41976
rect 5629 41967 5687 41973
rect 7282 41964 7288 41976
rect 7340 41964 7346 42016
rect 46474 41964 46480 42016
rect 46532 42004 46538 42016
rect 47765 42007 47823 42013
rect 47765 42004 47777 42007
rect 46532 41976 47777 42004
rect 46532 41964 46538 41976
rect 47765 41973 47777 41976
rect 47811 41973 47823 42007
rect 47765 41967 47823 41973
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 7282 41664 7288 41676
rect 7243 41636 7288 41664
rect 7282 41624 7288 41636
rect 7340 41624 7346 41676
rect 46474 41664 46480 41676
rect 46435 41636 46480 41664
rect 46474 41624 46480 41636
rect 46532 41624 46538 41676
rect 48222 41664 48228 41676
rect 48183 41636 48228 41664
rect 48222 41624 48228 41636
rect 48280 41624 48286 41676
rect 3050 41488 3056 41540
rect 3108 41528 3114 41540
rect 5445 41531 5503 41537
rect 5445 41528 5457 41531
rect 3108 41500 5457 41528
rect 3108 41488 3114 41500
rect 5445 41497 5457 41500
rect 5491 41497 5503 41531
rect 7098 41528 7104 41540
rect 7059 41500 7104 41528
rect 5445 41491 5503 41497
rect 7098 41488 7104 41500
rect 7156 41488 7162 41540
rect 46661 41531 46719 41537
rect 46661 41497 46673 41531
rect 46707 41528 46719 41531
rect 47118 41528 47124 41540
rect 46707 41500 47124 41528
rect 46707 41497 46719 41500
rect 46661 41491 46719 41497
rect 47118 41488 47124 41500
rect 47176 41488 47182 41540
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 6641 41259 6699 41265
rect 6641 41225 6653 41259
rect 6687 41256 6699 41259
rect 7098 41256 7104 41268
rect 6687 41228 7104 41256
rect 6687 41225 6699 41228
rect 6641 41219 6699 41225
rect 7098 41216 7104 41228
rect 7156 41216 7162 41268
rect 47118 41256 47124 41268
rect 47079 41228 47124 41256
rect 47118 41216 47124 41228
rect 47176 41216 47182 41268
rect 6086 41080 6092 41132
rect 6144 41120 6150 41132
rect 6549 41123 6607 41129
rect 6549 41120 6561 41123
rect 6144 41092 6561 41120
rect 6144 41080 6150 41092
rect 6549 41089 6561 41092
rect 6595 41120 6607 41123
rect 7374 41120 7380 41132
rect 6595 41092 7380 41120
rect 6595 41089 6607 41092
rect 6549 41083 6607 41089
rect 7374 41080 7380 41092
rect 7432 41080 7438 41132
rect 46934 41080 46940 41132
rect 46992 41120 46998 41132
rect 47213 41123 47271 41129
rect 47213 41120 47225 41123
rect 46992 41092 47225 41120
rect 46992 41080 46998 41092
rect 47213 41089 47225 41092
rect 47259 41089 47271 41123
rect 47213 41083 47271 41089
rect 46474 40876 46480 40928
rect 46532 40916 46538 40928
rect 47765 40919 47823 40925
rect 47765 40916 47777 40919
rect 46532 40888 47777 40916
rect 46532 40876 46538 40888
rect 47765 40885 47777 40888
rect 47811 40885 47823 40919
rect 47765 40879 47823 40885
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 46474 40576 46480 40588
rect 46435 40548 46480 40576
rect 46474 40536 46480 40548
rect 46532 40536 46538 40588
rect 14734 40468 14740 40520
rect 14792 40508 14798 40520
rect 15841 40511 15899 40517
rect 15841 40508 15853 40511
rect 14792 40480 15853 40508
rect 14792 40468 14798 40480
rect 15841 40477 15853 40480
rect 15887 40477 15899 40511
rect 15841 40471 15899 40477
rect 18325 40511 18383 40517
rect 18325 40477 18337 40511
rect 18371 40508 18383 40511
rect 19058 40508 19064 40520
rect 18371 40480 19064 40508
rect 18371 40477 18383 40480
rect 18325 40471 18383 40477
rect 19058 40468 19064 40480
rect 19116 40468 19122 40520
rect 23658 40508 23664 40520
rect 23619 40480 23664 40508
rect 23658 40468 23664 40480
rect 23716 40468 23722 40520
rect 23842 40508 23848 40520
rect 23803 40480 23848 40508
rect 23842 40468 23848 40480
rect 23900 40468 23906 40520
rect 16022 40440 16028 40452
rect 15983 40412 16028 40440
rect 16022 40400 16028 40412
rect 16080 40400 16086 40452
rect 17681 40443 17739 40449
rect 17681 40409 17693 40443
rect 17727 40440 17739 40443
rect 45554 40440 45560 40452
rect 17727 40412 45560 40440
rect 17727 40409 17739 40412
rect 17681 40403 17739 40409
rect 45554 40400 45560 40412
rect 45612 40400 45618 40452
rect 46661 40443 46719 40449
rect 46661 40409 46673 40443
rect 46707 40440 46719 40443
rect 47118 40440 47124 40452
rect 46707 40412 47124 40440
rect 46707 40409 46719 40412
rect 46661 40403 46719 40409
rect 47118 40400 47124 40412
rect 47176 40400 47182 40452
rect 48314 40440 48320 40452
rect 48275 40412 48320 40440
rect 48314 40400 48320 40412
rect 48372 40400 48378 40452
rect 17770 40332 17776 40384
rect 17828 40372 17834 40384
rect 18233 40375 18291 40381
rect 18233 40372 18245 40375
rect 17828 40344 18245 40372
rect 17828 40332 17834 40344
rect 18233 40341 18245 40344
rect 18279 40341 18291 40375
rect 18233 40335 18291 40341
rect 22278 40332 22284 40384
rect 22336 40372 22342 40384
rect 23753 40375 23811 40381
rect 23753 40372 23765 40375
rect 22336 40344 23765 40372
rect 22336 40332 22342 40344
rect 23753 40341 23765 40344
rect 23799 40341 23811 40375
rect 23753 40335 23811 40341
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 16022 40168 16028 40180
rect 15983 40140 16028 40168
rect 16022 40128 16028 40140
rect 16080 40128 16086 40180
rect 22281 40171 22339 40177
rect 22281 40137 22293 40171
rect 22327 40168 22339 40171
rect 24394 40168 24400 40180
rect 22327 40140 24400 40168
rect 22327 40137 22339 40140
rect 22281 40131 22339 40137
rect 24394 40128 24400 40140
rect 24452 40128 24458 40180
rect 3234 40060 3240 40112
rect 3292 40100 3298 40112
rect 8202 40100 8208 40112
rect 3292 40072 8208 40100
rect 3292 40060 3298 40072
rect 8202 40060 8208 40072
rect 8260 40060 8266 40112
rect 12986 40100 12992 40112
rect 12947 40072 12992 40100
rect 12986 40060 12992 40072
rect 13044 40060 13050 40112
rect 17770 40100 17776 40112
rect 17731 40072 17776 40100
rect 17770 40060 17776 40072
rect 17828 40060 17834 40112
rect 22097 40103 22155 40109
rect 22097 40069 22109 40103
rect 22143 40100 22155 40103
rect 22186 40100 22192 40112
rect 22143 40072 22192 40100
rect 22143 40069 22155 40072
rect 22097 40063 22155 40069
rect 22186 40060 22192 40072
rect 22244 40060 22250 40112
rect 24026 40100 24032 40112
rect 22388 40072 24032 40100
rect 15933 40035 15991 40041
rect 15933 40001 15945 40035
rect 15979 40032 15991 40035
rect 15979 40004 16068 40032
rect 15979 40001 15991 40004
rect 15933 39995 15991 40001
rect 14642 39964 14648 39976
rect 14603 39936 14648 39964
rect 14642 39924 14648 39936
rect 14700 39924 14706 39976
rect 14829 39967 14887 39973
rect 14829 39933 14841 39967
rect 14875 39964 14887 39967
rect 14918 39964 14924 39976
rect 14875 39936 14924 39964
rect 14875 39933 14887 39936
rect 14829 39927 14887 39933
rect 14918 39924 14924 39936
rect 14976 39924 14982 39976
rect 13078 39856 13084 39908
rect 13136 39896 13142 39908
rect 16040 39896 16068 40004
rect 21726 39992 21732 40044
rect 21784 40032 21790 40044
rect 22388 40041 22416 40072
rect 24026 40060 24032 40072
rect 24084 40060 24090 40112
rect 22005 40035 22063 40041
rect 22005 40032 22017 40035
rect 21784 40004 22017 40032
rect 21784 39992 21790 40004
rect 22005 40001 22017 40004
rect 22051 40001 22063 40035
rect 22005 39995 22063 40001
rect 22373 40035 22431 40041
rect 22373 40001 22385 40035
rect 22419 40001 22431 40035
rect 23845 40035 23903 40041
rect 23845 40032 23857 40035
rect 22373 39995 22431 40001
rect 22940 40004 23857 40032
rect 16942 39924 16948 39976
rect 17000 39964 17006 39976
rect 17589 39967 17647 39973
rect 17589 39964 17601 39967
rect 17000 39936 17601 39964
rect 17000 39924 17006 39936
rect 17589 39933 17601 39936
rect 17635 39933 17647 39967
rect 19242 39964 19248 39976
rect 19203 39936 19248 39964
rect 17589 39927 17647 39933
rect 19242 39924 19248 39936
rect 19300 39924 19306 39976
rect 22189 39967 22247 39973
rect 22189 39933 22201 39967
rect 22235 39964 22247 39967
rect 22278 39964 22284 39976
rect 22235 39936 22284 39964
rect 22235 39933 22247 39936
rect 22189 39927 22247 39933
rect 22278 39924 22284 39936
rect 22336 39924 22342 39976
rect 19058 39896 19064 39908
rect 13136 39868 19064 39896
rect 13136 39856 13142 39868
rect 19058 39856 19064 39868
rect 19116 39856 19122 39908
rect 20898 39856 20904 39908
rect 20956 39896 20962 39908
rect 22940 39896 22968 40004
rect 23845 40001 23857 40004
rect 23891 40032 23903 40035
rect 24765 40035 24823 40041
rect 23891 40004 24532 40032
rect 23891 40001 23903 40004
rect 23845 39995 23903 40001
rect 24504 39976 24532 40004
rect 24765 40001 24777 40035
rect 24811 40032 24823 40035
rect 24946 40032 24952 40044
rect 24811 40004 24952 40032
rect 24811 40001 24823 40004
rect 24765 39995 24823 40001
rect 24946 39992 24952 40004
rect 25004 39992 25010 40044
rect 47118 40032 47124 40044
rect 47079 40004 47124 40032
rect 47118 39992 47124 40004
rect 47176 39992 47182 40044
rect 47213 40035 47271 40041
rect 47213 40001 47225 40035
rect 47259 40032 47271 40035
rect 47394 40032 47400 40044
rect 47259 40004 47400 40032
rect 47259 40001 47271 40004
rect 47213 39995 47271 40001
rect 23934 39964 23940 39976
rect 23895 39936 23940 39964
rect 23934 39924 23940 39936
rect 23992 39924 23998 39976
rect 24486 39964 24492 39976
rect 24399 39936 24492 39964
rect 24486 39924 24492 39936
rect 24544 39924 24550 39976
rect 46382 39924 46388 39976
rect 46440 39964 46446 39976
rect 47228 39964 47256 39995
rect 47394 39992 47400 40004
rect 47452 39992 47458 40044
rect 46440 39936 47256 39964
rect 46440 39924 46446 39936
rect 20956 39868 22968 39896
rect 20956 39856 20962 39868
rect 23014 39856 23020 39908
rect 23072 39896 23078 39908
rect 23952 39896 23980 39924
rect 24673 39899 24731 39905
rect 24673 39896 24685 39899
rect 23072 39868 23796 39896
rect 23952 39868 24685 39896
rect 23072 39856 23078 39868
rect 23569 39831 23627 39837
rect 23569 39797 23581 39831
rect 23615 39828 23627 39831
rect 23658 39828 23664 39840
rect 23615 39800 23664 39828
rect 23615 39797 23627 39800
rect 23569 39791 23627 39797
rect 23658 39788 23664 39800
rect 23716 39788 23722 39840
rect 23768 39828 23796 39868
rect 24673 39865 24685 39868
rect 24719 39865 24731 39899
rect 24673 39859 24731 39865
rect 24581 39831 24639 39837
rect 24581 39828 24593 39831
rect 23768 39800 24593 39828
rect 24581 39797 24593 39800
rect 24627 39797 24639 39831
rect 24581 39791 24639 39797
rect 47949 39831 48007 39837
rect 47949 39797 47961 39831
rect 47995 39828 48007 39831
rect 48314 39828 48320 39840
rect 47995 39800 48320 39828
rect 47995 39797 48007 39800
rect 47949 39791 48007 39797
rect 48314 39788 48320 39800
rect 48372 39788 48378 39840
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 13173 39627 13231 39633
rect 13173 39593 13185 39627
rect 13219 39624 13231 39627
rect 14642 39624 14648 39636
rect 13219 39596 14648 39624
rect 13219 39593 13231 39596
rect 13173 39587 13231 39593
rect 14642 39584 14648 39596
rect 14700 39584 14706 39636
rect 23842 39584 23848 39636
rect 23900 39624 23906 39636
rect 24581 39627 24639 39633
rect 24581 39624 24593 39627
rect 23900 39596 24593 39624
rect 23900 39584 23906 39596
rect 24581 39593 24593 39596
rect 24627 39593 24639 39627
rect 24581 39587 24639 39593
rect 23750 39516 23756 39568
rect 23808 39556 23814 39568
rect 25501 39559 25559 39565
rect 25501 39556 25513 39559
rect 23808 39528 25513 39556
rect 23808 39516 23814 39528
rect 16022 39448 16028 39500
rect 16080 39488 16086 39500
rect 21453 39491 21511 39497
rect 21453 39488 21465 39491
rect 16080 39460 21465 39488
rect 16080 39448 16086 39460
rect 21453 39457 21465 39460
rect 21499 39457 21511 39491
rect 21453 39451 21511 39457
rect 22005 39491 22063 39497
rect 22005 39457 22017 39491
rect 22051 39488 22063 39491
rect 23014 39488 23020 39500
rect 22051 39460 23020 39488
rect 22051 39457 22063 39460
rect 22005 39451 22063 39457
rect 23014 39448 23020 39460
rect 23072 39448 23078 39500
rect 23860 39497 23888 39528
rect 25501 39525 25513 39528
rect 25547 39525 25559 39559
rect 25501 39519 25559 39525
rect 23845 39491 23903 39497
rect 23845 39457 23857 39491
rect 23891 39457 23903 39491
rect 46842 39488 46848 39500
rect 46803 39460 46848 39488
rect 23845 39451 23903 39457
rect 46842 39448 46848 39460
rect 46900 39448 46906 39500
rect 48314 39488 48320 39500
rect 48275 39460 48320 39488
rect 48314 39448 48320 39460
rect 48372 39448 48378 39500
rect 13078 39420 13084 39432
rect 13039 39392 13084 39420
rect 13078 39380 13084 39392
rect 13136 39380 13142 39432
rect 21726 39420 21732 39432
rect 21687 39392 21732 39420
rect 21726 39380 21732 39392
rect 21784 39380 21790 39432
rect 22370 39420 22376 39432
rect 22331 39392 22376 39420
rect 22370 39380 22376 39392
rect 22428 39380 22434 39432
rect 22741 39423 22799 39429
rect 22741 39389 22753 39423
rect 22787 39389 22799 39423
rect 23658 39420 23664 39432
rect 23619 39392 23664 39420
rect 22741 39383 22799 39389
rect 22186 39312 22192 39364
rect 22244 39352 22250 39364
rect 22756 39352 22784 39383
rect 23658 39380 23664 39392
rect 23716 39380 23722 39432
rect 23750 39380 23756 39432
rect 23808 39420 23814 39432
rect 23937 39423 23995 39429
rect 23808 39392 23853 39420
rect 23808 39380 23814 39392
rect 23937 39389 23949 39423
rect 23983 39420 23995 39423
rect 24026 39420 24032 39432
rect 23983 39392 24032 39420
rect 23983 39389 23995 39392
rect 23937 39383 23995 39389
rect 24026 39380 24032 39392
rect 24084 39380 24090 39432
rect 24486 39380 24492 39432
rect 24544 39420 24550 39432
rect 24765 39423 24823 39429
rect 24765 39420 24777 39423
rect 24544 39392 24777 39420
rect 24544 39380 24550 39392
rect 24765 39389 24777 39392
rect 24811 39420 24823 39423
rect 25409 39423 25467 39429
rect 25409 39420 25421 39423
rect 24811 39392 25421 39420
rect 24811 39389 24823 39392
rect 24765 39383 24823 39389
rect 25409 39389 25421 39392
rect 25455 39389 25467 39423
rect 25590 39420 25596 39432
rect 25551 39392 25596 39420
rect 25409 39383 25467 39389
rect 25590 39380 25596 39392
rect 25648 39380 25654 39432
rect 22244 39324 22784 39352
rect 22244 39312 22250 39324
rect 24946 39312 24952 39364
rect 25004 39352 25010 39364
rect 25608 39352 25636 39380
rect 25004 39324 25636 39352
rect 25004 39312 25010 39324
rect 47854 39312 47860 39364
rect 47912 39352 47918 39364
rect 48133 39355 48191 39361
rect 48133 39352 48145 39355
rect 47912 39324 48145 39352
rect 47912 39312 47918 39324
rect 48133 39321 48145 39324
rect 48179 39321 48191 39355
rect 48133 39315 48191 39321
rect 23477 39287 23535 39293
rect 23477 39253 23489 39287
rect 23523 39284 23535 39287
rect 23566 39284 23572 39296
rect 23523 39256 23572 39284
rect 23523 39253 23535 39256
rect 23477 39247 23535 39253
rect 23566 39244 23572 39256
rect 23624 39244 23630 39296
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 47854 39080 47860 39092
rect 47815 39052 47860 39080
rect 47854 39040 47860 39052
rect 47912 39040 47918 39092
rect 20898 39012 20904 39024
rect 20859 38984 20904 39012
rect 20898 38972 20904 38984
rect 20956 38972 20962 39024
rect 23750 38972 23756 39024
rect 23808 39012 23814 39024
rect 24581 39015 24639 39021
rect 24581 39012 24593 39015
rect 23808 38984 24593 39012
rect 23808 38972 23814 38984
rect 24581 38981 24593 38984
rect 24627 38981 24639 39015
rect 24581 38975 24639 38981
rect 24673 39015 24731 39021
rect 24673 38981 24685 39015
rect 24719 39012 24731 39015
rect 25590 39012 25596 39024
rect 24719 38984 25596 39012
rect 24719 38981 24731 38984
rect 24673 38975 24731 38981
rect 25590 38972 25596 38984
rect 25648 38972 25654 39024
rect 1670 38944 1676 38956
rect 1631 38916 1676 38944
rect 1670 38904 1676 38916
rect 1728 38904 1734 38956
rect 14734 38944 14740 38956
rect 14695 38916 14740 38944
rect 14734 38904 14740 38916
rect 14792 38904 14798 38956
rect 14918 38944 14924 38956
rect 14879 38916 14924 38944
rect 14918 38904 14924 38916
rect 14976 38904 14982 38956
rect 16022 38944 16028 38956
rect 15028 38916 16028 38944
rect 14826 38836 14832 38888
rect 14884 38876 14890 38888
rect 15028 38876 15056 38916
rect 16022 38904 16028 38916
rect 16080 38904 16086 38956
rect 16117 38947 16175 38953
rect 16117 38913 16129 38947
rect 16163 38944 16175 38947
rect 16942 38944 16948 38956
rect 16163 38916 16948 38944
rect 16163 38913 16175 38916
rect 16117 38907 16175 38913
rect 16942 38904 16948 38916
rect 17000 38904 17006 38956
rect 18325 38947 18383 38953
rect 18325 38913 18337 38947
rect 18371 38913 18383 38947
rect 18874 38944 18880 38956
rect 18325 38907 18383 38913
rect 18432 38916 18880 38944
rect 15933 38879 15991 38885
rect 15933 38876 15945 38879
rect 14884 38848 15056 38876
rect 15120 38848 15945 38876
rect 14884 38836 14890 38848
rect 1854 38808 1860 38820
rect 1815 38780 1860 38808
rect 1854 38768 1860 38780
rect 1912 38768 1918 38820
rect 15010 38700 15016 38752
rect 15068 38740 15074 38752
rect 15120 38749 15148 38848
rect 15933 38845 15945 38848
rect 15979 38845 15991 38879
rect 15933 38839 15991 38845
rect 16209 38879 16267 38885
rect 16209 38845 16221 38879
rect 16255 38876 16267 38879
rect 18046 38876 18052 38888
rect 16255 38848 18052 38876
rect 16255 38845 16267 38848
rect 16209 38839 16267 38845
rect 18046 38836 18052 38848
rect 18104 38836 18110 38888
rect 18340 38808 18368 38907
rect 18432 38885 18460 38916
rect 18874 38904 18880 38916
rect 18932 38944 18938 38956
rect 20533 38947 20591 38953
rect 20533 38944 20545 38947
rect 18932 38916 20545 38944
rect 18932 38904 18938 38916
rect 20533 38913 20545 38916
rect 20579 38913 20591 38947
rect 20533 38907 20591 38913
rect 22005 38947 22063 38953
rect 22005 38913 22017 38947
rect 22051 38913 22063 38947
rect 22005 38907 22063 38913
rect 22097 38947 22155 38953
rect 22097 38913 22109 38947
rect 22143 38944 22155 38947
rect 22186 38944 22192 38956
rect 22143 38916 22192 38944
rect 22143 38913 22155 38916
rect 22097 38907 22155 38913
rect 18417 38879 18475 38885
rect 18417 38845 18429 38879
rect 18463 38845 18475 38879
rect 20622 38876 20628 38888
rect 20583 38848 20628 38876
rect 18417 38839 18475 38845
rect 20622 38836 20628 38848
rect 20680 38836 20686 38888
rect 20809 38879 20867 38885
rect 20809 38845 20821 38879
rect 20855 38876 20867 38879
rect 21726 38876 21732 38888
rect 20855 38848 21732 38876
rect 20855 38845 20867 38848
rect 20809 38839 20867 38845
rect 21726 38836 21732 38848
rect 21784 38876 21790 38888
rect 22020 38876 22048 38907
rect 22186 38904 22192 38916
rect 22244 38904 22250 38956
rect 22278 38904 22284 38956
rect 22336 38944 22342 38956
rect 23566 38944 23572 38956
rect 22336 38916 22381 38944
rect 23527 38916 23572 38944
rect 22336 38904 22342 38916
rect 23566 38904 23572 38916
rect 23624 38904 23630 38956
rect 24394 38944 24400 38956
rect 24355 38916 24400 38944
rect 24394 38904 24400 38916
rect 24452 38904 24458 38956
rect 24765 38947 24823 38953
rect 24765 38913 24777 38947
rect 24811 38944 24823 38947
rect 28442 38944 28448 38956
rect 24811 38916 28448 38944
rect 24811 38913 24823 38916
rect 24765 38907 24823 38913
rect 23474 38876 23480 38888
rect 21784 38848 22048 38876
rect 23435 38848 23480 38876
rect 21784 38836 21790 38848
rect 23474 38836 23480 38848
rect 23532 38836 23538 38888
rect 23845 38879 23903 38885
rect 23845 38845 23857 38879
rect 23891 38845 23903 38879
rect 23845 38839 23903 38845
rect 19242 38808 19248 38820
rect 18340 38780 19248 38808
rect 19242 38768 19248 38780
rect 19300 38768 19306 38820
rect 22465 38811 22523 38817
rect 22465 38777 22477 38811
rect 22511 38808 22523 38811
rect 23566 38808 23572 38820
rect 22511 38780 23572 38808
rect 22511 38777 22523 38780
rect 22465 38771 22523 38777
rect 23566 38768 23572 38780
rect 23624 38808 23630 38820
rect 23750 38808 23756 38820
rect 23624 38780 23756 38808
rect 23624 38768 23630 38780
rect 23750 38768 23756 38780
rect 23808 38768 23814 38820
rect 23860 38808 23888 38839
rect 23934 38836 23940 38888
rect 23992 38876 23998 38888
rect 24486 38876 24492 38888
rect 23992 38848 24492 38876
rect 23992 38836 23998 38848
rect 24486 38836 24492 38848
rect 24544 38836 24550 38888
rect 24780 38808 24808 38907
rect 28442 38904 28448 38916
rect 28500 38904 28506 38956
rect 35710 38904 35716 38956
rect 35768 38944 35774 38956
rect 47578 38944 47584 38956
rect 35768 38916 47584 38944
rect 35768 38904 35774 38916
rect 47578 38904 47584 38916
rect 47636 38944 47642 38956
rect 47765 38947 47823 38953
rect 47765 38944 47777 38947
rect 47636 38916 47777 38944
rect 47636 38904 47642 38916
rect 47765 38913 47777 38916
rect 47811 38913 47823 38947
rect 47765 38907 47823 38913
rect 23860 38780 24808 38808
rect 23952 38752 23980 38780
rect 15105 38743 15163 38749
rect 15105 38740 15117 38743
rect 15068 38712 15117 38740
rect 15068 38700 15074 38712
rect 15105 38709 15117 38712
rect 15151 38709 15163 38743
rect 15105 38703 15163 38709
rect 15749 38743 15807 38749
rect 15749 38709 15761 38743
rect 15795 38740 15807 38743
rect 15930 38740 15936 38752
rect 15795 38712 15936 38740
rect 15795 38709 15807 38712
rect 15749 38703 15807 38709
rect 15930 38700 15936 38712
rect 15988 38700 15994 38752
rect 17954 38740 17960 38752
rect 17915 38712 17960 38740
rect 17954 38700 17960 38712
rect 18012 38700 18018 38752
rect 23293 38743 23351 38749
rect 23293 38709 23305 38743
rect 23339 38740 23351 38743
rect 23382 38740 23388 38752
rect 23339 38712 23388 38740
rect 23339 38709 23351 38712
rect 23293 38703 23351 38709
rect 23382 38700 23388 38712
rect 23440 38700 23446 38752
rect 23934 38700 23940 38752
rect 23992 38700 23998 38752
rect 24854 38700 24860 38752
rect 24912 38740 24918 38752
rect 24949 38743 25007 38749
rect 24949 38740 24961 38743
rect 24912 38712 24961 38740
rect 24912 38700 24918 38712
rect 24949 38709 24961 38712
rect 24995 38709 25007 38743
rect 24949 38703 25007 38709
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 13541 38539 13599 38545
rect 13541 38505 13553 38539
rect 13587 38536 13599 38539
rect 14274 38536 14280 38548
rect 13587 38508 14280 38536
rect 13587 38505 13599 38508
rect 13541 38499 13599 38505
rect 14274 38496 14280 38508
rect 14332 38536 14338 38548
rect 14918 38536 14924 38548
rect 14332 38508 14924 38536
rect 14332 38496 14338 38508
rect 14918 38496 14924 38508
rect 14976 38496 14982 38548
rect 16942 38536 16948 38548
rect 16903 38508 16948 38536
rect 16942 38496 16948 38508
rect 17000 38496 17006 38548
rect 18874 38536 18880 38548
rect 18835 38508 18880 38536
rect 18874 38496 18880 38508
rect 18932 38496 18938 38548
rect 22281 38539 22339 38545
rect 22281 38505 22293 38539
rect 22327 38536 22339 38539
rect 22370 38536 22376 38548
rect 22327 38508 22376 38536
rect 22327 38505 22339 38508
rect 22281 38499 22339 38505
rect 22370 38496 22376 38508
rect 22428 38496 22434 38548
rect 23293 38539 23351 38545
rect 23293 38505 23305 38539
rect 23339 38536 23351 38539
rect 23474 38536 23480 38548
rect 23339 38508 23480 38536
rect 23339 38505 23351 38508
rect 23293 38499 23351 38505
rect 23474 38496 23480 38508
rect 23532 38496 23538 38548
rect 25590 38496 25596 38548
rect 25648 38536 25654 38548
rect 25961 38539 26019 38545
rect 25961 38536 25973 38539
rect 25648 38508 25973 38536
rect 25648 38496 25654 38508
rect 25961 38505 25973 38508
rect 26007 38505 26019 38539
rect 25961 38499 26019 38505
rect 15102 38468 15108 38480
rect 15063 38440 15108 38468
rect 15102 38428 15108 38440
rect 15160 38428 15166 38480
rect 14752 38372 15608 38400
rect 4798 38292 4804 38344
rect 4856 38332 4862 38344
rect 6733 38335 6791 38341
rect 6733 38332 6745 38335
rect 4856 38304 6745 38332
rect 4856 38292 4862 38304
rect 6733 38301 6745 38304
rect 6779 38332 6791 38335
rect 8478 38332 8484 38344
rect 6779 38304 8484 38332
rect 6779 38301 6791 38304
rect 6733 38295 6791 38301
rect 8478 38292 8484 38304
rect 8536 38292 8542 38344
rect 12161 38335 12219 38341
rect 12161 38301 12173 38335
rect 12207 38332 12219 38335
rect 12894 38332 12900 38344
rect 12207 38304 12900 38332
rect 12207 38301 12219 38304
rect 12161 38295 12219 38301
rect 12894 38292 12900 38304
rect 12952 38332 12958 38344
rect 14752 38332 14780 38372
rect 12952 38304 14780 38332
rect 14829 38335 14887 38341
rect 12952 38292 12958 38304
rect 14829 38301 14841 38335
rect 14875 38332 14887 38335
rect 15010 38332 15016 38344
rect 14875 38304 15016 38332
rect 14875 38301 14887 38304
rect 14829 38295 14887 38301
rect 15010 38292 15016 38304
rect 15068 38292 15074 38344
rect 15580 38341 15608 38372
rect 15565 38335 15623 38341
rect 15565 38301 15577 38335
rect 15611 38332 15623 38335
rect 15654 38332 15660 38344
rect 15611 38304 15660 38332
rect 15611 38301 15623 38304
rect 15565 38295 15623 38301
rect 15654 38292 15660 38304
rect 15712 38332 15718 38344
rect 17497 38335 17555 38341
rect 17497 38332 17509 38335
rect 15712 38304 17509 38332
rect 15712 38292 15718 38304
rect 17497 38301 17509 38304
rect 17543 38301 17555 38335
rect 17497 38295 17555 38301
rect 22278 38292 22284 38344
rect 22336 38332 22342 38344
rect 22465 38335 22523 38341
rect 22465 38332 22477 38335
rect 22336 38304 22477 38332
rect 22336 38292 22342 38304
rect 22465 38301 22477 38304
rect 22511 38301 22523 38335
rect 23566 38332 23572 38344
rect 23527 38304 23572 38332
rect 22465 38295 22523 38301
rect 23566 38292 23572 38304
rect 23624 38292 23630 38344
rect 24578 38332 24584 38344
rect 24539 38304 24584 38332
rect 24578 38292 24584 38304
rect 24636 38292 24642 38344
rect 24854 38341 24860 38344
rect 24848 38332 24860 38341
rect 24815 38304 24860 38332
rect 24848 38295 24860 38304
rect 24854 38292 24860 38295
rect 24912 38292 24918 38344
rect 47673 38335 47731 38341
rect 47673 38301 47685 38335
rect 47719 38332 47731 38335
rect 48314 38332 48320 38344
rect 47719 38304 48320 38332
rect 47719 38301 47731 38304
rect 47673 38295 47731 38301
rect 48314 38292 48320 38304
rect 48372 38292 48378 38344
rect 12428 38267 12486 38273
rect 12428 38233 12440 38267
rect 12474 38264 12486 38267
rect 12802 38264 12808 38276
rect 12474 38236 12808 38264
rect 12474 38233 12486 38236
rect 12428 38227 12486 38233
rect 12802 38224 12808 38236
rect 12860 38224 12866 38276
rect 15838 38273 15844 38276
rect 15105 38267 15163 38273
rect 15105 38233 15117 38267
rect 15151 38233 15163 38267
rect 15105 38227 15163 38233
rect 15832 38227 15844 38273
rect 15896 38264 15902 38276
rect 17764 38267 17822 38273
rect 15896 38236 15932 38264
rect 6546 38196 6552 38208
rect 6507 38168 6552 38196
rect 6546 38156 6552 38168
rect 6604 38156 6610 38208
rect 14826 38156 14832 38208
rect 14884 38196 14890 38208
rect 14921 38199 14979 38205
rect 14921 38196 14933 38199
rect 14884 38168 14933 38196
rect 14884 38156 14890 38168
rect 14921 38165 14933 38168
rect 14967 38165 14979 38199
rect 15120 38196 15148 38227
rect 15838 38224 15844 38227
rect 15896 38224 15902 38236
rect 17764 38233 17776 38267
rect 17810 38264 17822 38267
rect 18690 38264 18696 38276
rect 17810 38236 18696 38264
rect 17810 38233 17822 38236
rect 17764 38227 17822 38233
rect 18690 38224 18696 38236
rect 18748 38224 18754 38276
rect 22649 38267 22707 38273
rect 22649 38233 22661 38267
rect 22695 38264 22707 38267
rect 23293 38267 23351 38273
rect 23293 38264 23305 38267
rect 22695 38236 23305 38264
rect 22695 38233 22707 38236
rect 22649 38227 22707 38233
rect 23293 38233 23305 38236
rect 23339 38264 23351 38267
rect 23658 38264 23664 38276
rect 23339 38236 23664 38264
rect 23339 38233 23351 38236
rect 23293 38227 23351 38233
rect 23658 38224 23664 38236
rect 23716 38224 23722 38276
rect 16942 38196 16948 38208
rect 15120 38168 16948 38196
rect 14921 38159 14979 38165
rect 16942 38156 16948 38168
rect 17000 38156 17006 38208
rect 23477 38199 23535 38205
rect 23477 38165 23489 38199
rect 23523 38196 23535 38199
rect 23842 38196 23848 38208
rect 23523 38168 23848 38196
rect 23523 38165 23535 38168
rect 23477 38159 23535 38165
rect 23842 38156 23848 38168
rect 23900 38156 23906 38208
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 5997 37995 6055 38001
rect 5997 37961 6009 37995
rect 6043 37961 6055 37995
rect 5997 37955 6055 37961
rect 6012 37924 6040 37955
rect 12802 37952 12808 38004
rect 12860 37992 12866 38004
rect 12897 37995 12955 38001
rect 12897 37992 12909 37995
rect 12860 37964 12909 37992
rect 12860 37952 12866 37964
rect 12897 37961 12909 37964
rect 12943 37961 12955 37995
rect 12897 37955 12955 37961
rect 13633 37995 13691 38001
rect 13633 37961 13645 37995
rect 13679 37961 13691 37995
rect 13633 37955 13691 37961
rect 14001 37995 14059 38001
rect 14001 37961 14013 37995
rect 14047 37992 14059 37995
rect 14829 37995 14887 38001
rect 14829 37992 14841 37995
rect 14047 37964 14841 37992
rect 14047 37961 14059 37964
rect 14001 37955 14059 37961
rect 14829 37961 14841 37964
rect 14875 37961 14887 37995
rect 15657 37995 15715 38001
rect 14829 37955 14887 37961
rect 14936 37964 15240 37992
rect 6794 37927 6852 37933
rect 6794 37924 6806 37927
rect 6012 37896 6806 37924
rect 6794 37893 6806 37896
rect 6840 37893 6852 37927
rect 6794 37887 6852 37893
rect 4798 37856 4804 37868
rect 4759 37828 4804 37856
rect 4798 37816 4804 37828
rect 4856 37816 4862 37868
rect 5810 37856 5816 37868
rect 5771 37828 5816 37856
rect 5810 37816 5816 37828
rect 5868 37816 5874 37868
rect 6546 37856 6552 37868
rect 6507 37828 6552 37856
rect 6546 37816 6552 37828
rect 6604 37816 6610 37868
rect 8110 37816 8116 37868
rect 8168 37856 8174 37868
rect 8478 37856 8484 37868
rect 8168 37828 8484 37856
rect 8168 37816 8174 37828
rect 8478 37816 8484 37828
rect 8536 37816 8542 37868
rect 13081 37859 13139 37865
rect 13081 37825 13093 37859
rect 13127 37856 13139 37859
rect 13648 37856 13676 37955
rect 14734 37884 14740 37936
rect 14792 37924 14798 37936
rect 14936 37924 14964 37964
rect 15212 37933 15240 37964
rect 15657 37961 15669 37995
rect 15703 37992 15715 37995
rect 15838 37992 15844 38004
rect 15703 37964 15844 37992
rect 15703 37961 15715 37964
rect 15657 37955 15715 37961
rect 15838 37952 15844 37964
rect 15896 37952 15902 38004
rect 18690 37992 18696 38004
rect 18651 37964 18696 37992
rect 18690 37952 18696 37964
rect 18748 37952 18754 38004
rect 24486 37992 24492 38004
rect 24447 37964 24492 37992
rect 24486 37952 24492 37964
rect 24544 37952 24550 38004
rect 14792 37896 14964 37924
rect 14997 37927 15055 37933
rect 14792 37884 14798 37896
rect 14997 37893 15009 37927
rect 15043 37924 15055 37927
rect 15197 37927 15255 37933
rect 15043 37893 15056 37924
rect 14997 37887 15056 37893
rect 15197 37893 15209 37927
rect 15243 37893 15255 37927
rect 15197 37887 15255 37893
rect 16301 37927 16359 37933
rect 16301 37893 16313 37927
rect 16347 37924 16359 37927
rect 16942 37924 16948 37936
rect 16347 37896 16948 37924
rect 16347 37893 16359 37896
rect 16301 37887 16359 37893
rect 13127 37828 13676 37856
rect 13127 37825 13139 37828
rect 13081 37819 13139 37825
rect 14826 37816 14832 37868
rect 14884 37856 14890 37868
rect 15028 37856 15056 37887
rect 16942 37884 16948 37896
rect 17000 37884 17006 37936
rect 17589 37927 17647 37933
rect 17589 37893 17601 37927
rect 17635 37924 17647 37927
rect 18325 37927 18383 37933
rect 18325 37924 18337 37927
rect 17635 37896 18337 37924
rect 17635 37893 17647 37896
rect 17589 37887 17647 37893
rect 18325 37893 18337 37896
rect 18371 37893 18383 37927
rect 18325 37887 18383 37893
rect 18417 37927 18475 37933
rect 18417 37893 18429 37927
rect 18463 37924 18475 37927
rect 18874 37924 18880 37936
rect 18463 37896 18880 37924
rect 18463 37893 18475 37896
rect 18417 37887 18475 37893
rect 18874 37884 18880 37896
rect 18932 37884 18938 37936
rect 18966 37884 18972 37936
rect 19024 37924 19030 37936
rect 24578 37924 24584 37936
rect 19024 37896 20484 37924
rect 19024 37884 19030 37896
rect 14884 37828 15056 37856
rect 14884 37816 14890 37828
rect 15102 37816 15108 37868
rect 15160 37856 15166 37868
rect 15841 37859 15899 37865
rect 15841 37856 15853 37859
rect 15160 37828 15853 37856
rect 15160 37816 15166 37828
rect 15841 37825 15853 37828
rect 15887 37825 15899 37859
rect 15841 37819 15899 37825
rect 15930 37816 15936 37868
rect 15988 37856 15994 37868
rect 17497 37859 17555 37865
rect 15988 37828 16033 37856
rect 15988 37816 15994 37828
rect 17497 37825 17509 37859
rect 17543 37825 17555 37859
rect 17497 37819 17555 37825
rect 17681 37859 17739 37865
rect 17681 37825 17693 37859
rect 17727 37856 17739 37859
rect 17954 37856 17960 37868
rect 17727 37828 17960 37856
rect 17727 37825 17739 37828
rect 17681 37819 17739 37825
rect 13814 37748 13820 37800
rect 13872 37788 13878 37800
rect 14093 37791 14151 37797
rect 14093 37788 14105 37791
rect 13872 37760 14105 37788
rect 13872 37748 13878 37760
rect 14093 37757 14105 37760
rect 14139 37757 14151 37791
rect 14274 37788 14280 37800
rect 14235 37760 14280 37788
rect 14093 37751 14151 37757
rect 14274 37748 14280 37760
rect 14332 37748 14338 37800
rect 16209 37791 16267 37797
rect 16209 37757 16221 37791
rect 16255 37757 16267 37791
rect 17512 37788 17540 37819
rect 17954 37816 17960 37828
rect 18012 37816 18018 37868
rect 18141 37859 18199 37865
rect 18141 37825 18153 37859
rect 18187 37856 18199 37859
rect 18230 37856 18236 37868
rect 18187 37828 18236 37856
rect 18187 37825 18199 37828
rect 18141 37819 18199 37825
rect 18230 37816 18236 37828
rect 18288 37816 18294 37868
rect 18509 37859 18567 37865
rect 18509 37825 18521 37859
rect 18555 37856 18567 37859
rect 18555 37828 18736 37856
rect 18555 37825 18567 37828
rect 18509 37819 18567 37825
rect 18598 37788 18604 37800
rect 17512 37760 18604 37788
rect 16209 37751 16267 37757
rect 16224 37720 16252 37751
rect 18598 37748 18604 37760
rect 18656 37748 18662 37800
rect 18138 37720 18144 37732
rect 16224 37692 18144 37720
rect 18138 37680 18144 37692
rect 18196 37720 18202 37732
rect 18708 37720 18736 37828
rect 19242 37816 19248 37868
rect 19300 37856 19306 37868
rect 20456 37865 20484 37896
rect 23124 37896 24584 37924
rect 23124 37865 23152 37896
rect 24578 37884 24584 37896
rect 24636 37884 24642 37936
rect 23382 37865 23388 37868
rect 19797 37859 19855 37865
rect 19797 37856 19809 37859
rect 19300 37828 19809 37856
rect 19300 37816 19306 37828
rect 19797 37825 19809 37828
rect 19843 37825 19855 37859
rect 19797 37819 19855 37825
rect 20441 37859 20499 37865
rect 20441 37825 20453 37859
rect 20487 37825 20499 37859
rect 20441 37819 20499 37825
rect 23109 37859 23167 37865
rect 23109 37825 23121 37859
rect 23155 37825 23167 37859
rect 23376 37856 23388 37865
rect 23343 37828 23388 37856
rect 23109 37819 23167 37825
rect 23376 37819 23388 37828
rect 23382 37816 23388 37819
rect 23440 37816 23446 37868
rect 46934 37816 46940 37868
rect 46992 37856 46998 37868
rect 47765 37859 47823 37865
rect 47765 37856 47777 37859
rect 46992 37828 47777 37856
rect 46992 37816 46998 37828
rect 47765 37825 47777 37828
rect 47811 37856 47823 37859
rect 48038 37856 48044 37868
rect 47811 37828 48044 37856
rect 47811 37825 47823 37828
rect 47765 37819 47823 37825
rect 48038 37816 48044 37828
rect 48096 37816 48102 37868
rect 19889 37791 19947 37797
rect 19889 37757 19901 37791
rect 19935 37788 19947 37791
rect 20622 37788 20628 37800
rect 19935 37760 20628 37788
rect 19935 37757 19947 37760
rect 19889 37751 19947 37757
rect 20622 37748 20628 37760
rect 20680 37748 20686 37800
rect 20714 37720 20720 37732
rect 18196 37692 20720 37720
rect 18196 37680 18202 37692
rect 20714 37680 20720 37692
rect 20772 37680 20778 37732
rect 4798 37652 4804 37664
rect 4759 37624 4804 37652
rect 4798 37612 4804 37624
rect 4856 37612 4862 37664
rect 7926 37652 7932 37664
rect 7887 37624 7932 37652
rect 7926 37612 7932 37624
rect 7984 37612 7990 37664
rect 8478 37652 8484 37664
rect 8439 37624 8484 37652
rect 8478 37612 8484 37624
rect 8536 37612 8542 37664
rect 15013 37655 15071 37661
rect 15013 37621 15025 37655
rect 15059 37652 15071 37655
rect 15102 37652 15108 37664
rect 15059 37624 15108 37652
rect 15059 37621 15071 37624
rect 15013 37615 15071 37621
rect 15102 37612 15108 37624
rect 15160 37612 15166 37664
rect 19426 37612 19432 37664
rect 19484 37652 19490 37664
rect 19521 37655 19579 37661
rect 19521 37652 19533 37655
rect 19484 37624 19533 37652
rect 19484 37612 19490 37624
rect 19521 37621 19533 37624
rect 19567 37652 19579 37655
rect 19794 37652 19800 37664
rect 19567 37624 19800 37652
rect 19567 37621 19579 37624
rect 19521 37615 19579 37621
rect 19794 37612 19800 37624
rect 19852 37652 19858 37664
rect 20533 37655 20591 37661
rect 20533 37652 20545 37655
rect 19852 37624 20545 37652
rect 19852 37612 19858 37624
rect 20533 37621 20545 37624
rect 20579 37621 20591 37655
rect 20533 37615 20591 37621
rect 20901 37655 20959 37661
rect 20901 37621 20913 37655
rect 20947 37652 20959 37655
rect 22278 37652 22284 37664
rect 20947 37624 22284 37652
rect 20947 37621 20959 37624
rect 20901 37615 20959 37621
rect 22278 37612 22284 37624
rect 22336 37612 22342 37664
rect 47857 37655 47915 37661
rect 47857 37621 47869 37655
rect 47903 37652 47915 37655
rect 48130 37652 48136 37664
rect 47903 37624 48136 37652
rect 47903 37621 47915 37624
rect 47857 37615 47915 37621
rect 48130 37612 48136 37624
rect 48188 37612 48194 37664
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 6181 37451 6239 37457
rect 6181 37417 6193 37451
rect 6227 37448 6239 37451
rect 6917 37451 6975 37457
rect 6917 37448 6929 37451
rect 6227 37420 6929 37448
rect 6227 37417 6239 37420
rect 6181 37411 6239 37417
rect 6917 37417 6929 37420
rect 6963 37417 6975 37451
rect 7926 37448 7932 37460
rect 7887 37420 7932 37448
rect 6917 37411 6975 37417
rect 7926 37408 7932 37420
rect 7984 37408 7990 37460
rect 18230 37448 18236 37460
rect 18191 37420 18236 37448
rect 18230 37408 18236 37420
rect 18288 37408 18294 37460
rect 20622 37448 20628 37460
rect 20583 37420 20628 37448
rect 20622 37408 20628 37420
rect 20680 37408 20686 37460
rect 5810 37340 5816 37392
rect 5868 37380 5874 37392
rect 6641 37383 6699 37389
rect 6641 37380 6653 37383
rect 5868 37352 6653 37380
rect 5868 37340 5874 37352
rect 6641 37349 6653 37352
rect 6687 37349 6699 37383
rect 6641 37343 6699 37349
rect 15933 37383 15991 37389
rect 15933 37349 15945 37383
rect 15979 37380 15991 37383
rect 16942 37380 16948 37392
rect 15979 37352 16948 37380
rect 15979 37349 15991 37352
rect 15933 37343 15991 37349
rect 16942 37340 16948 37352
rect 17000 37340 17006 37392
rect 1949 37315 2007 37321
rect 1949 37281 1961 37315
rect 1995 37312 2007 37315
rect 2682 37312 2688 37324
rect 1995 37284 2688 37312
rect 1995 37281 2007 37284
rect 1949 37275 2007 37281
rect 2682 37272 2688 37284
rect 2740 37272 2746 37324
rect 4798 37312 4804 37324
rect 4759 37284 4804 37312
rect 4798 37272 4804 37284
rect 4856 37272 4862 37324
rect 13725 37315 13783 37321
rect 13725 37281 13737 37315
rect 13771 37312 13783 37315
rect 13814 37312 13820 37324
rect 13771 37284 13820 37312
rect 13771 37281 13783 37284
rect 13725 37275 13783 37281
rect 13814 37272 13820 37284
rect 13872 37272 13878 37324
rect 14550 37272 14556 37324
rect 14608 37312 14614 37324
rect 15381 37315 15439 37321
rect 15381 37312 15393 37315
rect 14608 37284 15393 37312
rect 14608 37272 14614 37284
rect 15381 37281 15393 37284
rect 15427 37281 15439 37315
rect 15381 37275 15439 37281
rect 17954 37272 17960 37324
rect 18012 37312 18018 37324
rect 18693 37315 18751 37321
rect 18693 37312 18705 37315
rect 18012 37284 18705 37312
rect 18012 37272 18018 37284
rect 18693 37281 18705 37284
rect 18739 37312 18751 37315
rect 18966 37312 18972 37324
rect 18739 37284 18972 37312
rect 18739 37281 18751 37284
rect 18693 37275 18751 37281
rect 18966 37272 18972 37284
rect 19024 37272 19030 37324
rect 20073 37315 20131 37321
rect 20073 37281 20085 37315
rect 20119 37312 20131 37315
rect 20640 37312 20668 37408
rect 27893 37383 27951 37389
rect 27893 37349 27905 37383
rect 27939 37349 27951 37383
rect 27893 37343 27951 37349
rect 20119 37284 20668 37312
rect 20119 37281 20131 37284
rect 20073 37275 20131 37281
rect 4157 37247 4215 37253
rect 4157 37213 4169 37247
rect 4203 37244 4215 37247
rect 4890 37244 4896 37256
rect 4203 37216 4896 37244
rect 4203 37213 4215 37216
rect 4157 37207 4215 37213
rect 4890 37204 4896 37216
rect 4948 37204 4954 37256
rect 7098 37244 7104 37256
rect 7059 37216 7104 37244
rect 7098 37204 7104 37216
rect 7156 37244 7162 37256
rect 7653 37247 7711 37253
rect 7653 37244 7665 37247
rect 7156 37216 7665 37244
rect 7156 37204 7162 37216
rect 7653 37213 7665 37216
rect 7699 37213 7711 37247
rect 9309 37247 9367 37253
rect 9309 37244 9321 37247
rect 7653 37207 7711 37213
rect 8128 37216 9321 37244
rect 1670 37176 1676 37188
rect 1631 37148 1676 37176
rect 1670 37136 1676 37148
rect 1728 37136 1734 37188
rect 5046 37179 5104 37185
rect 5046 37176 5058 37179
rect 4356 37148 5058 37176
rect 4356 37117 4384 37148
rect 5046 37145 5058 37148
rect 5092 37145 5104 37179
rect 5046 37139 5104 37145
rect 8128 37117 8156 37216
rect 9309 37213 9321 37216
rect 9355 37213 9367 37247
rect 9309 37207 9367 37213
rect 12713 37247 12771 37253
rect 12713 37213 12725 37247
rect 12759 37244 12771 37247
rect 13357 37247 13415 37253
rect 13357 37244 13369 37247
rect 12759 37216 13369 37244
rect 12759 37213 12771 37216
rect 12713 37207 12771 37213
rect 13357 37213 13369 37216
rect 13403 37213 13415 37247
rect 13357 37207 13415 37213
rect 13541 37247 13599 37253
rect 13541 37213 13553 37247
rect 13587 37213 13599 37247
rect 13541 37207 13599 37213
rect 14645 37247 14703 37253
rect 14645 37213 14657 37247
rect 14691 37244 14703 37247
rect 14734 37244 14740 37256
rect 14691 37216 14740 37244
rect 14691 37213 14703 37216
rect 14645 37207 14703 37213
rect 13556 37176 13584 37207
rect 14734 37204 14740 37216
rect 14792 37204 14798 37256
rect 14918 37244 14924 37256
rect 14879 37216 14924 37244
rect 14918 37204 14924 37216
rect 14976 37204 14982 37256
rect 15010 37204 15016 37256
rect 15068 37244 15074 37256
rect 15565 37247 15623 37253
rect 15565 37244 15577 37247
rect 15068 37216 15577 37244
rect 15068 37204 15074 37216
rect 15565 37213 15577 37216
rect 15611 37213 15623 37247
rect 15565 37207 15623 37213
rect 18417 37247 18475 37253
rect 18417 37213 18429 37247
rect 18463 37213 18475 37247
rect 18598 37244 18604 37256
rect 18559 37216 18604 37244
rect 18417 37207 18475 37213
rect 14461 37179 14519 37185
rect 14461 37176 14473 37179
rect 13556 37148 14473 37176
rect 14461 37145 14473 37148
rect 14507 37145 14519 37179
rect 14461 37139 14519 37145
rect 14829 37179 14887 37185
rect 14829 37145 14841 37179
rect 14875 37176 14887 37179
rect 15102 37176 15108 37188
rect 14875 37148 15108 37176
rect 14875 37145 14887 37148
rect 14829 37139 14887 37145
rect 15102 37136 15108 37148
rect 15160 37176 15166 37188
rect 15749 37179 15807 37185
rect 15749 37176 15761 37179
rect 15160 37148 15761 37176
rect 15160 37136 15166 37148
rect 15749 37145 15761 37148
rect 15795 37176 15807 37179
rect 17034 37176 17040 37188
rect 15795 37148 17040 37176
rect 15795 37145 15807 37148
rect 15749 37139 15807 37145
rect 17034 37136 17040 37148
rect 17092 37176 17098 37188
rect 18432 37176 18460 37207
rect 18598 37204 18604 37216
rect 18656 37204 18662 37256
rect 19334 37204 19340 37256
rect 19392 37244 19398 37256
rect 19705 37247 19763 37253
rect 19705 37244 19717 37247
rect 19392 37216 19717 37244
rect 19392 37204 19398 37216
rect 19705 37213 19717 37216
rect 19751 37213 19763 37247
rect 19705 37207 19763 37213
rect 19794 37204 19800 37256
rect 19852 37244 19858 37256
rect 20165 37247 20223 37253
rect 19852 37216 19897 37244
rect 19852 37204 19858 37216
rect 20165 37213 20177 37247
rect 20211 37244 20223 37247
rect 20806 37244 20812 37256
rect 20211 37216 20812 37244
rect 20211 37213 20223 37216
rect 20165 37207 20223 37213
rect 20806 37204 20812 37216
rect 20864 37204 20870 37256
rect 22005 37247 22063 37253
rect 22005 37213 22017 37247
rect 22051 37244 22063 37247
rect 23842 37244 23848 37256
rect 22051 37216 23848 37244
rect 22051 37213 22063 37216
rect 22005 37207 22063 37213
rect 23842 37204 23848 37216
rect 23900 37244 23906 37256
rect 24578 37244 24584 37256
rect 23900 37216 24584 37244
rect 23900 37204 23906 37216
rect 24578 37204 24584 37216
rect 24636 37244 24642 37256
rect 27433 37247 27491 37253
rect 27433 37244 27445 37247
rect 24636 37216 27445 37244
rect 24636 37204 24642 37216
rect 27433 37213 27445 37216
rect 27479 37244 27491 37247
rect 27706 37244 27712 37256
rect 27479 37216 27712 37244
rect 27479 37213 27491 37216
rect 27433 37207 27491 37213
rect 27706 37204 27712 37216
rect 27764 37204 27770 37256
rect 17092 37148 19656 37176
rect 17092 37136 17098 37148
rect 4341 37111 4399 37117
rect 4341 37077 4353 37111
rect 4387 37077 4399 37111
rect 4341 37071 4399 37077
rect 8113 37111 8171 37117
rect 8113 37077 8125 37111
rect 8159 37077 8171 37111
rect 9122 37108 9128 37120
rect 9083 37080 9128 37108
rect 8113 37071 8171 37077
rect 9122 37068 9128 37080
rect 9180 37068 9186 37120
rect 12897 37111 12955 37117
rect 12897 37077 12909 37111
rect 12943 37108 12955 37111
rect 13170 37108 13176 37120
rect 12943 37080 13176 37108
rect 12943 37077 12955 37080
rect 12897 37071 12955 37077
rect 13170 37068 13176 37080
rect 13228 37068 13234 37120
rect 14918 37068 14924 37120
rect 14976 37108 14982 37120
rect 15657 37111 15715 37117
rect 15657 37108 15669 37111
rect 14976 37080 15669 37108
rect 14976 37068 14982 37080
rect 15657 37077 15669 37080
rect 15703 37077 15715 37111
rect 15657 37071 15715 37077
rect 18598 37068 18604 37120
rect 18656 37108 18662 37120
rect 19521 37111 19579 37117
rect 19521 37108 19533 37111
rect 18656 37080 19533 37108
rect 18656 37068 18662 37080
rect 19521 37077 19533 37080
rect 19567 37077 19579 37111
rect 19628 37108 19656 37148
rect 20898 37136 20904 37188
rect 20956 37176 20962 37188
rect 21738 37179 21796 37185
rect 21738 37176 21750 37179
rect 20956 37148 21750 37176
rect 20956 37136 20962 37148
rect 21738 37145 21750 37148
rect 21784 37145 21796 37179
rect 21738 37139 21796 37145
rect 22462 37136 22468 37188
rect 22520 37176 22526 37188
rect 23934 37176 23940 37188
rect 22520 37148 23940 37176
rect 22520 37136 22526 37148
rect 23934 37136 23940 37148
rect 23992 37136 23998 37188
rect 27188 37179 27246 37185
rect 27188 37145 27200 37179
rect 27234 37176 27246 37179
rect 27908 37176 27936 37343
rect 28442 37312 28448 37324
rect 28403 37284 28448 37312
rect 28442 37272 28448 37284
rect 28500 37272 28506 37324
rect 48130 37312 48136 37324
rect 48091 37284 48136 37312
rect 48130 37272 48136 37284
rect 48188 37272 48194 37324
rect 28074 37244 28080 37256
rect 28035 37216 28080 37244
rect 28074 37204 28080 37216
rect 28132 37204 28138 37256
rect 28166 37204 28172 37256
rect 28224 37244 28230 37256
rect 46474 37244 46480 37256
rect 28224 37216 28269 37244
rect 46435 37216 46480 37244
rect 28224 37204 28230 37216
rect 46474 37204 46480 37216
rect 46532 37204 46538 37256
rect 48314 37204 48320 37256
rect 48372 37244 48378 37256
rect 48372 37216 48417 37244
rect 48372 37204 48378 37216
rect 27234 37148 27936 37176
rect 28537 37179 28595 37185
rect 27234 37145 27246 37148
rect 27188 37139 27246 37145
rect 28537 37145 28549 37179
rect 28583 37145 28595 37179
rect 28537 37139 28595 37145
rect 24762 37108 24768 37120
rect 19628 37080 24768 37108
rect 19521 37071 19579 37077
rect 24762 37068 24768 37080
rect 24820 37068 24826 37120
rect 26050 37108 26056 37120
rect 25963 37080 26056 37108
rect 26050 37068 26056 37080
rect 26108 37108 26114 37120
rect 28552 37108 28580 37139
rect 26108 37080 28580 37108
rect 26108 37068 26114 37080
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 13814 36864 13820 36916
rect 13872 36904 13878 36916
rect 15565 36907 15623 36913
rect 15565 36904 15577 36907
rect 13872 36876 15577 36904
rect 13872 36864 13878 36876
rect 15565 36873 15577 36876
rect 15611 36873 15623 36907
rect 20898 36904 20904 36916
rect 20859 36876 20904 36904
rect 15565 36867 15623 36873
rect 20898 36864 20904 36876
rect 20956 36864 20962 36916
rect 22186 36864 22192 36916
rect 22244 36904 22250 36916
rect 22465 36907 22523 36913
rect 22465 36904 22477 36907
rect 22244 36876 22477 36904
rect 22244 36864 22250 36876
rect 22465 36873 22477 36876
rect 22511 36873 22523 36907
rect 22465 36867 22523 36873
rect 25501 36907 25559 36913
rect 25501 36873 25513 36907
rect 25547 36904 25559 36907
rect 28166 36904 28172 36916
rect 25547 36876 28172 36904
rect 25547 36873 25559 36876
rect 25501 36867 25559 36873
rect 28166 36864 28172 36876
rect 28224 36864 28230 36916
rect 8104 36839 8162 36845
rect 8104 36805 8116 36839
rect 8150 36836 8162 36839
rect 9122 36836 9128 36848
rect 8150 36808 9128 36836
rect 8150 36805 8162 36808
rect 8104 36799 8162 36805
rect 9122 36796 9128 36808
rect 9180 36796 9186 36848
rect 13170 36845 13176 36848
rect 13164 36836 13176 36845
rect 13131 36808 13176 36836
rect 13164 36799 13176 36808
rect 13170 36796 13176 36799
rect 13228 36796 13234 36848
rect 14734 36796 14740 36848
rect 14792 36836 14798 36848
rect 15381 36839 15439 36845
rect 15381 36836 15393 36839
rect 14792 36808 15393 36836
rect 14792 36796 14798 36808
rect 15381 36805 15393 36808
rect 15427 36805 15439 36839
rect 20622 36836 20628 36848
rect 20583 36808 20628 36836
rect 15381 36799 15439 36805
rect 20622 36796 20628 36808
rect 20680 36796 20686 36848
rect 21726 36796 21732 36848
rect 21784 36836 21790 36848
rect 22097 36839 22155 36845
rect 22097 36836 22109 36839
rect 21784 36808 22109 36836
rect 21784 36796 21790 36808
rect 22097 36805 22109 36808
rect 22143 36805 22155 36839
rect 22097 36799 22155 36805
rect 24765 36839 24823 36845
rect 24765 36805 24777 36839
rect 24811 36836 24823 36839
rect 24811 36808 25636 36836
rect 24811 36805 24823 36808
rect 24765 36799 24823 36805
rect 25608 36780 25636 36808
rect 4516 36771 4574 36777
rect 4516 36737 4528 36771
rect 4562 36768 4574 36771
rect 5994 36768 6000 36780
rect 4562 36740 6000 36768
rect 4562 36737 4574 36740
rect 4516 36731 4574 36737
rect 5994 36728 6000 36740
rect 6052 36728 6058 36780
rect 7837 36771 7895 36777
rect 7837 36737 7849 36771
rect 7883 36768 7895 36771
rect 8478 36768 8484 36780
rect 7883 36740 8484 36768
rect 7883 36737 7895 36740
rect 7837 36731 7895 36737
rect 8478 36728 8484 36740
rect 8536 36728 8542 36780
rect 12894 36768 12900 36780
rect 12855 36740 12900 36768
rect 12894 36728 12900 36740
rect 12952 36728 12958 36780
rect 14918 36728 14924 36780
rect 14976 36768 14982 36780
rect 15289 36771 15347 36777
rect 15289 36768 15301 36771
rect 14976 36740 15301 36768
rect 14976 36728 14982 36740
rect 15289 36737 15301 36740
rect 15335 36737 15347 36771
rect 15289 36731 15347 36737
rect 15657 36771 15715 36777
rect 15657 36737 15669 36771
rect 15703 36768 15715 36771
rect 18230 36768 18236 36780
rect 15703 36740 18236 36768
rect 15703 36737 15715 36740
rect 15657 36731 15715 36737
rect 18230 36728 18236 36740
rect 18288 36728 18294 36780
rect 19334 36728 19340 36780
rect 19392 36768 19398 36780
rect 19518 36768 19524 36780
rect 19392 36740 19524 36768
rect 19392 36728 19398 36740
rect 19518 36728 19524 36740
rect 19576 36728 19582 36780
rect 20349 36771 20407 36777
rect 20349 36768 20361 36771
rect 19904 36740 20361 36768
rect 4062 36660 4068 36712
rect 4120 36700 4126 36712
rect 4249 36703 4307 36709
rect 4249 36700 4261 36703
rect 4120 36672 4261 36700
rect 4120 36660 4126 36672
rect 4249 36669 4261 36672
rect 4295 36669 4307 36703
rect 4249 36663 4307 36669
rect 15473 36703 15531 36709
rect 15473 36669 15485 36703
rect 15519 36700 15531 36703
rect 16482 36700 16488 36712
rect 15519 36672 16488 36700
rect 15519 36669 15531 36672
rect 15473 36663 15531 36669
rect 16482 36660 16488 36672
rect 16540 36660 16546 36712
rect 19426 36700 19432 36712
rect 19387 36672 19432 36700
rect 19426 36660 19432 36672
rect 19484 36660 19490 36712
rect 19904 36709 19932 36740
rect 20349 36737 20361 36740
rect 20395 36737 20407 36771
rect 20349 36731 20407 36737
rect 20533 36771 20591 36777
rect 20533 36737 20545 36771
rect 20579 36737 20591 36771
rect 20714 36768 20720 36780
rect 20675 36740 20720 36768
rect 20533 36731 20591 36737
rect 19889 36703 19947 36709
rect 19889 36669 19901 36703
rect 19935 36669 19947 36703
rect 19889 36663 19947 36669
rect 14277 36635 14335 36641
rect 14277 36601 14289 36635
rect 14323 36632 14335 36635
rect 14734 36632 14740 36644
rect 14323 36604 14740 36632
rect 14323 36601 14335 36604
rect 14277 36595 14335 36601
rect 14734 36592 14740 36604
rect 14792 36592 14798 36644
rect 17310 36592 17316 36644
rect 17368 36632 17374 36644
rect 20346 36632 20352 36644
rect 17368 36604 20352 36632
rect 17368 36592 17374 36604
rect 20346 36592 20352 36604
rect 20404 36632 20410 36644
rect 20548 36632 20576 36731
rect 20714 36728 20720 36740
rect 20772 36728 20778 36780
rect 21542 36728 21548 36780
rect 21600 36768 21606 36780
rect 22005 36771 22063 36777
rect 22005 36768 22017 36771
rect 21600 36740 22017 36768
rect 21600 36728 21606 36740
rect 22005 36737 22017 36740
rect 22051 36737 22063 36771
rect 22278 36768 22284 36780
rect 22239 36740 22284 36768
rect 22005 36731 22063 36737
rect 22278 36728 22284 36740
rect 22336 36728 22342 36780
rect 24673 36771 24731 36777
rect 24673 36737 24685 36771
rect 24719 36737 24731 36771
rect 24946 36768 24952 36780
rect 24907 36740 24952 36768
rect 24673 36731 24731 36737
rect 20732 36700 20760 36728
rect 22462 36700 22468 36712
rect 20732 36672 22468 36700
rect 22462 36660 22468 36672
rect 22520 36660 22526 36712
rect 24688 36700 24716 36731
rect 24946 36728 24952 36740
rect 25004 36728 25010 36780
rect 25409 36771 25467 36777
rect 25409 36737 25421 36771
rect 25455 36737 25467 36771
rect 25590 36768 25596 36780
rect 25551 36740 25596 36768
rect 25409 36731 25467 36737
rect 24854 36700 24860 36712
rect 24688 36672 24860 36700
rect 24854 36660 24860 36672
rect 24912 36660 24918 36712
rect 25424 36700 25452 36731
rect 25590 36728 25596 36740
rect 25648 36728 25654 36780
rect 27706 36768 27712 36780
rect 27667 36740 27712 36768
rect 27706 36728 27712 36740
rect 27764 36728 27770 36780
rect 27982 36777 27988 36780
rect 27976 36731 27988 36777
rect 28040 36768 28046 36780
rect 28040 36740 28076 36768
rect 27982 36728 27988 36731
rect 28040 36728 28046 36740
rect 25424 36672 25820 36700
rect 25682 36632 25688 36644
rect 20404 36604 25688 36632
rect 20404 36592 20410 36604
rect 25682 36592 25688 36604
rect 25740 36592 25746 36644
rect 5442 36524 5448 36576
rect 5500 36564 5506 36576
rect 5629 36567 5687 36573
rect 5629 36564 5641 36567
rect 5500 36536 5641 36564
rect 5500 36524 5506 36536
rect 5629 36533 5641 36536
rect 5675 36533 5687 36567
rect 9214 36564 9220 36576
rect 9175 36536 9220 36564
rect 5629 36527 5687 36533
rect 9214 36524 9220 36536
rect 9272 36524 9278 36576
rect 23934 36524 23940 36576
rect 23992 36564 23998 36576
rect 24673 36567 24731 36573
rect 24673 36564 24685 36567
rect 23992 36536 24685 36564
rect 23992 36524 23998 36536
rect 24673 36533 24685 36536
rect 24719 36533 24731 36567
rect 24673 36527 24731 36533
rect 24762 36524 24768 36576
rect 24820 36564 24826 36576
rect 25792 36564 25820 36672
rect 24820 36536 25820 36564
rect 24820 36524 24826 36536
rect 27706 36524 27712 36576
rect 27764 36564 27770 36576
rect 29089 36567 29147 36573
rect 29089 36564 29101 36567
rect 27764 36536 29101 36564
rect 27764 36524 27770 36536
rect 29089 36533 29101 36536
rect 29135 36533 29147 36567
rect 29089 36527 29147 36533
rect 47949 36567 48007 36573
rect 47949 36533 47961 36567
rect 47995 36564 48007 36567
rect 48314 36564 48320 36576
rect 47995 36536 48320 36564
rect 47995 36533 48007 36536
rect 47949 36527 48007 36533
rect 48314 36524 48320 36536
rect 48372 36524 48378 36576
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 4062 36320 4068 36372
rect 4120 36360 4126 36372
rect 4341 36363 4399 36369
rect 4341 36360 4353 36363
rect 4120 36332 4353 36360
rect 4120 36320 4126 36332
rect 4341 36329 4353 36332
rect 4387 36329 4399 36363
rect 4341 36323 4399 36329
rect 4890 36320 4896 36372
rect 4948 36360 4954 36372
rect 5077 36363 5135 36369
rect 5077 36360 5089 36363
rect 4948 36332 5089 36360
rect 4948 36320 4954 36332
rect 5077 36329 5089 36332
rect 5123 36329 5135 36363
rect 5442 36360 5448 36372
rect 5403 36332 5448 36360
rect 5077 36323 5135 36329
rect 5442 36320 5448 36332
rect 5500 36320 5506 36372
rect 5994 36360 6000 36372
rect 5955 36332 6000 36360
rect 5994 36320 6000 36332
rect 6052 36320 6058 36372
rect 9214 36360 9220 36372
rect 9175 36332 9220 36360
rect 9214 36320 9220 36332
rect 9272 36320 9278 36372
rect 17310 36360 17316 36372
rect 17271 36332 17316 36360
rect 17310 36320 17316 36332
rect 17368 36320 17374 36372
rect 19518 36320 19524 36372
rect 19576 36360 19582 36372
rect 21361 36363 21419 36369
rect 21361 36360 21373 36363
rect 19576 36332 21373 36360
rect 19576 36320 19582 36332
rect 21361 36329 21373 36332
rect 21407 36329 21419 36363
rect 21361 36323 21419 36329
rect 23937 36363 23995 36369
rect 23937 36329 23949 36363
rect 23983 36360 23995 36363
rect 24854 36360 24860 36372
rect 23983 36332 24860 36360
rect 23983 36329 23995 36332
rect 23937 36323 23995 36329
rect 24854 36320 24860 36332
rect 24912 36320 24918 36372
rect 26326 36320 26332 36372
rect 26384 36360 26390 36372
rect 26513 36363 26571 36369
rect 26513 36360 26525 36363
rect 26384 36332 26525 36360
rect 26384 36320 26390 36332
rect 26513 36329 26525 36332
rect 26559 36329 26571 36363
rect 26513 36323 26571 36329
rect 26697 36363 26755 36369
rect 26697 36329 26709 36363
rect 26743 36329 26755 36363
rect 27982 36360 27988 36372
rect 27943 36332 27988 36360
rect 26697 36323 26755 36329
rect 24872 36292 24900 36320
rect 26712 36292 26740 36323
rect 27982 36320 27988 36332
rect 28040 36320 28046 36372
rect 28074 36292 28080 36304
rect 24872 36264 25820 36292
rect 26712 36264 28080 36292
rect 4890 36184 4896 36236
rect 4948 36224 4954 36236
rect 5350 36224 5356 36236
rect 4948 36196 5356 36224
rect 4948 36184 4954 36196
rect 5350 36184 5356 36196
rect 5408 36184 5414 36236
rect 9585 36227 9643 36233
rect 9585 36193 9597 36227
rect 9631 36193 9643 36227
rect 21726 36224 21732 36236
rect 21687 36196 21732 36224
rect 9585 36187 9643 36193
rect 4525 36159 4583 36165
rect 4525 36125 4537 36159
rect 4571 36156 4583 36159
rect 4982 36156 4988 36168
rect 4571 36128 4988 36156
rect 4571 36125 4583 36128
rect 4525 36119 4583 36125
rect 4982 36116 4988 36128
rect 5040 36116 5046 36168
rect 5537 36159 5595 36165
rect 5537 36125 5549 36159
rect 5583 36125 5595 36159
rect 6178 36156 6184 36168
rect 6139 36128 6184 36156
rect 5537 36119 5595 36125
rect 5552 36088 5580 36119
rect 6178 36116 6184 36128
rect 6236 36116 6242 36168
rect 8110 36156 8116 36168
rect 8071 36128 8116 36156
rect 8110 36116 8116 36128
rect 8168 36116 8174 36168
rect 9125 36159 9183 36165
rect 9125 36156 9137 36159
rect 8220 36128 9137 36156
rect 7098 36088 7104 36100
rect 5552 36060 7104 36088
rect 7098 36048 7104 36060
rect 7156 36088 7162 36100
rect 8220 36088 8248 36128
rect 9125 36125 9137 36128
rect 9171 36156 9183 36159
rect 9214 36156 9220 36168
rect 9171 36128 9220 36156
rect 9171 36125 9183 36128
rect 9125 36119 9183 36125
rect 9214 36116 9220 36128
rect 9272 36116 9278 36168
rect 9600 36156 9628 36187
rect 21726 36184 21732 36196
rect 21784 36184 21790 36236
rect 23860 36196 24992 36224
rect 10229 36159 10287 36165
rect 10229 36156 10241 36159
rect 9600 36128 10241 36156
rect 10229 36125 10241 36128
rect 10275 36125 10287 36159
rect 17034 36156 17040 36168
rect 16995 36128 17040 36156
rect 10229 36119 10287 36125
rect 17034 36116 17040 36128
rect 17092 36116 17098 36168
rect 21542 36156 21548 36168
rect 21503 36128 21548 36156
rect 21542 36116 21548 36128
rect 21600 36116 21606 36168
rect 23474 36116 23480 36168
rect 23532 36156 23538 36168
rect 23860 36165 23888 36196
rect 24964 36165 24992 36196
rect 25792 36165 25820 36264
rect 28074 36252 28080 36264
rect 28132 36252 28138 36304
rect 46842 36224 46848 36236
rect 46803 36196 46848 36224
rect 46842 36184 46848 36196
rect 46900 36184 46906 36236
rect 48314 36224 48320 36236
rect 48275 36196 48320 36224
rect 48314 36184 48320 36196
rect 48372 36184 48378 36236
rect 23845 36159 23903 36165
rect 23845 36156 23857 36159
rect 23532 36128 23857 36156
rect 23532 36116 23538 36128
rect 23845 36125 23857 36128
rect 23891 36125 23903 36159
rect 23845 36119 23903 36125
rect 24029 36159 24087 36165
rect 24029 36125 24041 36159
rect 24075 36156 24087 36159
rect 24949 36159 25007 36165
rect 24075 36128 24808 36156
rect 24075 36125 24087 36128
rect 24029 36119 24087 36125
rect 7156 36060 8248 36088
rect 8389 36091 8447 36097
rect 7156 36048 7162 36060
rect 8389 36057 8401 36091
rect 8435 36088 8447 36091
rect 9582 36088 9588 36100
rect 8435 36060 9588 36088
rect 8435 36057 8447 36060
rect 8389 36051 8447 36057
rect 9582 36048 9588 36060
rect 9640 36048 9646 36100
rect 24780 36097 24808 36128
rect 24949 36125 24961 36159
rect 24995 36125 25007 36159
rect 24949 36119 25007 36125
rect 25133 36159 25191 36165
rect 25133 36125 25145 36159
rect 25179 36156 25191 36159
rect 25593 36159 25651 36165
rect 25593 36156 25605 36159
rect 25179 36128 25605 36156
rect 25179 36125 25191 36128
rect 25133 36119 25191 36125
rect 25593 36125 25605 36128
rect 25639 36125 25651 36159
rect 25593 36119 25651 36125
rect 25777 36159 25835 36165
rect 25777 36125 25789 36159
rect 25823 36125 25835 36159
rect 27430 36156 27436 36168
rect 27391 36128 27436 36156
rect 25777 36119 25835 36125
rect 24765 36091 24823 36097
rect 24765 36057 24777 36091
rect 24811 36057 24823 36091
rect 24964 36088 24992 36119
rect 27430 36116 27436 36128
rect 27488 36116 27494 36168
rect 27706 36156 27712 36168
rect 27667 36128 27712 36156
rect 27706 36116 27712 36128
rect 27764 36116 27770 36168
rect 27801 36159 27859 36165
rect 27801 36125 27813 36159
rect 27847 36156 27859 36159
rect 28442 36156 28448 36168
rect 27847 36128 28448 36156
rect 27847 36125 27859 36128
rect 27801 36119 27859 36125
rect 28442 36116 28448 36128
rect 28500 36116 28506 36168
rect 25222 36088 25228 36100
rect 24964 36060 25228 36088
rect 24765 36051 24823 36057
rect 10042 36020 10048 36032
rect 10003 35992 10048 36020
rect 10042 35980 10048 35992
rect 10100 35980 10106 36032
rect 24780 36020 24808 36051
rect 25222 36048 25228 36060
rect 25280 36048 25286 36100
rect 25685 36091 25743 36097
rect 25685 36057 25697 36091
rect 25731 36088 25743 36091
rect 26142 36088 26148 36100
rect 25731 36060 26148 36088
rect 25731 36057 25743 36060
rect 25685 36051 25743 36057
rect 26142 36048 26148 36060
rect 26200 36088 26206 36100
rect 26329 36091 26387 36097
rect 26329 36088 26341 36091
rect 26200 36060 26341 36088
rect 26200 36048 26206 36060
rect 26329 36057 26341 36060
rect 26375 36057 26387 36091
rect 26329 36051 26387 36057
rect 27617 36091 27675 36097
rect 27617 36057 27629 36091
rect 27663 36057 27675 36091
rect 48130 36088 48136 36100
rect 48091 36060 48136 36088
rect 27617 36051 27675 36057
rect 25038 36020 25044 36032
rect 24780 35992 25044 36020
rect 25038 35980 25044 35992
rect 25096 36020 25102 36032
rect 26050 36020 26056 36032
rect 25096 35992 26056 36020
rect 25096 35980 25102 35992
rect 26050 35980 26056 35992
rect 26108 35980 26114 36032
rect 26510 35980 26516 36032
rect 26568 36029 26574 36032
rect 26568 36023 26587 36029
rect 26575 35989 26587 36023
rect 27632 36020 27660 36051
rect 48130 36048 48136 36060
rect 48188 36048 48194 36100
rect 27798 36020 27804 36032
rect 27632 35992 27804 36020
rect 26568 35983 26587 35989
rect 26568 35980 26574 35983
rect 27798 35980 27804 35992
rect 27856 35980 27862 36032
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 5629 35819 5687 35825
rect 5629 35785 5641 35819
rect 5675 35816 5687 35819
rect 6178 35816 6184 35828
rect 5675 35788 6184 35816
rect 5675 35785 5687 35788
rect 5629 35779 5687 35785
rect 6178 35776 6184 35788
rect 6236 35776 6242 35828
rect 14090 35816 14096 35828
rect 14051 35788 14096 35816
rect 14090 35776 14096 35788
rect 14148 35776 14154 35828
rect 21361 35819 21419 35825
rect 21361 35785 21373 35819
rect 21407 35816 21419 35819
rect 21726 35816 21732 35828
rect 21407 35788 21732 35816
rect 21407 35785 21419 35788
rect 21361 35779 21419 35785
rect 21726 35776 21732 35788
rect 21784 35776 21790 35828
rect 24026 35776 24032 35828
rect 24084 35816 24090 35828
rect 24762 35816 24768 35828
rect 24084 35788 24768 35816
rect 24084 35776 24090 35788
rect 24762 35776 24768 35788
rect 24820 35776 24826 35828
rect 24854 35776 24860 35828
rect 24912 35816 24918 35828
rect 24949 35819 25007 35825
rect 24949 35816 24961 35819
rect 24912 35788 24961 35816
rect 24912 35776 24918 35788
rect 24949 35785 24961 35788
rect 24995 35785 25007 35819
rect 24949 35779 25007 35785
rect 25222 35776 25228 35828
rect 25280 35816 25286 35828
rect 28718 35816 28724 35828
rect 25280 35788 28724 35816
rect 25280 35776 25286 35788
rect 28718 35776 28724 35788
rect 28776 35776 28782 35828
rect 47857 35819 47915 35825
rect 47857 35785 47869 35819
rect 47903 35816 47915 35819
rect 48130 35816 48136 35828
rect 47903 35788 48136 35816
rect 47903 35785 47915 35788
rect 47857 35779 47915 35785
rect 48130 35776 48136 35788
rect 48188 35776 48194 35828
rect 9340 35751 9398 35757
rect 9340 35717 9352 35751
rect 9386 35748 9398 35751
rect 10042 35748 10048 35760
rect 9386 35720 10048 35748
rect 9386 35717 9398 35720
rect 9340 35711 9398 35717
rect 10042 35708 10048 35720
rect 10100 35708 10106 35760
rect 15930 35748 15936 35760
rect 14384 35720 15936 35748
rect 5166 35680 5172 35692
rect 5127 35652 5172 35680
rect 5166 35640 5172 35652
rect 5224 35640 5230 35692
rect 9582 35680 9588 35692
rect 9543 35652 9588 35680
rect 9582 35640 9588 35652
rect 9640 35640 9646 35692
rect 14090 35683 14148 35689
rect 14090 35649 14102 35683
rect 14136 35680 14148 35683
rect 14384 35680 14412 35720
rect 15930 35708 15936 35720
rect 15988 35708 15994 35760
rect 25774 35748 25780 35760
rect 22296 35720 25780 35748
rect 14550 35680 14556 35692
rect 14136 35652 14412 35680
rect 14511 35652 14556 35680
rect 14136 35649 14148 35652
rect 14090 35643 14148 35649
rect 14550 35640 14556 35652
rect 14608 35640 14614 35692
rect 18141 35683 18199 35689
rect 18141 35649 18153 35683
rect 18187 35680 18199 35683
rect 19242 35680 19248 35692
rect 18187 35652 19248 35680
rect 18187 35649 18199 35652
rect 18141 35643 18199 35649
rect 19242 35640 19248 35652
rect 19300 35640 19306 35692
rect 21269 35683 21327 35689
rect 21269 35649 21281 35683
rect 21315 35680 21327 35683
rect 22002 35680 22008 35692
rect 21315 35652 22008 35680
rect 21315 35649 21327 35652
rect 21269 35643 21327 35649
rect 22002 35640 22008 35652
rect 22060 35640 22066 35692
rect 22296 35689 22324 35720
rect 25774 35708 25780 35720
rect 25832 35708 25838 35760
rect 26510 35748 26516 35760
rect 26423 35720 26516 35748
rect 22281 35683 22339 35689
rect 22281 35649 22293 35683
rect 22327 35649 22339 35683
rect 22281 35643 22339 35649
rect 23293 35683 23351 35689
rect 23293 35649 23305 35683
rect 23339 35680 23351 35683
rect 23474 35680 23480 35692
rect 23339 35652 23480 35680
rect 23339 35649 23351 35652
rect 23293 35643 23351 35649
rect 23474 35640 23480 35652
rect 23532 35640 23538 35692
rect 24765 35683 24823 35689
rect 24765 35649 24777 35683
rect 24811 35680 24823 35683
rect 24946 35680 24952 35692
rect 24811 35652 24952 35680
rect 24811 35649 24823 35652
rect 24765 35643 24823 35649
rect 24946 35640 24952 35652
rect 25004 35640 25010 35692
rect 25041 35683 25099 35689
rect 25041 35649 25053 35683
rect 25087 35680 25099 35683
rect 25590 35680 25596 35692
rect 25087 35652 25596 35680
rect 25087 35649 25099 35652
rect 25041 35643 25099 35649
rect 25590 35640 25596 35652
rect 25648 35680 25654 35692
rect 25961 35683 26019 35689
rect 25961 35680 25973 35683
rect 25648 35652 25973 35680
rect 25648 35640 25654 35652
rect 25961 35649 25973 35652
rect 26007 35649 26019 35683
rect 26142 35680 26148 35692
rect 26103 35652 26148 35680
rect 25961 35643 26019 35649
rect 26142 35640 26148 35652
rect 26200 35640 26206 35692
rect 26326 35680 26332 35692
rect 26287 35652 26332 35680
rect 26326 35640 26332 35652
rect 26384 35640 26390 35692
rect 26436 35689 26464 35720
rect 26510 35708 26516 35720
rect 26568 35748 26574 35760
rect 27157 35751 27215 35757
rect 27157 35748 27169 35751
rect 26568 35720 27169 35748
rect 26568 35708 26574 35720
rect 27157 35717 27169 35720
rect 27203 35717 27215 35751
rect 27157 35711 27215 35717
rect 26421 35683 26479 35689
rect 26421 35649 26433 35683
rect 26467 35649 26479 35683
rect 26421 35643 26479 35649
rect 27338 35640 27344 35692
rect 27396 35680 27402 35692
rect 27433 35683 27491 35689
rect 27433 35680 27445 35683
rect 27396 35652 27445 35680
rect 27396 35640 27402 35652
rect 27433 35649 27445 35652
rect 27479 35649 27491 35683
rect 27433 35643 27491 35649
rect 32309 35683 32367 35689
rect 32309 35649 32321 35683
rect 32355 35680 32367 35683
rect 32398 35680 32404 35692
rect 32355 35652 32404 35680
rect 32355 35649 32367 35652
rect 32309 35643 32367 35649
rect 32398 35640 32404 35652
rect 32456 35640 32462 35692
rect 32576 35683 32634 35689
rect 32576 35649 32588 35683
rect 32622 35680 32634 35683
rect 33042 35680 33048 35692
rect 32622 35652 33048 35680
rect 32622 35649 32634 35652
rect 32576 35643 32634 35649
rect 33042 35640 33048 35652
rect 33100 35640 33106 35692
rect 34790 35640 34796 35692
rect 34848 35680 34854 35692
rect 35253 35683 35311 35689
rect 35253 35680 35265 35683
rect 34848 35652 35265 35680
rect 34848 35640 34854 35652
rect 35253 35649 35265 35652
rect 35299 35649 35311 35683
rect 35253 35643 35311 35649
rect 35437 35683 35495 35689
rect 35437 35649 35449 35683
rect 35483 35649 35495 35683
rect 35437 35643 35495 35649
rect 17954 35572 17960 35624
rect 18012 35612 18018 35624
rect 18049 35615 18107 35621
rect 18049 35612 18061 35615
rect 18012 35584 18061 35612
rect 18012 35572 18018 35584
rect 18049 35581 18061 35584
rect 18095 35581 18107 35615
rect 23198 35612 23204 35624
rect 23159 35584 23204 35612
rect 18049 35575 18107 35581
rect 23198 35572 23204 35584
rect 23256 35572 23262 35624
rect 24118 35612 24124 35624
rect 23308 35584 24124 35612
rect 17678 35504 17684 35556
rect 17736 35544 17742 35556
rect 17773 35547 17831 35553
rect 17773 35544 17785 35547
rect 17736 35516 17785 35544
rect 17736 35504 17742 35516
rect 17773 35513 17785 35516
rect 17819 35513 17831 35547
rect 23308 35544 23336 35584
rect 24118 35572 24124 35584
rect 24176 35572 24182 35624
rect 27062 35572 27068 35624
rect 27120 35612 27126 35624
rect 27157 35615 27215 35621
rect 27157 35612 27169 35615
rect 27120 35584 27169 35612
rect 27120 35572 27126 35584
rect 27157 35581 27169 35584
rect 27203 35581 27215 35615
rect 27157 35575 27215 35581
rect 34698 35572 34704 35624
rect 34756 35612 34762 35624
rect 35452 35612 35480 35643
rect 47118 35640 47124 35692
rect 47176 35680 47182 35692
rect 47765 35683 47823 35689
rect 47765 35680 47777 35683
rect 47176 35652 47777 35680
rect 47176 35640 47182 35652
rect 47765 35649 47777 35652
rect 47811 35649 47823 35683
rect 47765 35643 47823 35649
rect 34756 35584 35480 35612
rect 34756 35572 34762 35584
rect 17773 35507 17831 35513
rect 18064 35516 23336 35544
rect 23661 35547 23719 35553
rect 18064 35488 18092 35516
rect 23661 35513 23673 35547
rect 23707 35544 23719 35547
rect 24762 35544 24768 35556
rect 23707 35516 24768 35544
rect 23707 35513 23719 35516
rect 23661 35507 23719 35513
rect 24762 35504 24768 35516
rect 24820 35504 24826 35556
rect 24946 35504 24952 35556
rect 25004 35544 25010 35556
rect 26050 35544 26056 35556
rect 25004 35516 26056 35544
rect 25004 35504 25010 35516
rect 26050 35504 26056 35516
rect 26108 35504 26114 35556
rect 5442 35476 5448 35488
rect 5403 35448 5448 35476
rect 5442 35436 5448 35448
rect 5500 35436 5506 35488
rect 8110 35436 8116 35488
rect 8168 35476 8174 35488
rect 8205 35479 8263 35485
rect 8205 35476 8217 35479
rect 8168 35448 8217 35476
rect 8168 35436 8174 35448
rect 8205 35445 8217 35448
rect 8251 35445 8263 35479
rect 8205 35439 8263 35445
rect 13909 35479 13967 35485
rect 13909 35445 13921 35479
rect 13955 35476 13967 35479
rect 13998 35476 14004 35488
rect 13955 35448 14004 35476
rect 13955 35445 13967 35448
rect 13909 35439 13967 35445
rect 13998 35436 14004 35448
rect 14056 35436 14062 35488
rect 14458 35476 14464 35488
rect 14419 35448 14464 35476
rect 14458 35436 14464 35448
rect 14516 35436 14522 35488
rect 18046 35436 18052 35488
rect 18104 35436 18110 35488
rect 21450 35436 21456 35488
rect 21508 35476 21514 35488
rect 22189 35479 22247 35485
rect 22189 35476 22201 35479
rect 21508 35448 22201 35476
rect 21508 35436 21514 35448
rect 22189 35445 22201 35448
rect 22235 35445 22247 35479
rect 22189 35439 22247 35445
rect 23750 35436 23756 35488
rect 23808 35476 23814 35488
rect 24581 35479 24639 35485
rect 24581 35476 24593 35479
rect 23808 35448 24593 35476
rect 23808 35436 23814 35448
rect 24581 35445 24593 35448
rect 24627 35445 24639 35479
rect 24581 35439 24639 35445
rect 25130 35436 25136 35488
rect 25188 35476 25194 35488
rect 27341 35479 27399 35485
rect 27341 35476 27353 35479
rect 25188 35448 27353 35476
rect 25188 35436 25194 35448
rect 27341 35445 27353 35448
rect 27387 35476 27399 35479
rect 27706 35476 27712 35488
rect 27387 35448 27712 35476
rect 27387 35445 27399 35448
rect 27341 35439 27399 35445
rect 27706 35436 27712 35448
rect 27764 35476 27770 35488
rect 28626 35476 28632 35488
rect 27764 35448 28632 35476
rect 27764 35436 27770 35448
rect 28626 35436 28632 35448
rect 28684 35436 28690 35488
rect 33502 35436 33508 35488
rect 33560 35476 33566 35488
rect 33689 35479 33747 35485
rect 33689 35476 33701 35479
rect 33560 35448 33701 35476
rect 33560 35436 33566 35448
rect 33689 35445 33701 35448
rect 33735 35445 33747 35479
rect 33689 35439 33747 35445
rect 35345 35479 35403 35485
rect 35345 35445 35357 35479
rect 35391 35476 35403 35479
rect 35434 35476 35440 35488
rect 35391 35448 35440 35476
rect 35391 35445 35403 35448
rect 35345 35439 35403 35445
rect 35434 35436 35440 35448
rect 35492 35436 35498 35488
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 5442 35232 5448 35284
rect 5500 35272 5506 35284
rect 5721 35275 5779 35281
rect 5721 35272 5733 35275
rect 5500 35244 5733 35272
rect 5500 35232 5506 35244
rect 5721 35241 5733 35244
rect 5767 35241 5779 35275
rect 5721 35235 5779 35241
rect 20993 35275 21051 35281
rect 20993 35241 21005 35275
rect 21039 35272 21051 35275
rect 21542 35272 21548 35284
rect 21039 35244 21548 35272
rect 21039 35241 21051 35244
rect 20993 35235 21051 35241
rect 21542 35232 21548 35244
rect 21600 35232 21606 35284
rect 22557 35275 22615 35281
rect 22557 35241 22569 35275
rect 22603 35272 22615 35275
rect 23198 35272 23204 35284
rect 22603 35244 23204 35272
rect 22603 35241 22615 35244
rect 22557 35235 22615 35241
rect 23198 35232 23204 35244
rect 23256 35272 23262 35284
rect 25038 35272 25044 35284
rect 23256 35244 23980 35272
rect 24999 35244 25044 35272
rect 23256 35232 23262 35244
rect 8294 35164 8300 35216
rect 8352 35164 8358 35216
rect 17037 35207 17095 35213
rect 17037 35173 17049 35207
rect 17083 35204 17095 35207
rect 17954 35204 17960 35216
rect 17083 35176 17960 35204
rect 17083 35173 17095 35176
rect 17037 35167 17095 35173
rect 17954 35164 17960 35176
rect 18012 35164 18018 35216
rect 23952 35204 23980 35244
rect 25038 35232 25044 35244
rect 25096 35232 25102 35284
rect 25130 35232 25136 35284
rect 25188 35272 25194 35284
rect 25774 35272 25780 35284
rect 25188 35244 25233 35272
rect 25735 35244 25780 35272
rect 25188 35232 25194 35244
rect 25774 35232 25780 35244
rect 25832 35232 25838 35284
rect 26237 35275 26295 35281
rect 26237 35241 26249 35275
rect 26283 35241 26295 35275
rect 26237 35235 26295 35241
rect 27341 35275 27399 35281
rect 27341 35241 27353 35275
rect 27387 35272 27399 35275
rect 27430 35272 27436 35284
rect 27387 35244 27436 35272
rect 27387 35241 27399 35244
rect 27341 35235 27399 35241
rect 24949 35207 25007 35213
rect 24949 35204 24961 35207
rect 23952 35176 24961 35204
rect 24949 35173 24961 35176
rect 24995 35173 25007 35207
rect 26252 35204 26280 35235
rect 27430 35232 27436 35244
rect 27488 35232 27494 35284
rect 33042 35272 33048 35284
rect 33003 35244 33048 35272
rect 33042 35232 33048 35244
rect 33100 35232 33106 35284
rect 35866 35244 38976 35272
rect 28353 35207 28411 35213
rect 28353 35204 28365 35207
rect 26252 35176 28365 35204
rect 24949 35167 25007 35173
rect 8312 35136 8340 35164
rect 8389 35139 8447 35145
rect 8389 35136 8401 35139
rect 8312 35108 8401 35136
rect 8389 35105 8401 35108
rect 8435 35105 8447 35139
rect 15654 35136 15660 35148
rect 15615 35108 15660 35136
rect 8389 35099 8447 35105
rect 15654 35096 15660 35108
rect 15712 35096 15718 35148
rect 17494 35096 17500 35148
rect 17552 35136 17558 35148
rect 17773 35139 17831 35145
rect 17773 35136 17785 35139
rect 17552 35108 17785 35136
rect 17552 35096 17558 35108
rect 17773 35105 17785 35108
rect 17819 35105 17831 35139
rect 20806 35136 20812 35148
rect 20767 35108 20812 35136
rect 17773 35099 17831 35105
rect 20806 35096 20812 35108
rect 20864 35096 20870 35148
rect 21450 35136 21456 35148
rect 20916 35108 21456 35136
rect 4338 35068 4344 35080
rect 4299 35040 4344 35068
rect 4338 35028 4344 35040
rect 4396 35028 4402 35080
rect 8110 35028 8116 35080
rect 8168 35068 8174 35080
rect 8297 35071 8355 35077
rect 8297 35068 8309 35071
rect 8168 35040 8309 35068
rect 8168 35028 8174 35040
rect 8297 35037 8309 35040
rect 8343 35037 8355 35071
rect 8297 35031 8355 35037
rect 16666 35028 16672 35080
rect 16724 35068 16730 35080
rect 17678 35068 17684 35080
rect 16724 35040 17684 35068
rect 16724 35028 16730 35040
rect 17678 35028 17684 35040
rect 17736 35028 17742 35080
rect 17865 35071 17923 35077
rect 17865 35037 17877 35071
rect 17911 35037 17923 35071
rect 17865 35031 17923 35037
rect 17957 35071 18015 35077
rect 17957 35037 17969 35071
rect 18003 35068 18015 35071
rect 18046 35068 18052 35080
rect 18003 35040 18052 35068
rect 18003 35037 18015 35040
rect 17957 35031 18015 35037
rect 4608 35003 4666 35009
rect 4608 34969 4620 35003
rect 4654 35000 4666 35003
rect 5718 35000 5724 35012
rect 4654 34972 5724 35000
rect 4654 34969 4666 34972
rect 4608 34963 4666 34969
rect 5718 34960 5724 34972
rect 5776 34960 5782 35012
rect 15924 35003 15982 35009
rect 15924 34969 15936 35003
rect 15970 35000 15982 35003
rect 16850 35000 16856 35012
rect 15970 34972 16856 35000
rect 15970 34969 15982 34972
rect 15924 34963 15982 34969
rect 16850 34960 16856 34972
rect 16908 34960 16914 35012
rect 17218 35000 17224 35012
rect 16960 34972 17224 35000
rect 7098 34892 7104 34944
rect 7156 34932 7162 34944
rect 7929 34935 7987 34941
rect 7929 34932 7941 34935
rect 7156 34904 7941 34932
rect 7156 34892 7162 34904
rect 7929 34901 7941 34904
rect 7975 34901 7987 34935
rect 7929 34895 7987 34901
rect 16574 34892 16580 34944
rect 16632 34932 16638 34944
rect 16960 34932 16988 34972
rect 17218 34960 17224 34972
rect 17276 35000 17282 35012
rect 17880 35000 17908 35031
rect 18046 35028 18052 35040
rect 18104 35028 18110 35080
rect 20625 35071 20683 35077
rect 20625 35037 20637 35071
rect 20671 35068 20683 35071
rect 20916 35068 20944 35108
rect 21450 35096 21456 35108
rect 21508 35096 21514 35148
rect 26142 35136 26148 35148
rect 26103 35108 26148 35136
rect 26142 35096 26148 35108
rect 26200 35096 26206 35148
rect 27614 35136 27620 35148
rect 27575 35108 27620 35136
rect 27614 35096 27620 35108
rect 27672 35096 27678 35148
rect 20671 35040 20944 35068
rect 20993 35071 21051 35077
rect 20671 35037 20683 35040
rect 20625 35031 20683 35037
rect 20993 35037 21005 35071
rect 21039 35068 21051 35071
rect 21039 35040 23796 35068
rect 21039 35037 21051 35040
rect 20993 35031 21051 35037
rect 17276 34972 17908 35000
rect 17276 34960 17282 34972
rect 20898 34960 20904 35012
rect 20956 35000 20962 35012
rect 21821 35003 21879 35009
rect 20956 34972 21680 35000
rect 20956 34960 20962 34972
rect 16632 34904 16988 34932
rect 16632 34892 16638 34904
rect 17126 34892 17132 34944
rect 17184 34932 17190 34944
rect 17497 34935 17555 34941
rect 17497 34932 17509 34935
rect 17184 34904 17509 34932
rect 17184 34892 17190 34904
rect 17497 34901 17509 34904
rect 17543 34901 17555 34935
rect 20714 34932 20720 34944
rect 20675 34904 20720 34932
rect 17497 34895 17555 34901
rect 20714 34892 20720 34904
rect 20772 34892 20778 34944
rect 21542 34932 21548 34944
rect 21503 34904 21548 34932
rect 21542 34892 21548 34904
rect 21600 34892 21606 34944
rect 21652 34932 21680 34972
rect 21821 34969 21833 35003
rect 21867 35000 21879 35003
rect 23474 35000 23480 35012
rect 21867 34972 23480 35000
rect 21867 34969 21879 34972
rect 21821 34963 21879 34969
rect 23474 34960 23480 34972
rect 23532 34960 23538 35012
rect 23658 35000 23664 35012
rect 23716 35009 23722 35012
rect 23628 34972 23664 35000
rect 23658 34960 23664 34972
rect 23716 34963 23728 35009
rect 23768 35000 23796 35040
rect 23842 35028 23848 35080
rect 23900 35068 23906 35080
rect 23937 35071 23995 35077
rect 23937 35068 23949 35071
rect 23900 35040 23949 35068
rect 23900 35028 23906 35040
rect 23937 35037 23949 35040
rect 23983 35037 23995 35071
rect 24857 35071 24915 35077
rect 24857 35068 24869 35071
rect 23937 35031 23995 35037
rect 24688 35040 24869 35068
rect 24581 35003 24639 35009
rect 24581 35000 24593 35003
rect 23768 34972 24593 35000
rect 24581 34969 24593 34972
rect 24627 34969 24639 35003
rect 24581 34963 24639 34969
rect 23716 34960 23722 34963
rect 24688 34932 24716 35040
rect 24857 35037 24869 35040
rect 24903 35037 24915 35071
rect 24857 35031 24915 35037
rect 25317 35071 25375 35077
rect 25317 35037 25329 35071
rect 25363 35068 25375 35071
rect 25866 35068 25872 35080
rect 25363 35040 25872 35068
rect 25363 35037 25375 35040
rect 25317 35031 25375 35037
rect 25866 35028 25872 35040
rect 25924 35028 25930 35080
rect 25961 35071 26019 35077
rect 25961 35037 25973 35071
rect 26007 35037 26019 35071
rect 25961 35031 26019 35037
rect 24854 34932 24860 34944
rect 21652 34904 24860 34932
rect 24854 34892 24860 34904
rect 24912 34892 24918 34944
rect 25976 34932 26004 35031
rect 26234 35028 26240 35080
rect 26292 35068 26298 35080
rect 26292 35040 26337 35068
rect 26292 35028 26298 35040
rect 27522 35028 27528 35080
rect 27580 35068 27586 35080
rect 27724 35077 27752 35176
rect 28353 35173 28365 35176
rect 28399 35173 28411 35207
rect 28353 35167 28411 35173
rect 32306 35164 32312 35216
rect 32364 35204 32370 35216
rect 35866 35204 35894 35244
rect 32364 35176 35894 35204
rect 32364 35164 32370 35176
rect 28626 35136 28632 35148
rect 28587 35108 28632 35136
rect 28626 35096 28632 35108
rect 28684 35096 28690 35148
rect 33502 35136 33508 35148
rect 31864 35108 32444 35136
rect 33463 35108 33508 35136
rect 27709 35071 27767 35077
rect 27709 35068 27721 35071
rect 27580 35040 27721 35068
rect 27580 35028 27586 35040
rect 27709 35037 27721 35040
rect 27755 35037 27767 35071
rect 28718 35068 28724 35080
rect 28679 35040 28724 35068
rect 27709 35031 27767 35037
rect 28718 35028 28724 35040
rect 28776 35028 28782 35080
rect 29730 35028 29736 35080
rect 29788 35068 29794 35080
rect 29825 35071 29883 35077
rect 29825 35068 29837 35071
rect 29788 35040 29837 35068
rect 29788 35028 29794 35040
rect 29825 35037 29837 35040
rect 29871 35037 29883 35071
rect 29825 35031 29883 35037
rect 30466 35028 30472 35080
rect 30524 35068 30530 35080
rect 31864 35068 31892 35108
rect 30524 35040 31892 35068
rect 31941 35071 31999 35077
rect 30524 35028 30530 35040
rect 31941 35037 31953 35071
rect 31987 35037 31999 35071
rect 31941 35031 31999 35037
rect 32125 35071 32183 35077
rect 32125 35037 32137 35071
rect 32171 35068 32183 35071
rect 32306 35068 32312 35080
rect 32171 35040 32312 35068
rect 32171 35037 32183 35040
rect 32125 35031 32183 35037
rect 29362 34960 29368 35012
rect 29420 35000 29426 35012
rect 30070 35003 30128 35009
rect 30070 35000 30082 35003
rect 29420 34972 30082 35000
rect 29420 34960 29426 34972
rect 30070 34969 30082 34972
rect 30116 34969 30128 35003
rect 30070 34963 30128 34969
rect 30190 34960 30196 35012
rect 30248 35000 30254 35012
rect 31956 35000 31984 35031
rect 32306 35028 32312 35040
rect 32364 35028 32370 35080
rect 32416 35077 32444 35108
rect 33502 35096 33508 35108
rect 33560 35096 33566 35148
rect 35342 35096 35348 35148
rect 35400 35136 35406 35148
rect 36909 35139 36967 35145
rect 36909 35136 36921 35139
rect 35400 35108 36921 35136
rect 35400 35096 35406 35108
rect 36909 35105 36921 35108
rect 36955 35105 36967 35139
rect 36909 35099 36967 35105
rect 32401 35071 32459 35077
rect 32401 35037 32413 35071
rect 32447 35037 32459 35071
rect 32401 35031 32459 35037
rect 32585 35071 32643 35077
rect 32585 35037 32597 35071
rect 32631 35068 32643 35071
rect 33229 35071 33287 35077
rect 33229 35068 33241 35071
rect 32631 35040 33241 35068
rect 32631 35037 32643 35040
rect 32585 35031 32643 35037
rect 33229 35037 33241 35040
rect 33275 35037 33287 35071
rect 33413 35071 33471 35077
rect 33413 35068 33425 35071
rect 33229 35031 33287 35037
rect 33336 35040 33425 35068
rect 32674 35000 32680 35012
rect 30248 34972 31892 35000
rect 31956 34972 32680 35000
rect 30248 34960 30254 34972
rect 27154 34932 27160 34944
rect 25976 34904 27160 34932
rect 27154 34892 27160 34904
rect 27212 34892 27218 34944
rect 31202 34932 31208 34944
rect 31163 34904 31208 34932
rect 31202 34892 31208 34904
rect 31260 34892 31266 34944
rect 31864 34932 31892 34972
rect 32674 34960 32680 34972
rect 32732 34960 32738 35012
rect 33336 34932 33364 35040
rect 33413 35037 33425 35040
rect 33459 35037 33471 35071
rect 33413 35031 33471 35037
rect 35713 35071 35771 35077
rect 35713 35037 35725 35071
rect 35759 35068 35771 35071
rect 35802 35068 35808 35080
rect 35759 35040 35808 35068
rect 35759 35037 35771 35040
rect 35713 35031 35771 35037
rect 35802 35028 35808 35040
rect 35860 35028 35866 35080
rect 35986 35028 35992 35080
rect 36044 35068 36050 35080
rect 36173 35071 36231 35077
rect 36173 35068 36185 35071
rect 36044 35040 36185 35068
rect 36044 35028 36050 35040
rect 36173 35037 36185 35040
rect 36219 35037 36231 35071
rect 36173 35031 36231 35037
rect 36357 35071 36415 35077
rect 36357 35037 36369 35071
rect 36403 35068 36415 35071
rect 36998 35068 37004 35080
rect 36403 35040 37004 35068
rect 36403 35037 36415 35040
rect 36357 35031 36415 35037
rect 36998 35028 37004 35040
rect 37056 35028 37062 35080
rect 38654 35028 38660 35080
rect 38712 35068 38718 35080
rect 38948 35077 38976 35244
rect 38749 35071 38807 35077
rect 38749 35068 38761 35071
rect 38712 35040 38761 35068
rect 38712 35028 38718 35040
rect 38749 35037 38761 35040
rect 38795 35037 38807 35071
rect 38749 35031 38807 35037
rect 38933 35071 38991 35077
rect 38933 35037 38945 35071
rect 38979 35068 38991 35071
rect 39022 35068 39028 35080
rect 38979 35040 39028 35068
rect 38979 35037 38991 35040
rect 38933 35031 38991 35037
rect 39022 35028 39028 35040
rect 39080 35028 39086 35080
rect 39206 35068 39212 35080
rect 39167 35040 39212 35068
rect 39206 35028 39212 35040
rect 39264 35028 39270 35080
rect 34698 34960 34704 35012
rect 34756 35000 34762 35012
rect 35437 35003 35495 35009
rect 35437 35000 35449 35003
rect 34756 34972 35449 35000
rect 34756 34960 34762 34972
rect 35437 34969 35449 34972
rect 35483 34969 35495 35003
rect 35618 35000 35624 35012
rect 35579 34972 35624 35000
rect 35437 34963 35495 34969
rect 35618 34960 35624 34972
rect 35676 35000 35682 35012
rect 36814 35000 36820 35012
rect 35676 34972 36820 35000
rect 35676 34960 35682 34972
rect 36814 34960 36820 34972
rect 36872 34960 36878 35012
rect 36906 34960 36912 35012
rect 36964 35000 36970 35012
rect 37154 35003 37212 35009
rect 37154 35000 37166 35003
rect 36964 34972 37166 35000
rect 36964 34960 36970 34972
rect 37154 34969 37166 34972
rect 37200 34969 37212 35003
rect 37154 34963 37212 34969
rect 34422 34932 34428 34944
rect 31864 34904 34428 34932
rect 34422 34892 34428 34904
rect 34480 34892 34486 34944
rect 35526 34932 35532 34944
rect 35487 34904 35532 34932
rect 35526 34892 35532 34904
rect 35584 34892 35590 34944
rect 36262 34932 36268 34944
rect 36223 34904 36268 34932
rect 36262 34892 36268 34904
rect 36320 34892 36326 34944
rect 37642 34892 37648 34944
rect 37700 34932 37706 34944
rect 38289 34935 38347 34941
rect 38289 34932 38301 34935
rect 37700 34904 38301 34932
rect 37700 34892 37706 34904
rect 38289 34901 38301 34904
rect 38335 34901 38347 34935
rect 38289 34895 38347 34901
rect 38930 34892 38936 34944
rect 38988 34932 38994 34944
rect 39393 34935 39451 34941
rect 39393 34932 39405 34935
rect 38988 34904 39405 34932
rect 38988 34892 38994 34904
rect 39393 34901 39405 34904
rect 39439 34901 39451 34935
rect 39393 34895 39451 34901
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 1765 34731 1823 34737
rect 1765 34697 1777 34731
rect 1811 34728 1823 34731
rect 1946 34728 1952 34740
rect 1811 34700 1952 34728
rect 1811 34697 1823 34700
rect 1765 34691 1823 34697
rect 1946 34688 1952 34700
rect 2004 34688 2010 34740
rect 4338 34688 4344 34740
rect 4396 34728 4402 34740
rect 4433 34731 4491 34737
rect 4433 34728 4445 34731
rect 4396 34700 4445 34728
rect 4396 34688 4402 34700
rect 4433 34697 4445 34700
rect 4479 34697 4491 34731
rect 5718 34728 5724 34740
rect 5679 34700 5724 34728
rect 4433 34691 4491 34697
rect 5718 34688 5724 34700
rect 5776 34688 5782 34740
rect 7742 34728 7748 34740
rect 6886 34700 7748 34728
rect 6886 34660 6914 34700
rect 7742 34688 7748 34700
rect 7800 34688 7806 34740
rect 8018 34688 8024 34740
rect 8076 34728 8082 34740
rect 9033 34731 9091 34737
rect 8076 34700 8984 34728
rect 8076 34688 8082 34700
rect 5276 34632 6914 34660
rect 7116 34632 8340 34660
rect 1578 34592 1584 34604
rect 1539 34564 1584 34592
rect 1578 34552 1584 34564
rect 1636 34552 1642 34604
rect 4617 34595 4675 34601
rect 4617 34561 4629 34595
rect 4663 34592 4675 34595
rect 4798 34592 4804 34604
rect 4663 34564 4804 34592
rect 4663 34561 4675 34564
rect 4617 34555 4675 34561
rect 4798 34552 4804 34564
rect 4856 34592 4862 34604
rect 4982 34592 4988 34604
rect 4856 34564 4988 34592
rect 4856 34552 4862 34564
rect 4982 34552 4988 34564
rect 5040 34552 5046 34604
rect 5276 34601 5304 34632
rect 5077 34595 5135 34601
rect 5077 34561 5089 34595
rect 5123 34561 5135 34595
rect 5077 34555 5135 34561
rect 5261 34595 5319 34601
rect 5261 34561 5273 34595
rect 5307 34561 5319 34595
rect 5902 34592 5908 34604
rect 5863 34564 5908 34592
rect 5261 34555 5319 34561
rect 5092 34524 5120 34555
rect 5902 34552 5908 34564
rect 5960 34552 5966 34604
rect 5166 34524 5172 34536
rect 5079 34496 5172 34524
rect 4982 34416 4988 34468
rect 5040 34456 5046 34468
rect 5092 34456 5120 34496
rect 5166 34484 5172 34496
rect 5224 34524 5230 34536
rect 7116 34533 7144 34632
rect 7377 34595 7435 34601
rect 7377 34561 7389 34595
rect 7423 34592 7435 34595
rect 7742 34592 7748 34604
rect 7423 34564 7748 34592
rect 7423 34561 7435 34564
rect 7377 34555 7435 34561
rect 7742 34552 7748 34564
rect 7800 34552 7806 34604
rect 7101 34527 7159 34533
rect 7101 34524 7113 34527
rect 5224 34496 7113 34524
rect 5224 34484 5230 34496
rect 7101 34493 7113 34496
rect 7147 34493 7159 34527
rect 7101 34487 7159 34493
rect 7282 34484 7288 34536
rect 7340 34524 7346 34536
rect 8110 34524 8116 34536
rect 7340 34496 8116 34524
rect 7340 34484 7346 34496
rect 8110 34484 8116 34496
rect 8168 34484 8174 34536
rect 5040 34428 5120 34456
rect 8312 34456 8340 34632
rect 8849 34595 8907 34601
rect 8849 34561 8861 34595
rect 8895 34561 8907 34595
rect 8956 34592 8984 34700
rect 9033 34697 9045 34731
rect 9079 34728 9091 34731
rect 9674 34728 9680 34740
rect 9079 34700 9680 34728
rect 9079 34697 9091 34700
rect 9033 34691 9091 34697
rect 9674 34688 9680 34700
rect 9732 34688 9738 34740
rect 14458 34728 14464 34740
rect 10980 34700 14464 34728
rect 9677 34595 9735 34601
rect 9677 34592 9689 34595
rect 8956 34564 9689 34592
rect 8849 34555 8907 34561
rect 9677 34561 9689 34564
rect 9723 34592 9735 34595
rect 10980 34592 11008 34700
rect 14458 34688 14464 34700
rect 14516 34728 14522 34740
rect 16117 34731 16175 34737
rect 14516 34700 15056 34728
rect 14516 34688 14522 34700
rect 13722 34620 13728 34672
rect 13780 34660 13786 34672
rect 13780 34632 14872 34660
rect 13780 34620 13786 34632
rect 9723 34564 11008 34592
rect 9723 34561 9735 34564
rect 9677 34555 9735 34561
rect 8864 34524 8892 34555
rect 13998 34552 14004 34604
rect 14056 34601 14062 34604
rect 14292 34601 14320 34632
rect 14056 34592 14068 34601
rect 14277 34595 14335 34601
rect 14056 34564 14101 34592
rect 14056 34555 14068 34564
rect 14277 34561 14289 34595
rect 14323 34561 14335 34595
rect 14277 34555 14335 34561
rect 14737 34595 14795 34601
rect 14737 34561 14749 34595
rect 14783 34561 14795 34595
rect 14737 34555 14795 34561
rect 14056 34552 14062 34555
rect 9766 34524 9772 34536
rect 8864 34496 9772 34524
rect 9766 34484 9772 34496
rect 9824 34484 9830 34536
rect 14752 34524 14780 34555
rect 14292 34496 14780 34524
rect 14844 34524 14872 34632
rect 15028 34601 15056 34700
rect 16117 34697 16129 34731
rect 16163 34728 16175 34731
rect 16574 34728 16580 34740
rect 16163 34700 16580 34728
rect 16163 34697 16175 34700
rect 16117 34691 16175 34697
rect 16574 34688 16580 34700
rect 16632 34688 16638 34740
rect 16850 34728 16856 34740
rect 16811 34700 16856 34728
rect 16850 34688 16856 34700
rect 16908 34688 16914 34740
rect 20898 34728 20904 34740
rect 20859 34700 20904 34728
rect 20898 34688 20904 34700
rect 20956 34688 20962 34740
rect 22373 34731 22431 34737
rect 22373 34697 22385 34731
rect 22419 34728 22431 34731
rect 23474 34728 23480 34740
rect 22419 34700 23480 34728
rect 22419 34697 22431 34700
rect 22373 34691 22431 34697
rect 23474 34688 23480 34700
rect 23532 34688 23538 34740
rect 23658 34728 23664 34740
rect 23619 34700 23664 34728
rect 23658 34688 23664 34700
rect 23716 34688 23722 34740
rect 24857 34731 24915 34737
rect 24857 34697 24869 34731
rect 24903 34728 24915 34731
rect 24946 34728 24952 34740
rect 24903 34700 24952 34728
rect 24903 34697 24915 34700
rect 24857 34691 24915 34697
rect 24946 34688 24952 34700
rect 25004 34688 25010 34740
rect 26326 34688 26332 34740
rect 26384 34728 26390 34740
rect 27157 34731 27215 34737
rect 27157 34728 27169 34731
rect 26384 34700 27169 34728
rect 26384 34688 26390 34700
rect 27157 34697 27169 34700
rect 27203 34697 27215 34731
rect 29362 34728 29368 34740
rect 29323 34700 29368 34728
rect 27157 34691 27215 34697
rect 29362 34688 29368 34700
rect 29420 34688 29426 34740
rect 33873 34731 33931 34737
rect 33873 34697 33885 34731
rect 33919 34728 33931 34731
rect 35986 34728 35992 34740
rect 33919 34700 34652 34728
rect 35947 34700 35992 34728
rect 33919 34697 33931 34700
rect 33873 34691 33931 34697
rect 17494 34660 17500 34672
rect 16040 34632 17500 34660
rect 16040 34601 16068 34632
rect 17494 34620 17500 34632
rect 17552 34620 17558 34672
rect 21542 34660 21548 34672
rect 20732 34632 21548 34660
rect 15013 34595 15071 34601
rect 15013 34561 15025 34595
rect 15059 34561 15071 34595
rect 15013 34555 15071 34561
rect 16025 34595 16083 34601
rect 16025 34561 16037 34595
rect 16071 34561 16083 34595
rect 16025 34555 16083 34561
rect 16301 34595 16359 34601
rect 16301 34561 16313 34595
rect 16347 34592 16359 34595
rect 16666 34592 16672 34604
rect 16347 34564 16672 34592
rect 16347 34561 16359 34564
rect 16301 34555 16359 34561
rect 16666 34552 16672 34564
rect 16724 34552 16730 34604
rect 17126 34592 17132 34604
rect 17087 34564 17132 34592
rect 17126 34552 17132 34564
rect 17184 34552 17190 34604
rect 17405 34595 17463 34601
rect 17405 34561 17417 34595
rect 17451 34592 17463 34595
rect 18138 34592 18144 34604
rect 17451 34564 18144 34592
rect 17451 34561 17463 34564
rect 17405 34555 17463 34561
rect 18138 34552 18144 34564
rect 18196 34552 18202 34604
rect 18414 34592 18420 34604
rect 18375 34564 18420 34592
rect 18414 34552 18420 34564
rect 18472 34552 18478 34604
rect 18509 34595 18567 34601
rect 18509 34561 18521 34595
rect 18555 34592 18567 34595
rect 18598 34592 18604 34604
rect 18555 34564 18604 34592
rect 18555 34561 18567 34564
rect 18509 34555 18567 34561
rect 18598 34552 18604 34564
rect 18656 34552 18662 34604
rect 18693 34595 18751 34601
rect 18693 34561 18705 34595
rect 18739 34592 18751 34595
rect 18782 34592 18788 34604
rect 18739 34564 18788 34592
rect 18739 34561 18751 34564
rect 18693 34555 18751 34561
rect 18782 34552 18788 34564
rect 18840 34552 18846 34604
rect 19242 34552 19248 34604
rect 19300 34592 19306 34604
rect 20732 34601 20760 34632
rect 21542 34620 21548 34632
rect 21600 34620 21606 34672
rect 23934 34660 23940 34672
rect 23895 34632 23940 34660
rect 23934 34620 23940 34632
rect 23992 34620 23998 34672
rect 24026 34620 24032 34672
rect 24084 34660 24090 34672
rect 24167 34663 24225 34669
rect 24084 34632 24129 34660
rect 24084 34620 24090 34632
rect 24167 34629 24179 34663
rect 24213 34660 24225 34663
rect 25774 34660 25780 34672
rect 24213 34632 25780 34660
rect 24213 34629 24225 34632
rect 24167 34623 24225 34629
rect 25774 34620 25780 34632
rect 25832 34620 25838 34672
rect 32306 34660 32312 34672
rect 30760 34632 32312 34660
rect 30760 34604 30788 34632
rect 32306 34620 32312 34632
rect 32364 34620 32370 34672
rect 33502 34620 33508 34672
rect 33560 34660 33566 34672
rect 34517 34663 34575 34669
rect 34517 34660 34529 34663
rect 33560 34632 34529 34660
rect 33560 34620 33566 34632
rect 20717 34595 20775 34601
rect 20717 34592 20729 34595
rect 19300 34564 20729 34592
rect 19300 34552 19306 34564
rect 20717 34561 20729 34564
rect 20763 34561 20775 34595
rect 20717 34555 20775 34561
rect 20806 34552 20812 34604
rect 20864 34592 20870 34604
rect 21818 34592 21824 34604
rect 20864 34564 21824 34592
rect 20864 34552 20870 34564
rect 21818 34552 21824 34564
rect 21876 34592 21882 34604
rect 22373 34595 22431 34601
rect 22373 34592 22385 34595
rect 21876 34564 22385 34592
rect 21876 34552 21882 34564
rect 22373 34561 22385 34564
rect 22419 34561 22431 34595
rect 22373 34555 22431 34561
rect 23750 34552 23756 34604
rect 23808 34592 23814 34604
rect 23845 34595 23903 34601
rect 23845 34592 23857 34595
rect 23808 34564 23857 34592
rect 23808 34552 23814 34564
rect 23845 34561 23857 34564
rect 23891 34561 23903 34595
rect 24762 34592 24768 34604
rect 24723 34564 24768 34592
rect 23845 34555 23903 34561
rect 24762 34552 24768 34564
rect 24820 34552 24826 34604
rect 24854 34552 24860 34604
rect 24912 34592 24918 34604
rect 27062 34592 27068 34604
rect 24912 34564 27068 34592
rect 24912 34552 24918 34564
rect 26206 34536 26234 34564
rect 27062 34552 27068 34564
rect 27120 34552 27126 34604
rect 27154 34552 27160 34604
rect 27212 34592 27218 34604
rect 27341 34595 27399 34601
rect 27341 34592 27353 34595
rect 27212 34564 27353 34592
rect 27212 34552 27218 34564
rect 27341 34561 27353 34564
rect 27387 34561 27399 34595
rect 27522 34592 27528 34604
rect 27483 34564 27528 34592
rect 27341 34555 27399 34561
rect 27522 34552 27528 34564
rect 27580 34552 27586 34604
rect 29549 34595 29607 34601
rect 29549 34561 29561 34595
rect 29595 34592 29607 34595
rect 30285 34595 30343 34601
rect 30285 34592 30297 34595
rect 29595 34564 30297 34592
rect 29595 34561 29607 34564
rect 29549 34555 29607 34561
rect 30285 34561 30297 34564
rect 30331 34561 30343 34595
rect 30466 34592 30472 34604
rect 30427 34564 30472 34592
rect 30285 34555 30343 34561
rect 30466 34552 30472 34564
rect 30524 34552 30530 34604
rect 30742 34592 30748 34604
rect 30655 34564 30748 34592
rect 30742 34552 30748 34564
rect 30800 34552 30806 34604
rect 30926 34592 30932 34604
rect 30887 34564 30932 34592
rect 30926 34552 30932 34564
rect 30984 34592 30990 34604
rect 32490 34592 32496 34604
rect 30984 34564 32496 34592
rect 30984 34552 30990 34564
rect 32490 34552 32496 34564
rect 32548 34552 32554 34604
rect 33410 34552 33416 34604
rect 33468 34592 33474 34604
rect 33689 34595 33747 34601
rect 33689 34592 33701 34595
rect 33468 34564 33701 34592
rect 33468 34552 33474 34564
rect 33689 34561 33701 34564
rect 33735 34592 33747 34595
rect 33778 34592 33784 34604
rect 33735 34564 33784 34592
rect 33735 34561 33747 34564
rect 33689 34555 33747 34561
rect 33778 34552 33784 34564
rect 33836 34552 33842 34604
rect 33888 34601 33916 34632
rect 34517 34629 34529 34632
rect 34563 34629 34575 34663
rect 34624 34660 34652 34700
rect 35986 34688 35992 34700
rect 36044 34688 36050 34740
rect 36906 34728 36912 34740
rect 36867 34700 36912 34728
rect 36906 34688 36912 34700
rect 36964 34688 36970 34740
rect 36998 34688 37004 34740
rect 37056 34728 37062 34740
rect 37553 34731 37611 34737
rect 37553 34728 37565 34731
rect 37056 34700 37565 34728
rect 37056 34688 37062 34700
rect 37553 34697 37565 34700
rect 37599 34697 37611 34731
rect 37553 34691 37611 34697
rect 34790 34660 34796 34672
rect 34624 34632 34796 34660
rect 34517 34623 34575 34629
rect 34790 34620 34796 34632
rect 34848 34620 34854 34672
rect 35802 34660 35808 34672
rect 35763 34632 35808 34660
rect 35802 34620 35808 34632
rect 35860 34660 35866 34672
rect 38556 34663 38614 34669
rect 35860 34632 37688 34660
rect 35860 34620 35866 34632
rect 33873 34595 33931 34601
rect 33873 34561 33885 34595
rect 33919 34561 33931 34595
rect 33873 34555 33931 34561
rect 33962 34552 33968 34604
rect 34020 34592 34026 34604
rect 34333 34595 34391 34601
rect 34333 34592 34345 34595
rect 34020 34564 34345 34592
rect 34020 34552 34026 34564
rect 34333 34561 34345 34564
rect 34379 34561 34391 34595
rect 34333 34555 34391 34561
rect 34422 34552 34428 34604
rect 34480 34592 34486 34604
rect 35618 34592 35624 34604
rect 34480 34564 35480 34592
rect 35579 34564 35624 34592
rect 34480 34552 34486 34564
rect 15378 34524 15384 34536
rect 14844 34496 15384 34524
rect 9214 34456 9220 34468
rect 8312 34428 9220 34456
rect 5040 34416 5046 34428
rect 9214 34416 9220 34428
rect 9272 34416 9278 34468
rect 5166 34388 5172 34400
rect 5127 34360 5172 34388
rect 5166 34348 5172 34360
rect 5224 34348 5230 34400
rect 7006 34348 7012 34400
rect 7064 34388 7070 34400
rect 7193 34391 7251 34397
rect 7193 34388 7205 34391
rect 7064 34360 7205 34388
rect 7064 34348 7070 34360
rect 7193 34357 7205 34360
rect 7239 34357 7251 34391
rect 7193 34351 7251 34357
rect 9398 34348 9404 34400
rect 9456 34388 9462 34400
rect 9585 34391 9643 34397
rect 9585 34388 9597 34391
rect 9456 34360 9597 34388
rect 9456 34348 9462 34360
rect 9585 34357 9597 34360
rect 9631 34357 9643 34391
rect 9585 34351 9643 34357
rect 12434 34348 12440 34400
rect 12492 34388 12498 34400
rect 12897 34391 12955 34397
rect 12897 34388 12909 34391
rect 12492 34360 12909 34388
rect 12492 34348 12498 34360
rect 12897 34357 12909 34360
rect 12943 34388 12955 34391
rect 14292 34388 14320 34496
rect 15378 34484 15384 34496
rect 15436 34524 15442 34536
rect 15654 34524 15660 34536
rect 15436 34496 15660 34524
rect 15436 34484 15442 34496
rect 15654 34484 15660 34496
rect 15712 34484 15718 34536
rect 17037 34527 17095 34533
rect 17037 34524 17049 34527
rect 16316 34496 17049 34524
rect 16316 34465 16344 34496
rect 17037 34493 17049 34496
rect 17083 34493 17095 34527
rect 17037 34487 17095 34493
rect 17497 34527 17555 34533
rect 17497 34493 17509 34527
rect 17543 34524 17555 34527
rect 17954 34524 17960 34536
rect 17543 34496 17960 34524
rect 17543 34493 17555 34496
rect 17497 34487 17555 34493
rect 17954 34484 17960 34496
rect 18012 34524 18018 34536
rect 18874 34524 18880 34536
rect 18012 34496 18880 34524
rect 18012 34484 18018 34496
rect 18874 34484 18880 34496
rect 18932 34484 18938 34536
rect 22002 34524 22008 34536
rect 21963 34496 22008 34524
rect 22002 34484 22008 34496
rect 22060 34484 22066 34536
rect 22557 34527 22615 34533
rect 22557 34524 22569 34527
rect 22112 34496 22569 34524
rect 16301 34459 16359 34465
rect 16301 34425 16313 34459
rect 16347 34425 16359 34459
rect 16301 34419 16359 34425
rect 20714 34416 20720 34468
rect 20772 34456 20778 34468
rect 22112 34456 22140 34496
rect 22557 34493 22569 34496
rect 22603 34493 22615 34527
rect 22557 34487 22615 34493
rect 23198 34484 23204 34536
rect 23256 34524 23262 34536
rect 24305 34527 24363 34533
rect 24305 34524 24317 34527
rect 23256 34496 24317 34524
rect 23256 34484 23262 34496
rect 24305 34493 24317 34496
rect 24351 34493 24363 34527
rect 26206 34496 26240 34536
rect 24305 34487 24363 34493
rect 26234 34484 26240 34496
rect 26292 34484 26298 34536
rect 29825 34527 29883 34533
rect 29825 34493 29837 34527
rect 29871 34524 29883 34527
rect 31018 34524 31024 34536
rect 29871 34496 31024 34524
rect 29871 34493 29883 34496
rect 29825 34487 29883 34493
rect 31018 34484 31024 34496
rect 31076 34524 31082 34536
rect 31202 34524 31208 34536
rect 31076 34496 31208 34524
rect 31076 34484 31082 34496
rect 31202 34484 31208 34496
rect 31260 34484 31266 34536
rect 32398 34484 32404 34536
rect 32456 34524 32462 34536
rect 35342 34524 35348 34536
rect 32456 34496 35348 34524
rect 32456 34484 32462 34496
rect 35342 34484 35348 34496
rect 35400 34484 35406 34536
rect 35452 34524 35480 34564
rect 35618 34552 35624 34564
rect 35676 34552 35682 34604
rect 36464 34601 36492 34632
rect 37660 34604 37688 34632
rect 38556 34629 38568 34663
rect 38602 34660 38614 34663
rect 38746 34660 38752 34672
rect 38602 34632 38752 34660
rect 38602 34629 38614 34632
rect 38556 34623 38614 34629
rect 38746 34620 38752 34632
rect 38804 34620 38810 34672
rect 36449 34595 36507 34601
rect 36449 34561 36461 34595
rect 36495 34561 36507 34595
rect 36449 34555 36507 34561
rect 36725 34595 36783 34601
rect 36725 34561 36737 34595
rect 36771 34561 36783 34595
rect 36725 34555 36783 34561
rect 36541 34527 36599 34533
rect 36541 34524 36553 34527
rect 35452 34496 36553 34524
rect 36541 34493 36553 34496
rect 36587 34524 36599 34527
rect 36740 34524 36768 34555
rect 36814 34552 36820 34604
rect 36872 34592 36878 34604
rect 37461 34595 37519 34601
rect 37461 34592 37473 34595
rect 36872 34564 37473 34592
rect 36872 34552 36878 34564
rect 37461 34561 37473 34564
rect 37507 34561 37519 34595
rect 37642 34592 37648 34604
rect 37603 34564 37648 34592
rect 37461 34555 37519 34561
rect 37642 34552 37648 34564
rect 37700 34552 37706 34604
rect 39114 34592 39120 34604
rect 37936 34564 39120 34592
rect 37550 34524 37556 34536
rect 36587 34496 36676 34524
rect 36740 34496 37556 34524
rect 36587 34493 36599 34496
rect 36541 34487 36599 34493
rect 34698 34456 34704 34468
rect 20772 34428 22140 34456
rect 34659 34428 34704 34456
rect 20772 34416 20778 34428
rect 34698 34416 34704 34428
rect 34756 34416 34762 34468
rect 36648 34456 36676 34496
rect 37550 34484 37556 34496
rect 37608 34484 37614 34536
rect 37936 34524 37964 34564
rect 39114 34552 39120 34564
rect 39172 34552 39178 34604
rect 37660 34496 37964 34524
rect 37660 34456 37688 34496
rect 38010 34484 38016 34536
rect 38068 34524 38074 34536
rect 38289 34527 38347 34533
rect 38289 34524 38301 34527
rect 38068 34496 38301 34524
rect 38068 34484 38074 34496
rect 38289 34493 38301 34496
rect 38335 34493 38347 34527
rect 38289 34487 38347 34493
rect 36648 34428 37688 34456
rect 18414 34388 18420 34400
rect 12943 34360 14320 34388
rect 18375 34360 18420 34388
rect 12943 34357 12955 34360
rect 12897 34351 12955 34357
rect 18414 34348 18420 34360
rect 18472 34348 18478 34400
rect 27246 34348 27252 34400
rect 27304 34388 27310 34400
rect 27341 34391 27399 34397
rect 27341 34388 27353 34391
rect 27304 34360 27353 34388
rect 27304 34348 27310 34360
rect 27341 34357 27353 34360
rect 27387 34357 27399 34391
rect 27341 34351 27399 34357
rect 29733 34391 29791 34397
rect 29733 34357 29745 34391
rect 29779 34388 29791 34391
rect 30190 34388 30196 34400
rect 29779 34360 30196 34388
rect 29779 34357 29791 34360
rect 29733 34351 29791 34357
rect 30190 34348 30196 34360
rect 30248 34348 30254 34400
rect 39666 34388 39672 34400
rect 39627 34360 39672 34388
rect 39666 34348 39672 34360
rect 39724 34348 39730 34400
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 14090 34144 14096 34196
rect 14148 34184 14154 34196
rect 14461 34187 14519 34193
rect 14461 34184 14473 34187
rect 14148 34156 14473 34184
rect 14148 34144 14154 34156
rect 14461 34153 14473 34156
rect 14507 34153 14519 34187
rect 14461 34147 14519 34153
rect 17494 34144 17500 34196
rect 17552 34184 17558 34196
rect 18325 34187 18383 34193
rect 18325 34184 18337 34187
rect 17552 34156 18337 34184
rect 17552 34144 17558 34156
rect 18325 34153 18337 34156
rect 18371 34153 18383 34187
rect 18325 34147 18383 34153
rect 18874 34144 18880 34196
rect 18932 34184 18938 34196
rect 19797 34187 19855 34193
rect 19797 34184 19809 34187
rect 18932 34156 19809 34184
rect 18932 34144 18938 34156
rect 19797 34153 19809 34156
rect 19843 34153 19855 34187
rect 19797 34147 19855 34153
rect 20714 34144 20720 34196
rect 20772 34184 20778 34196
rect 20809 34187 20867 34193
rect 20809 34184 20821 34187
rect 20772 34156 20821 34184
rect 20772 34144 20778 34156
rect 20809 34153 20821 34156
rect 20855 34153 20867 34187
rect 20809 34147 20867 34153
rect 20993 34187 21051 34193
rect 20993 34153 21005 34187
rect 21039 34153 21051 34187
rect 27246 34184 27252 34196
rect 27207 34156 27252 34184
rect 20993 34147 21051 34153
rect 17770 34116 17776 34128
rect 16868 34088 17776 34116
rect 5166 34008 5172 34060
rect 5224 34008 5230 34060
rect 9398 34048 9404 34060
rect 9359 34020 9404 34048
rect 9398 34008 9404 34020
rect 9456 34008 9462 34060
rect 15378 34048 15384 34060
rect 15339 34020 15384 34048
rect 15378 34008 15384 34020
rect 15436 34008 15442 34060
rect 4154 33980 4160 33992
rect 4115 33952 4160 33980
rect 4154 33940 4160 33952
rect 4212 33940 4218 33992
rect 4424 33983 4482 33989
rect 4424 33949 4436 33983
rect 4470 33980 4482 33983
rect 5184 33980 5212 34008
rect 7006 33980 7012 33992
rect 4470 33952 5212 33980
rect 6967 33952 7012 33980
rect 4470 33949 4482 33952
rect 4424 33943 4482 33949
rect 7006 33940 7012 33952
rect 7064 33940 7070 33992
rect 7282 33980 7288 33992
rect 7243 33952 7288 33980
rect 7282 33940 7288 33952
rect 7340 33940 7346 33992
rect 8018 33980 8024 33992
rect 7979 33952 8024 33980
rect 8018 33940 8024 33952
rect 8076 33940 8082 33992
rect 9674 33989 9680 33992
rect 9668 33980 9680 33989
rect 9635 33952 9680 33980
rect 9668 33943 9680 33952
rect 9674 33940 9680 33943
rect 9732 33940 9738 33992
rect 12066 33980 12072 33992
rect 12027 33952 12072 33980
rect 12066 33940 12072 33952
rect 12124 33940 12130 33992
rect 12434 33940 12440 33992
rect 12492 33980 12498 33992
rect 13541 33983 13599 33989
rect 13541 33980 13553 33983
rect 12492 33952 13553 33980
rect 12492 33940 12498 33952
rect 13541 33949 13553 33952
rect 13587 33949 13599 33983
rect 13541 33943 13599 33949
rect 14277 33983 14335 33989
rect 14277 33949 14289 33983
rect 14323 33949 14335 33983
rect 14277 33943 14335 33949
rect 14461 33983 14519 33989
rect 14461 33949 14473 33983
rect 14507 33980 14519 33983
rect 16868 33980 16896 34088
rect 17770 34076 17776 34088
rect 17828 34076 17834 34128
rect 18138 34076 18144 34128
rect 18196 34116 18202 34128
rect 19242 34116 19248 34128
rect 18196 34088 19248 34116
rect 18196 34076 18202 34088
rect 19242 34076 19248 34088
rect 19300 34116 19306 34128
rect 19300 34088 19840 34116
rect 19300 34076 19306 34088
rect 18414 34048 18420 34060
rect 17420 34020 18420 34048
rect 17420 33989 17448 34020
rect 18414 34008 18420 34020
rect 18472 34008 18478 34060
rect 19334 34008 19340 34060
rect 19392 34048 19398 34060
rect 19613 34051 19671 34057
rect 19613 34048 19625 34051
rect 19392 34020 19625 34048
rect 19392 34008 19398 34020
rect 19613 34017 19625 34020
rect 19659 34017 19671 34051
rect 19613 34011 19671 34017
rect 14507 33952 16896 33980
rect 17405 33983 17463 33989
rect 14507 33949 14519 33952
rect 14461 33943 14519 33949
rect 17405 33949 17417 33983
rect 17451 33949 17463 33983
rect 17405 33943 17463 33949
rect 7193 33915 7251 33921
rect 7193 33881 7205 33915
rect 7239 33912 7251 33915
rect 7742 33912 7748 33924
rect 7239 33884 7748 33912
rect 7239 33881 7251 33884
rect 7193 33875 7251 33881
rect 7742 33872 7748 33884
rect 7800 33872 7806 33924
rect 14292 33912 14320 33943
rect 17494 33940 17500 33992
rect 17552 33980 17558 33992
rect 17770 33989 17776 33992
rect 17727 33983 17776 33989
rect 17552 33952 17597 33980
rect 17552 33940 17558 33952
rect 17727 33949 17739 33983
rect 17773 33949 17776 33983
rect 17727 33943 17776 33949
rect 17770 33940 17776 33943
rect 17828 33940 17834 33992
rect 17865 33983 17923 33989
rect 17865 33949 17877 33983
rect 17911 33982 17923 33983
rect 17911 33954 18000 33982
rect 18506 33980 18512 33992
rect 17911 33949 17923 33954
rect 17865 33943 17923 33949
rect 13464 33884 14320 33912
rect 15648 33915 15706 33921
rect 5258 33804 5264 33856
rect 5316 33844 5322 33856
rect 5537 33847 5595 33853
rect 5537 33844 5549 33847
rect 5316 33816 5549 33844
rect 5316 33804 5322 33816
rect 5537 33813 5549 33816
rect 5583 33813 5595 33847
rect 6822 33844 6828 33856
rect 6783 33816 6828 33844
rect 5537 33807 5595 33813
rect 6822 33804 6828 33816
rect 6880 33804 6886 33856
rect 7374 33804 7380 33856
rect 7432 33844 7438 33856
rect 7837 33847 7895 33853
rect 7837 33844 7849 33847
rect 7432 33816 7849 33844
rect 7432 33804 7438 33816
rect 7837 33813 7849 33816
rect 7883 33813 7895 33847
rect 7837 33807 7895 33813
rect 10318 33804 10324 33856
rect 10376 33844 10382 33856
rect 10781 33847 10839 33853
rect 10781 33844 10793 33847
rect 10376 33816 10793 33844
rect 10376 33804 10382 33816
rect 10781 33813 10793 33816
rect 10827 33813 10839 33847
rect 12250 33844 12256 33856
rect 12211 33816 12256 33844
rect 10781 33807 10839 33813
rect 12250 33804 12256 33816
rect 12308 33804 12314 33856
rect 12342 33804 12348 33856
rect 12400 33844 12406 33856
rect 13464 33853 13492 33884
rect 15648 33881 15660 33915
rect 15694 33912 15706 33915
rect 17221 33915 17279 33921
rect 17221 33912 17233 33915
rect 15694 33884 17233 33912
rect 15694 33881 15706 33884
rect 15648 33875 15706 33881
rect 17221 33881 17233 33884
rect 17267 33881 17279 33915
rect 17221 33875 17279 33881
rect 17310 33872 17316 33924
rect 17368 33912 17374 33924
rect 17589 33915 17647 33921
rect 17589 33912 17601 33915
rect 17368 33884 17601 33912
rect 17368 33872 17374 33884
rect 17589 33881 17601 33884
rect 17635 33881 17647 33915
rect 17589 33875 17647 33881
rect 17972 33912 18000 33954
rect 18467 33952 18512 33980
rect 18506 33940 18512 33952
rect 18564 33940 18570 33992
rect 18782 33980 18788 33992
rect 18743 33952 18788 33980
rect 18782 33940 18788 33952
rect 18840 33940 18846 33992
rect 19426 33980 19432 33992
rect 19387 33952 19432 33980
rect 19426 33940 19432 33952
rect 19484 33940 19490 33992
rect 19705 33983 19763 33989
rect 19705 33949 19717 33983
rect 19751 33949 19763 33983
rect 19812 33980 19840 34088
rect 21008 34048 21036 34147
rect 27246 34144 27252 34156
rect 27304 34144 27310 34196
rect 27614 34184 27620 34196
rect 27575 34156 27620 34184
rect 27614 34144 27620 34156
rect 27672 34144 27678 34196
rect 31202 34144 31208 34196
rect 31260 34184 31266 34196
rect 31260 34156 35894 34184
rect 31260 34144 31266 34156
rect 25682 34076 25688 34128
rect 25740 34116 25746 34128
rect 27798 34116 27804 34128
rect 25740 34088 27804 34116
rect 25740 34076 25746 34088
rect 27798 34076 27804 34088
rect 27856 34076 27862 34128
rect 35434 34116 35440 34128
rect 35395 34088 35440 34116
rect 35434 34076 35440 34088
rect 35492 34076 35498 34128
rect 35526 34076 35532 34128
rect 35584 34076 35590 34128
rect 35866 34116 35894 34156
rect 36262 34144 36268 34196
rect 36320 34184 36326 34196
rect 36357 34187 36415 34193
rect 36357 34184 36369 34187
rect 36320 34156 36369 34184
rect 36320 34144 36326 34156
rect 36357 34153 36369 34156
rect 36403 34153 36415 34187
rect 36357 34147 36415 34153
rect 37550 34144 37556 34196
rect 37608 34184 37614 34196
rect 37645 34187 37703 34193
rect 37645 34184 37657 34187
rect 37608 34156 37657 34184
rect 37608 34144 37614 34156
rect 37645 34153 37657 34156
rect 37691 34153 37703 34187
rect 39206 34184 39212 34196
rect 37645 34147 37703 34153
rect 37844 34156 39212 34184
rect 37844 34116 37872 34156
rect 39206 34144 39212 34156
rect 39264 34184 39270 34196
rect 40310 34184 40316 34196
rect 39264 34156 40316 34184
rect 39264 34144 39270 34156
rect 40310 34144 40316 34156
rect 40368 34144 40374 34196
rect 39022 34116 39028 34128
rect 35866 34088 37872 34116
rect 26602 34048 26608 34060
rect 20180 34020 21036 34048
rect 26252 34020 26608 34048
rect 20180 33992 20208 34020
rect 19889 33983 19947 33989
rect 19889 33980 19901 33983
rect 19812 33952 19901 33980
rect 19705 33943 19763 33949
rect 19889 33949 19901 33952
rect 19935 33949 19947 33983
rect 19889 33943 19947 33949
rect 19720 33912 19748 33943
rect 20162 33940 20168 33992
rect 20220 33940 20226 33992
rect 22002 33980 22008 33992
rect 21008 33952 22008 33980
rect 21008 33912 21036 33952
rect 22002 33940 22008 33952
rect 22060 33940 22066 33992
rect 23474 33940 23480 33992
rect 23532 33980 23538 33992
rect 26252 33989 26280 34020
rect 26602 34008 26608 34020
rect 26660 34048 26666 34060
rect 27246 34048 27252 34060
rect 26660 34020 27252 34048
rect 26660 34008 26666 34020
rect 27246 34008 27252 34020
rect 27304 34008 27310 34060
rect 32398 34048 32404 34060
rect 32359 34020 32404 34048
rect 32398 34008 32404 34020
rect 32456 34008 32462 34060
rect 35544 34048 35572 34076
rect 35360 34020 35572 34048
rect 36541 34051 36599 34057
rect 26237 33983 26295 33989
rect 26237 33980 26249 33983
rect 23532 33952 26249 33980
rect 23532 33940 23538 33952
rect 26237 33949 26249 33952
rect 26283 33949 26295 33983
rect 27154 33980 27160 33992
rect 27115 33952 27160 33980
rect 26237 33943 26295 33949
rect 27154 33940 27160 33952
rect 27212 33940 27218 33992
rect 27430 33980 27436 33992
rect 27391 33952 27436 33980
rect 27430 33940 27436 33952
rect 27488 33940 27494 33992
rect 30098 33980 30104 33992
rect 30059 33952 30104 33980
rect 30098 33940 30104 33952
rect 30156 33940 30162 33992
rect 30190 33940 30196 33992
rect 30248 33980 30254 33992
rect 30285 33983 30343 33989
rect 30285 33980 30297 33983
rect 30248 33952 30297 33980
rect 30248 33940 30254 33952
rect 30285 33949 30297 33952
rect 30331 33949 30343 33983
rect 30285 33943 30343 33949
rect 30374 33940 30380 33992
rect 30432 33980 30438 33992
rect 30432 33952 30477 33980
rect 30432 33940 30438 33952
rect 34790 33940 34796 33992
rect 34848 33980 34854 33992
rect 35360 33989 35388 34020
rect 36541 34017 36553 34051
rect 36587 34048 36599 34051
rect 36998 34048 37004 34060
rect 36587 34020 37004 34048
rect 36587 34017 36599 34020
rect 36541 34011 36599 34017
rect 36998 34008 37004 34020
rect 37056 34008 37062 34060
rect 35161 33983 35219 33989
rect 35161 33980 35173 33983
rect 34848 33952 35173 33980
rect 34848 33940 34854 33952
rect 35161 33949 35173 33952
rect 35207 33949 35219 33983
rect 35161 33943 35219 33949
rect 35345 33983 35403 33989
rect 35345 33949 35357 33983
rect 35391 33949 35403 33983
rect 35345 33943 35403 33949
rect 35529 33983 35587 33989
rect 35529 33949 35541 33983
rect 35575 33949 35587 33983
rect 35529 33943 35587 33949
rect 35621 33983 35679 33989
rect 35621 33949 35633 33983
rect 35667 33980 35679 33983
rect 36262 33980 36268 33992
rect 35667 33952 36268 33980
rect 35667 33949 35679 33952
rect 35621 33943 35679 33949
rect 21174 33912 21180 33924
rect 17972 33884 19748 33912
rect 20180 33884 21036 33912
rect 21135 33884 21180 33912
rect 13449 33847 13507 33853
rect 13449 33844 13461 33847
rect 12400 33816 13461 33844
rect 12400 33804 12406 33816
rect 13449 33813 13461 33816
rect 13495 33813 13507 33847
rect 13449 33807 13507 33813
rect 16761 33847 16819 33853
rect 16761 33813 16773 33847
rect 16807 33844 16819 33847
rect 17770 33844 17776 33856
rect 16807 33816 17776 33844
rect 16807 33813 16819 33816
rect 16761 33807 16819 33813
rect 17770 33804 17776 33816
rect 17828 33844 17834 33856
rect 17972 33844 18000 33884
rect 18690 33844 18696 33856
rect 17828 33816 18000 33844
rect 18651 33816 18696 33844
rect 17828 33804 17834 33816
rect 18690 33804 18696 33816
rect 18748 33804 18754 33856
rect 20180 33853 20208 33884
rect 21174 33872 21180 33884
rect 21232 33872 21238 33924
rect 26053 33915 26111 33921
rect 26053 33881 26065 33915
rect 26099 33912 26111 33915
rect 27172 33912 27200 33940
rect 26099 33884 27200 33912
rect 32668 33915 32726 33921
rect 26099 33881 26111 33884
rect 26053 33875 26111 33881
rect 32668 33881 32680 33915
rect 32714 33912 32726 33915
rect 32766 33912 32772 33924
rect 32714 33884 32772 33912
rect 32714 33881 32726 33884
rect 32668 33875 32726 33881
rect 32766 33872 32772 33884
rect 32824 33872 32830 33924
rect 35544 33912 35572 33943
rect 36262 33940 36268 33952
rect 36320 33940 36326 33992
rect 37844 33989 37872 34088
rect 38120 34088 39028 34116
rect 38120 33989 38148 34088
rect 39022 34076 39028 34088
rect 39080 34116 39086 34128
rect 39942 34116 39948 34128
rect 39080 34088 39948 34116
rect 39080 34076 39086 34088
rect 39942 34076 39948 34088
rect 40000 34076 40006 34128
rect 38746 34048 38752 34060
rect 38707 34020 38752 34048
rect 38746 34008 38752 34020
rect 38804 34008 38810 34060
rect 39206 34048 39212 34060
rect 39119 34020 39212 34048
rect 39206 34008 39212 34020
rect 39264 34048 39270 34060
rect 39666 34048 39672 34060
rect 39264 34020 39672 34048
rect 39264 34008 39270 34020
rect 39666 34008 39672 34020
rect 39724 34008 39730 34060
rect 37829 33983 37887 33989
rect 37829 33949 37841 33983
rect 37875 33949 37887 33983
rect 37829 33943 37887 33949
rect 38105 33983 38163 33989
rect 38105 33949 38117 33983
rect 38151 33949 38163 33983
rect 38105 33943 38163 33949
rect 38289 33983 38347 33989
rect 38289 33949 38301 33983
rect 38335 33949 38347 33983
rect 38930 33980 38936 33992
rect 38891 33952 38936 33980
rect 38289 33943 38347 33949
rect 36170 33912 36176 33924
rect 35544 33884 36176 33912
rect 36170 33872 36176 33884
rect 36228 33872 36234 33924
rect 36372 33884 37320 33912
rect 20990 33853 20996 33856
rect 20165 33847 20223 33853
rect 20165 33813 20177 33847
rect 20211 33813 20223 33847
rect 20165 33807 20223 33813
rect 20977 33847 20996 33853
rect 20977 33813 20989 33847
rect 20977 33807 20996 33813
rect 20990 33804 20996 33807
rect 21048 33804 21054 33856
rect 25590 33804 25596 33856
rect 25648 33844 25654 33856
rect 25869 33847 25927 33853
rect 25869 33844 25881 33847
rect 25648 33816 25881 33844
rect 25648 33804 25654 33816
rect 25869 33813 25881 33816
rect 25915 33813 25927 33847
rect 25869 33807 25927 33813
rect 29917 33847 29975 33853
rect 29917 33813 29929 33847
rect 29963 33844 29975 33847
rect 30006 33844 30012 33856
rect 29963 33816 30012 33844
rect 29963 33813 29975 33816
rect 29917 33807 29975 33813
rect 30006 33804 30012 33816
rect 30064 33804 30070 33856
rect 33410 33804 33416 33856
rect 33468 33844 33474 33856
rect 33781 33847 33839 33853
rect 33781 33844 33793 33847
rect 33468 33816 33793 33844
rect 33468 33804 33474 33816
rect 33781 33813 33793 33816
rect 33827 33813 33839 33847
rect 33781 33807 33839 33813
rect 35805 33847 35863 33853
rect 35805 33813 35817 33847
rect 35851 33844 35863 33847
rect 36372 33844 36400 33884
rect 36538 33844 36544 33856
rect 35851 33816 36400 33844
rect 36499 33816 36544 33844
rect 35851 33813 35863 33816
rect 35805 33807 35863 33813
rect 36538 33804 36544 33816
rect 36596 33804 36602 33856
rect 37292 33844 37320 33884
rect 37366 33872 37372 33924
rect 37424 33912 37430 33924
rect 38304 33912 38332 33943
rect 38930 33940 38936 33952
rect 38988 33940 38994 33992
rect 39114 33940 39120 33992
rect 39172 33980 39178 33992
rect 40402 33980 40408 33992
rect 39172 33952 40408 33980
rect 39172 33940 39178 33952
rect 40402 33940 40408 33952
rect 40460 33940 40466 33992
rect 37424 33884 38332 33912
rect 37424 33872 37430 33884
rect 37734 33844 37740 33856
rect 37292 33816 37740 33844
rect 37734 33804 37740 33816
rect 37792 33804 37798 33856
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 4154 33600 4160 33652
rect 4212 33640 4218 33652
rect 4341 33643 4399 33649
rect 4341 33640 4353 33643
rect 4212 33612 4353 33640
rect 4212 33600 4218 33612
rect 4341 33609 4353 33612
rect 4387 33609 4399 33643
rect 4341 33603 4399 33609
rect 5445 33643 5503 33649
rect 5445 33609 5457 33643
rect 5491 33640 5503 33643
rect 5902 33640 5908 33652
rect 5491 33612 5908 33640
rect 5491 33609 5503 33612
rect 5445 33603 5503 33609
rect 5902 33600 5908 33612
rect 5960 33600 5966 33652
rect 6917 33643 6975 33649
rect 6917 33609 6929 33643
rect 6963 33609 6975 33643
rect 6917 33603 6975 33609
rect 9677 33643 9735 33649
rect 9677 33609 9689 33643
rect 9723 33640 9735 33643
rect 9766 33640 9772 33652
rect 9723 33612 9772 33640
rect 9723 33609 9735 33612
rect 9677 33603 9735 33609
rect 6932 33572 6960 33603
rect 9766 33600 9772 33612
rect 9824 33600 9830 33652
rect 18782 33600 18788 33652
rect 18840 33640 18846 33652
rect 19429 33643 19487 33649
rect 19429 33640 19441 33643
rect 18840 33612 19441 33640
rect 18840 33600 18846 33612
rect 19429 33609 19441 33612
rect 19475 33609 19487 33643
rect 21174 33640 21180 33652
rect 21135 33612 21180 33640
rect 19429 33603 19487 33609
rect 21174 33600 21180 33612
rect 21232 33600 21238 33652
rect 27154 33600 27160 33652
rect 27212 33600 27218 33652
rect 27430 33600 27436 33652
rect 27488 33640 27494 33652
rect 28077 33643 28135 33649
rect 28077 33640 28089 33643
rect 27488 33612 28089 33640
rect 27488 33600 27494 33612
rect 28077 33609 28089 33612
rect 28123 33609 28135 33643
rect 28077 33603 28135 33609
rect 30098 33600 30104 33652
rect 30156 33640 30162 33652
rect 30561 33643 30619 33649
rect 30561 33640 30573 33643
rect 30156 33612 30573 33640
rect 30156 33600 30162 33612
rect 30561 33609 30573 33612
rect 30607 33609 30619 33643
rect 32766 33640 32772 33652
rect 32727 33612 32772 33640
rect 30561 33603 30619 33609
rect 32766 33600 32772 33612
rect 32824 33600 32830 33652
rect 7622 33575 7680 33581
rect 7622 33572 7634 33575
rect 6932 33544 7634 33572
rect 7622 33541 7634 33544
rect 7668 33541 7680 33575
rect 7622 33535 7680 33541
rect 7742 33532 7748 33584
rect 7800 33572 7806 33584
rect 10229 33575 10287 33581
rect 10229 33572 10241 33575
rect 7800 33544 10241 33572
rect 7800 33532 7806 33544
rect 10229 33541 10241 33544
rect 10275 33541 10287 33575
rect 10229 33535 10287 33541
rect 12250 33532 12256 33584
rect 12308 33572 12314 33584
rect 12814 33575 12872 33581
rect 12814 33572 12826 33575
rect 12308 33544 12826 33572
rect 12308 33532 12314 33544
rect 12814 33541 12826 33544
rect 12860 33541 12872 33575
rect 17770 33572 17776 33584
rect 12814 33535 12872 33541
rect 17144 33544 17776 33572
rect 4525 33507 4583 33513
rect 4525 33473 4537 33507
rect 4571 33504 4583 33507
rect 4798 33504 4804 33516
rect 4571 33476 4804 33504
rect 4571 33473 4583 33476
rect 4525 33467 4583 33473
rect 4798 33464 4804 33476
rect 4856 33464 4862 33516
rect 4982 33504 4988 33516
rect 4943 33476 4988 33504
rect 4982 33464 4988 33476
rect 5040 33464 5046 33516
rect 6733 33507 6791 33513
rect 6733 33473 6745 33507
rect 6779 33504 6791 33507
rect 7190 33504 7196 33516
rect 6779 33476 7196 33504
rect 6779 33473 6791 33476
rect 6733 33467 6791 33473
rect 7190 33464 7196 33476
rect 7248 33464 7254 33516
rect 7374 33504 7380 33516
rect 7335 33476 7380 33504
rect 7374 33464 7380 33476
rect 7432 33464 7438 33516
rect 9214 33504 9220 33516
rect 9175 33476 9220 33504
rect 9214 33464 9220 33476
rect 9272 33464 9278 33516
rect 10318 33504 10324 33516
rect 10279 33476 10324 33504
rect 10318 33464 10324 33476
rect 10376 33464 10382 33516
rect 13081 33507 13139 33513
rect 13081 33473 13093 33507
rect 13127 33504 13139 33507
rect 13170 33504 13176 33516
rect 13127 33476 13176 33504
rect 13127 33473 13139 33476
rect 13081 33467 13139 33473
rect 13170 33464 13176 33476
rect 13228 33504 13234 33516
rect 13722 33504 13728 33516
rect 13228 33476 13728 33504
rect 13228 33464 13234 33476
rect 13722 33464 13728 33476
rect 13780 33464 13786 33516
rect 17144 33513 17172 33544
rect 17770 33532 17776 33544
rect 17828 33532 17834 33584
rect 17957 33575 18015 33581
rect 17957 33541 17969 33575
rect 18003 33572 18015 33575
rect 18138 33572 18144 33584
rect 18003 33544 18144 33572
rect 18003 33541 18015 33544
rect 17957 33535 18015 33541
rect 17129 33507 17187 33513
rect 17129 33473 17141 33507
rect 17175 33473 17187 33507
rect 17129 33467 17187 33473
rect 17313 33507 17371 33513
rect 17313 33473 17325 33507
rect 17359 33504 17371 33507
rect 17972 33504 18000 33535
rect 18138 33532 18144 33544
rect 18196 33532 18202 33584
rect 20990 33572 20996 33584
rect 18800 33544 20996 33572
rect 17359 33476 18000 33504
rect 17359 33473 17371 33476
rect 17313 33467 17371 33473
rect 18046 33464 18052 33516
rect 18104 33504 18110 33516
rect 18506 33504 18512 33516
rect 18104 33476 18512 33504
rect 18104 33464 18110 33476
rect 18506 33464 18512 33476
rect 18564 33504 18570 33516
rect 18800 33513 18828 33544
rect 20990 33532 20996 33544
rect 21048 33532 21054 33584
rect 25590 33572 25596 33584
rect 25551 33544 25596 33572
rect 25590 33532 25596 33544
rect 25648 33532 25654 33584
rect 25682 33532 25688 33584
rect 25740 33572 25746 33584
rect 27172 33572 27200 33600
rect 25740 33544 25785 33572
rect 26436 33544 27200 33572
rect 27341 33575 27399 33581
rect 25740 33532 25746 33544
rect 18693 33507 18751 33513
rect 18693 33504 18705 33507
rect 18564 33476 18705 33504
rect 18564 33464 18570 33476
rect 18693 33473 18705 33476
rect 18739 33473 18751 33507
rect 18693 33467 18751 33473
rect 18785 33507 18843 33513
rect 18785 33473 18797 33507
rect 18831 33473 18843 33507
rect 18785 33467 18843 33473
rect 18877 33507 18935 33513
rect 18877 33473 18889 33507
rect 18923 33473 18935 33507
rect 18877 33467 18935 33473
rect 17678 33396 17684 33448
rect 17736 33436 17742 33448
rect 18892 33436 18920 33467
rect 19334 33464 19340 33516
rect 19392 33504 19398 33516
rect 19613 33507 19671 33513
rect 19613 33504 19625 33507
rect 19392 33476 19625 33504
rect 19392 33464 19398 33476
rect 19613 33473 19625 33476
rect 19659 33473 19671 33507
rect 19613 33467 19671 33473
rect 19702 33464 19708 33516
rect 19760 33504 19766 33516
rect 20162 33504 20168 33516
rect 19760 33476 19805 33504
rect 20123 33476 20168 33504
rect 19760 33464 19766 33476
rect 20162 33464 20168 33476
rect 20220 33464 20226 33516
rect 20349 33507 20407 33513
rect 20349 33473 20361 33507
rect 20395 33504 20407 33507
rect 20438 33504 20444 33516
rect 20395 33476 20444 33504
rect 20395 33473 20407 33476
rect 20349 33467 20407 33473
rect 20438 33464 20444 33476
rect 20496 33464 20502 33516
rect 21082 33504 21088 33516
rect 21043 33476 21088 33504
rect 21082 33464 21088 33476
rect 21140 33464 21146 33516
rect 21266 33504 21272 33516
rect 21227 33476 21272 33504
rect 21266 33464 21272 33476
rect 21324 33464 21330 33516
rect 24673 33507 24731 33513
rect 24673 33473 24685 33507
rect 24719 33504 24731 33507
rect 24854 33504 24860 33516
rect 24719 33476 24860 33504
rect 24719 33473 24731 33476
rect 24673 33467 24731 33473
rect 24854 33464 24860 33476
rect 24912 33464 24918 33516
rect 25501 33507 25559 33513
rect 25501 33473 25513 33507
rect 25547 33504 25559 33507
rect 25774 33504 25780 33516
rect 25832 33513 25838 33516
rect 26436 33513 26464 33544
rect 27341 33541 27353 33575
rect 27387 33572 27399 33575
rect 28718 33572 28724 33584
rect 27387 33544 28724 33572
rect 27387 33541 27399 33544
rect 27341 33535 27399 33541
rect 25832 33507 25861 33513
rect 25547 33476 25636 33504
rect 25547 33473 25559 33476
rect 25501 33467 25559 33473
rect 17736 33408 18920 33436
rect 19429 33439 19487 33445
rect 17736 33396 17742 33408
rect 19429 33405 19441 33439
rect 19475 33436 19487 33439
rect 20898 33436 20904 33448
rect 19475 33408 20904 33436
rect 19475 33405 19487 33408
rect 19429 33399 19487 33405
rect 20898 33396 20904 33408
rect 20956 33396 20962 33448
rect 23842 33436 23848 33448
rect 23803 33408 23848 33436
rect 23842 33396 23848 33408
rect 23900 33396 23906 33448
rect 17954 33328 17960 33380
rect 18012 33368 18018 33380
rect 18506 33368 18512 33380
rect 18012 33340 18512 33368
rect 18012 33328 18018 33340
rect 18506 33328 18512 33340
rect 18564 33328 18570 33380
rect 18690 33328 18696 33380
rect 18748 33368 18754 33380
rect 20257 33371 20315 33377
rect 20257 33368 20269 33371
rect 18748 33340 20269 33368
rect 18748 33328 18754 33340
rect 20257 33337 20269 33340
rect 20303 33337 20315 33371
rect 20257 33331 20315 33337
rect 24670 33328 24676 33380
rect 24728 33368 24734 33380
rect 25608 33368 25636 33476
rect 25700 33476 25780 33504
rect 25700 33448 25728 33476
rect 25774 33464 25780 33476
rect 25849 33504 25861 33507
rect 25961 33507 26019 33513
rect 25849 33476 25925 33504
rect 25849 33473 25861 33476
rect 25832 33467 25861 33473
rect 25961 33473 25973 33507
rect 26007 33504 26019 33507
rect 26421 33507 26479 33513
rect 26007 33476 26234 33504
rect 26007 33473 26019 33476
rect 25961 33467 26019 33473
rect 25832 33464 25838 33467
rect 25682 33396 25688 33448
rect 25740 33396 25746 33448
rect 26206 33436 26234 33476
rect 26421 33473 26433 33507
rect 26467 33473 26479 33507
rect 26602 33504 26608 33516
rect 26563 33476 26608 33504
rect 26421 33467 26479 33473
rect 26602 33464 26608 33476
rect 26660 33464 26666 33516
rect 27157 33507 27215 33513
rect 27157 33473 27169 33507
rect 27203 33504 27215 33507
rect 27246 33504 27252 33516
rect 27203 33476 27252 33504
rect 27203 33473 27215 33476
rect 27157 33467 27215 33473
rect 27246 33464 27252 33476
rect 27304 33464 27310 33516
rect 28184 33513 28212 33544
rect 28718 33532 28724 33544
rect 28776 33532 28782 33584
rect 30742 33572 30748 33584
rect 30116 33544 30748 33572
rect 30116 33513 30144 33544
rect 30742 33532 30748 33544
rect 30800 33532 30806 33584
rect 35434 33572 35440 33584
rect 35360 33544 35440 33572
rect 27985 33507 28043 33513
rect 27985 33473 27997 33507
rect 28031 33473 28043 33507
rect 27985 33467 28043 33473
rect 28169 33507 28227 33513
rect 28169 33473 28181 33507
rect 28215 33504 28227 33507
rect 29917 33507 29975 33513
rect 28215 33476 28249 33504
rect 28215 33473 28227 33476
rect 28169 33467 28227 33473
rect 29917 33473 29929 33507
rect 29963 33473 29975 33507
rect 29917 33467 29975 33473
rect 30101 33507 30159 33513
rect 30101 33473 30113 33507
rect 30147 33473 30159 33507
rect 30101 33467 30159 33473
rect 30377 33507 30435 33513
rect 30377 33473 30389 33507
rect 30423 33504 30435 33507
rect 30466 33504 30472 33516
rect 30423 33476 30472 33504
rect 30423 33473 30435 33476
rect 30377 33467 30435 33473
rect 26326 33436 26332 33448
rect 26206 33408 26332 33436
rect 26326 33396 26332 33408
rect 26384 33436 26390 33448
rect 27264 33436 27292 33464
rect 28000 33436 28028 33467
rect 26384 33408 28028 33436
rect 26384 33396 26390 33408
rect 26513 33371 26571 33377
rect 26513 33368 26525 33371
rect 24728 33340 25452 33368
rect 25608 33340 26525 33368
rect 24728 33328 24734 33340
rect 5258 33300 5264 33312
rect 5219 33272 5264 33300
rect 5258 33260 5264 33272
rect 5316 33260 5322 33312
rect 8757 33303 8815 33309
rect 8757 33269 8769 33303
rect 8803 33300 8815 33303
rect 9309 33303 9367 33309
rect 9309 33300 9321 33303
rect 8803 33272 9321 33300
rect 8803 33269 8815 33272
rect 8757 33263 8815 33269
rect 9309 33269 9321 33272
rect 9355 33269 9367 33303
rect 11698 33300 11704 33312
rect 11659 33272 11704 33300
rect 9309 33263 9367 33269
rect 11698 33260 11704 33272
rect 11756 33260 11762 33312
rect 17218 33300 17224 33312
rect 17179 33272 17224 33300
rect 17218 33260 17224 33272
rect 17276 33260 17282 33312
rect 18138 33300 18144 33312
rect 18099 33272 18144 33300
rect 18138 33260 18144 33272
rect 18196 33260 18202 33312
rect 25222 33260 25228 33312
rect 25280 33300 25286 33312
rect 25317 33303 25375 33309
rect 25317 33300 25329 33303
rect 25280 33272 25329 33300
rect 25280 33260 25286 33272
rect 25317 33269 25329 33272
rect 25363 33269 25375 33303
rect 25424 33300 25452 33340
rect 26513 33337 26525 33340
rect 26559 33337 26571 33371
rect 29086 33368 29092 33380
rect 26513 33331 26571 33337
rect 27356 33340 29092 33368
rect 27356 33300 27384 33340
rect 29086 33328 29092 33340
rect 29144 33368 29150 33380
rect 29932 33368 29960 33467
rect 30466 33464 30472 33476
rect 30524 33504 30530 33516
rect 31202 33504 31208 33516
rect 30524 33476 31208 33504
rect 30524 33464 30530 33476
rect 31202 33464 31208 33476
rect 31260 33464 31266 33516
rect 32950 33504 32956 33516
rect 32911 33476 32956 33504
rect 32950 33464 32956 33476
rect 33008 33464 33014 33516
rect 35360 33513 35388 33544
rect 35434 33532 35440 33544
rect 35492 33532 35498 33584
rect 35345 33507 35403 33513
rect 35345 33473 35357 33507
rect 35391 33473 35403 33507
rect 46934 33504 46940 33516
rect 46895 33476 46940 33504
rect 35345 33467 35403 33473
rect 46934 33464 46940 33476
rect 46992 33464 46998 33516
rect 35437 33439 35495 33445
rect 35437 33405 35449 33439
rect 35483 33436 35495 33439
rect 36538 33436 36544 33448
rect 35483 33408 36544 33436
rect 35483 33405 35495 33408
rect 35437 33399 35495 33405
rect 36538 33396 36544 33408
rect 36596 33396 36602 33448
rect 29144 33340 29960 33368
rect 29144 33328 29150 33340
rect 34606 33328 34612 33380
rect 34664 33368 34670 33380
rect 34977 33371 35035 33377
rect 34977 33368 34989 33371
rect 34664 33340 34989 33368
rect 34664 33328 34670 33340
rect 34977 33337 34989 33340
rect 35023 33337 35035 33371
rect 46934 33368 46940 33380
rect 34977 33331 35035 33337
rect 45526 33340 46940 33368
rect 27522 33300 27528 33312
rect 25424 33272 27384 33300
rect 27483 33272 27528 33300
rect 25317 33263 25375 33269
rect 27522 33260 27528 33272
rect 27580 33260 27586 33312
rect 29638 33260 29644 33312
rect 29696 33300 29702 33312
rect 45526 33300 45554 33340
rect 46934 33328 46940 33340
rect 46992 33328 46998 33380
rect 47026 33300 47032 33312
rect 29696 33272 45554 33300
rect 46987 33272 47032 33300
rect 29696 33260 29702 33272
rect 47026 33260 47032 33272
rect 47084 33260 47090 33312
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 2682 33056 2688 33108
rect 2740 33096 2746 33108
rect 7377 33099 7435 33105
rect 2740 33068 7144 33096
rect 2740 33056 2746 33068
rect 4982 32988 4988 33040
rect 5040 33028 5046 33040
rect 5261 33031 5319 33037
rect 5261 33028 5273 33031
rect 5040 33000 5273 33028
rect 5040 32988 5046 33000
rect 5261 32997 5273 33000
rect 5307 32997 5319 33031
rect 5261 32991 5319 32997
rect 3786 32852 3792 32904
rect 3844 32892 3850 32904
rect 3973 32895 4031 32901
rect 3973 32892 3985 32895
rect 3844 32864 3985 32892
rect 3844 32852 3850 32864
rect 3973 32861 3985 32864
rect 4019 32861 4031 32895
rect 5994 32892 6000 32904
rect 5955 32864 6000 32892
rect 3973 32855 4031 32861
rect 5994 32852 6000 32864
rect 6052 32852 6058 32904
rect 6264 32895 6322 32901
rect 6264 32861 6276 32895
rect 6310 32892 6322 32895
rect 6822 32892 6828 32904
rect 6310 32864 6828 32892
rect 6310 32861 6322 32864
rect 6264 32855 6322 32861
rect 6822 32852 6828 32864
rect 6880 32852 6886 32904
rect 5442 32824 5448 32836
rect 5403 32796 5448 32824
rect 5442 32784 5448 32796
rect 5500 32784 5506 32836
rect 7116 32824 7144 33068
rect 7377 33065 7389 33099
rect 7423 33096 7435 33099
rect 8021 33099 8079 33105
rect 8021 33096 8033 33099
rect 7423 33068 8033 33096
rect 7423 33065 7435 33068
rect 7377 33059 7435 33065
rect 8021 33065 8033 33068
rect 8067 33065 8079 33099
rect 8021 33059 8079 33065
rect 20257 33099 20315 33105
rect 20257 33065 20269 33099
rect 20303 33096 20315 33099
rect 21082 33096 21088 33108
rect 20303 33068 21088 33096
rect 20303 33065 20315 33068
rect 20257 33059 20315 33065
rect 21082 33056 21088 33068
rect 21140 33056 21146 33108
rect 26326 33096 26332 33108
rect 26287 33068 26332 33096
rect 26326 33056 26332 33068
rect 26384 33056 26390 33108
rect 27154 33056 27160 33108
rect 27212 33096 27218 33108
rect 27433 33099 27491 33105
rect 27433 33096 27445 33099
rect 27212 33068 27445 33096
rect 27212 33056 27218 33068
rect 27433 33065 27445 33068
rect 27479 33065 27491 33099
rect 27433 33059 27491 33065
rect 30374 33056 30380 33108
rect 30432 33096 30438 33108
rect 31113 33099 31171 33105
rect 31113 33096 31125 33099
rect 30432 33068 31125 33096
rect 30432 33056 30438 33068
rect 31113 33065 31125 33068
rect 31159 33096 31171 33099
rect 31386 33096 31392 33108
rect 31159 33068 31392 33096
rect 31159 33065 31171 33068
rect 31113 33059 31171 33065
rect 31386 33056 31392 33068
rect 31444 33096 31450 33108
rect 31444 33068 31616 33096
rect 31444 33056 31450 33068
rect 7190 32988 7196 33040
rect 7248 33028 7254 33040
rect 7837 33031 7895 33037
rect 7837 33028 7849 33031
rect 7248 33000 7849 33028
rect 7248 32988 7254 33000
rect 7837 32997 7849 33000
rect 7883 32997 7895 33031
rect 7837 32991 7895 32997
rect 9398 32920 9404 32972
rect 9456 32960 9462 32972
rect 10321 32963 10379 32969
rect 10321 32960 10333 32963
rect 9456 32932 10333 32960
rect 9456 32920 9462 32932
rect 10321 32929 10333 32932
rect 10367 32929 10379 32963
rect 10321 32923 10379 32929
rect 12805 32963 12863 32969
rect 12805 32929 12817 32963
rect 12851 32960 12863 32963
rect 12851 32932 15332 32960
rect 12851 32929 12863 32932
rect 12805 32923 12863 32929
rect 8297 32895 8355 32901
rect 8297 32861 8309 32895
rect 8343 32892 8355 32895
rect 9214 32892 9220 32904
rect 8343 32864 9220 32892
rect 8343 32861 8355 32864
rect 8297 32855 8355 32861
rect 9214 32852 9220 32864
rect 9272 32852 9278 32904
rect 10137 32895 10195 32901
rect 10137 32861 10149 32895
rect 10183 32892 10195 32895
rect 11698 32892 11704 32904
rect 10183 32864 11704 32892
rect 10183 32861 10195 32864
rect 10137 32855 10195 32861
rect 11698 32852 11704 32864
rect 11756 32892 11762 32904
rect 12529 32895 12587 32901
rect 12529 32892 12541 32895
rect 11756 32864 12541 32892
rect 11756 32852 11762 32864
rect 12529 32861 12541 32864
rect 12575 32861 12587 32895
rect 12529 32855 12587 32861
rect 13725 32895 13783 32901
rect 13725 32861 13737 32895
rect 13771 32892 13783 32895
rect 14274 32892 14280 32904
rect 13771 32864 14280 32892
rect 13771 32861 13783 32864
rect 13725 32855 13783 32861
rect 14274 32852 14280 32864
rect 14332 32852 14338 32904
rect 15304 32892 15332 32932
rect 15378 32920 15384 32972
rect 15436 32960 15442 32972
rect 17589 32963 17647 32969
rect 17589 32960 17601 32963
rect 15436 32932 17601 32960
rect 15436 32920 15442 32932
rect 17589 32929 17601 32932
rect 17635 32929 17647 32963
rect 20717 32963 20775 32969
rect 20717 32960 20729 32963
rect 17589 32923 17647 32929
rect 20088 32932 20729 32960
rect 15562 32892 15568 32904
rect 15304 32864 15568 32892
rect 15562 32852 15568 32864
rect 15620 32852 15626 32904
rect 19242 32852 19248 32904
rect 19300 32892 19306 32904
rect 20088 32901 20116 32932
rect 20717 32929 20729 32932
rect 20763 32929 20775 32963
rect 20717 32923 20775 32929
rect 21085 32963 21143 32969
rect 21085 32929 21097 32963
rect 21131 32960 21143 32963
rect 21266 32960 21272 32972
rect 21131 32932 21272 32960
rect 21131 32929 21143 32932
rect 21085 32923 21143 32929
rect 21266 32920 21272 32932
rect 21324 32920 21330 32972
rect 22465 32963 22523 32969
rect 22465 32960 22477 32963
rect 21744 32932 22477 32960
rect 20073 32895 20131 32901
rect 20073 32892 20085 32895
rect 19300 32864 20085 32892
rect 19300 32852 19306 32864
rect 20073 32861 20085 32864
rect 20119 32861 20131 32895
rect 20073 32855 20131 32861
rect 20257 32895 20315 32901
rect 20257 32861 20269 32895
rect 20303 32861 20315 32895
rect 20257 32855 20315 32861
rect 20901 32895 20959 32901
rect 20901 32861 20913 32895
rect 20947 32861 20959 32895
rect 20901 32855 20959 32861
rect 12621 32827 12679 32833
rect 12621 32824 12633 32827
rect 7116 32796 12633 32824
rect 12621 32793 12633 32796
rect 12667 32824 12679 32827
rect 14826 32824 14832 32836
rect 12667 32796 14832 32824
rect 12667 32793 12679 32796
rect 12621 32787 12679 32793
rect 14826 32784 14832 32796
rect 14884 32784 14890 32836
rect 18322 32784 18328 32836
rect 18380 32824 18386 32836
rect 18417 32827 18475 32833
rect 18417 32824 18429 32827
rect 18380 32796 18429 32824
rect 18380 32784 18386 32796
rect 18417 32793 18429 32796
rect 18463 32793 18475 32827
rect 18417 32787 18475 32793
rect 19702 32784 19708 32836
rect 19760 32824 19766 32836
rect 20272 32824 20300 32855
rect 20916 32824 20944 32855
rect 21174 32852 21180 32904
rect 21232 32892 21238 32904
rect 21744 32901 21772 32932
rect 22465 32929 22477 32932
rect 22511 32929 22523 32963
rect 22465 32923 22523 32929
rect 22649 32963 22707 32969
rect 22649 32929 22661 32963
rect 22695 32929 22707 32963
rect 22649 32923 22707 32929
rect 21729 32895 21787 32901
rect 21729 32892 21741 32895
rect 21232 32864 21741 32892
rect 21232 32852 21238 32864
rect 21729 32861 21741 32864
rect 21775 32861 21787 32895
rect 21729 32855 21787 32861
rect 21818 32852 21824 32904
rect 21876 32892 21882 32904
rect 22373 32895 22431 32901
rect 22373 32892 22385 32895
rect 21876 32864 22385 32892
rect 21876 32852 21882 32864
rect 22373 32861 22385 32864
rect 22419 32861 22431 32895
rect 22664 32892 22692 32923
rect 23842 32920 23848 32972
rect 23900 32960 23906 32972
rect 24949 32963 25007 32969
rect 24949 32960 24961 32963
rect 23900 32932 24961 32960
rect 23900 32920 23906 32932
rect 24949 32929 24961 32932
rect 24995 32929 25007 32963
rect 27430 32960 27436 32972
rect 24949 32923 25007 32929
rect 27356 32932 27436 32960
rect 23937 32895 23995 32901
rect 23937 32892 23949 32895
rect 22664 32864 23949 32892
rect 22373 32855 22431 32861
rect 23937 32861 23949 32864
rect 23983 32892 23995 32895
rect 24026 32892 24032 32904
rect 23983 32864 24032 32892
rect 23983 32861 23995 32864
rect 23937 32855 23995 32861
rect 24026 32852 24032 32864
rect 24084 32852 24090 32904
rect 25222 32901 25228 32904
rect 25216 32892 25228 32901
rect 25183 32864 25228 32892
rect 25216 32855 25228 32864
rect 25222 32852 25228 32855
rect 25280 32852 25286 32904
rect 27356 32901 27384 32932
rect 27430 32920 27436 32932
rect 27488 32920 27494 32972
rect 28350 32920 28356 32972
rect 28408 32960 28414 32972
rect 29730 32960 29736 32972
rect 28408 32932 29736 32960
rect 28408 32920 28414 32932
rect 29730 32920 29736 32932
rect 29788 32920 29794 32972
rect 31588 32969 31616 33068
rect 32950 33056 32956 33108
rect 33008 33096 33014 33108
rect 33045 33099 33103 33105
rect 33045 33096 33057 33099
rect 33008 33068 33057 33096
rect 33008 33056 33014 33068
rect 33045 33065 33057 33068
rect 33091 33065 33103 33099
rect 40402 33096 40408 33108
rect 40363 33068 40408 33096
rect 33045 33059 33103 33065
rect 40402 33056 40408 33068
rect 40460 33056 40466 33108
rect 46750 33028 46756 33040
rect 45756 33000 46756 33028
rect 31573 32963 31631 32969
rect 31573 32929 31585 32963
rect 31619 32929 31631 32963
rect 31573 32923 31631 32929
rect 33689 32963 33747 32969
rect 33689 32929 33701 32963
rect 33735 32960 33747 32963
rect 35250 32960 35256 32972
rect 33735 32932 35256 32960
rect 33735 32929 33747 32932
rect 33689 32923 33747 32929
rect 35250 32920 35256 32932
rect 35308 32920 35314 32972
rect 27341 32895 27399 32901
rect 27341 32861 27353 32895
rect 27387 32861 27399 32895
rect 27522 32892 27528 32904
rect 27483 32864 27528 32892
rect 27341 32855 27399 32861
rect 27522 32852 27528 32864
rect 27580 32852 27586 32904
rect 30006 32901 30012 32904
rect 30000 32892 30012 32901
rect 29967 32864 30012 32892
rect 30000 32855 30012 32864
rect 30006 32852 30012 32855
rect 30064 32852 30070 32904
rect 31757 32895 31815 32901
rect 31757 32892 31769 32895
rect 31588 32864 31769 32892
rect 31588 32836 31616 32864
rect 31757 32861 31769 32864
rect 31803 32861 31815 32895
rect 33410 32892 33416 32904
rect 33371 32864 33416 32892
rect 31757 32855 31815 32861
rect 33410 32852 33416 32864
rect 33468 32852 33474 32904
rect 35345 32895 35403 32901
rect 35345 32861 35357 32895
rect 35391 32861 35403 32895
rect 35345 32855 35403 32861
rect 35529 32895 35587 32901
rect 35529 32861 35541 32895
rect 35575 32892 35587 32895
rect 36170 32892 36176 32904
rect 35575 32864 36176 32892
rect 35575 32861 35587 32864
rect 35529 32855 35587 32861
rect 23382 32824 23388 32836
rect 19760 32796 23388 32824
rect 19760 32784 19766 32796
rect 23382 32784 23388 32796
rect 23440 32784 23446 32836
rect 31570 32784 31576 32836
rect 31628 32784 31634 32836
rect 33134 32784 33140 32836
rect 33192 32824 33198 32836
rect 35360 32824 35388 32855
rect 36170 32852 36176 32864
rect 36228 32852 36234 32904
rect 38930 32892 38936 32904
rect 38891 32864 38936 32892
rect 38930 32852 38936 32864
rect 38988 32852 38994 32904
rect 39114 32892 39120 32904
rect 39075 32864 39120 32892
rect 39114 32852 39120 32864
rect 39172 32852 39178 32904
rect 40218 32892 40224 32904
rect 40179 32864 40224 32892
rect 40218 32852 40224 32864
rect 40276 32852 40282 32904
rect 40497 32895 40555 32901
rect 40497 32861 40509 32895
rect 40543 32892 40555 32895
rect 41322 32892 41328 32904
rect 40543 32864 41328 32892
rect 40543 32861 40555 32864
rect 40497 32855 40555 32861
rect 41322 32852 41328 32864
rect 41380 32852 41386 32904
rect 45756 32901 45784 33000
rect 46750 32988 46756 33000
rect 46808 33028 46814 33040
rect 47118 33028 47124 33040
rect 46808 33000 47124 33028
rect 46808 32988 46814 33000
rect 47118 32988 47124 33000
rect 47176 32988 47182 33040
rect 46661 32963 46719 32969
rect 46661 32929 46673 32963
rect 46707 32960 46719 32963
rect 47026 32960 47032 32972
rect 46707 32932 47032 32960
rect 46707 32929 46719 32932
rect 46661 32923 46719 32929
rect 47026 32920 47032 32932
rect 47084 32920 47090 32972
rect 45741 32895 45799 32901
rect 45741 32861 45753 32895
rect 45787 32861 45799 32895
rect 46474 32892 46480 32904
rect 46435 32864 46480 32892
rect 45741 32855 45799 32861
rect 46474 32852 46480 32864
rect 46532 32852 46538 32904
rect 36354 32824 36360 32836
rect 33192 32796 36360 32824
rect 33192 32784 33198 32796
rect 36354 32784 36360 32796
rect 36412 32784 36418 32836
rect 48314 32824 48320 32836
rect 48275 32796 48320 32824
rect 48314 32784 48320 32796
rect 48372 32784 48378 32836
rect 9766 32756 9772 32768
rect 9727 32728 9772 32756
rect 9766 32716 9772 32728
rect 9824 32716 9830 32768
rect 10229 32759 10287 32765
rect 10229 32725 10241 32759
rect 10275 32756 10287 32759
rect 10318 32756 10324 32768
rect 10275 32728 10324 32756
rect 10275 32725 10287 32728
rect 10229 32719 10287 32725
rect 10318 32716 10324 32728
rect 10376 32716 10382 32768
rect 12158 32756 12164 32768
rect 12119 32728 12164 32756
rect 12158 32716 12164 32728
rect 12216 32716 12222 32768
rect 13538 32756 13544 32768
rect 13499 32728 13544 32756
rect 13538 32716 13544 32728
rect 13596 32716 13602 32768
rect 20438 32716 20444 32768
rect 20496 32756 20502 32768
rect 21545 32759 21603 32765
rect 21545 32756 21557 32759
rect 20496 32728 21557 32756
rect 20496 32716 20502 32728
rect 21545 32725 21557 32728
rect 21591 32725 21603 32759
rect 21545 32719 21603 32725
rect 22186 32716 22192 32768
rect 22244 32756 22250 32768
rect 22649 32759 22707 32765
rect 22649 32756 22661 32759
rect 22244 32728 22661 32756
rect 22244 32716 22250 32728
rect 22649 32725 22661 32728
rect 22695 32725 22707 32759
rect 22649 32719 22707 32725
rect 23937 32759 23995 32765
rect 23937 32725 23949 32759
rect 23983 32756 23995 32759
rect 24118 32756 24124 32768
rect 23983 32728 24124 32756
rect 23983 32725 23995 32728
rect 23937 32719 23995 32725
rect 24118 32716 24124 32728
rect 24176 32756 24182 32768
rect 25222 32756 25228 32768
rect 24176 32728 25228 32756
rect 24176 32716 24182 32728
rect 25222 32716 25228 32728
rect 25280 32716 25286 32768
rect 31941 32759 31999 32765
rect 31941 32725 31953 32759
rect 31987 32756 31999 32759
rect 33042 32756 33048 32768
rect 31987 32728 33048 32756
rect 31987 32725 31999 32728
rect 31941 32719 31999 32725
rect 33042 32716 33048 32728
rect 33100 32716 33106 32768
rect 33505 32759 33563 32765
rect 33505 32725 33517 32759
rect 33551 32756 33563 32759
rect 33594 32756 33600 32768
rect 33551 32728 33600 32756
rect 33551 32725 33563 32728
rect 33505 32719 33563 32725
rect 33594 32716 33600 32728
rect 33652 32716 33658 32768
rect 35437 32759 35495 32765
rect 35437 32725 35449 32759
rect 35483 32756 35495 32759
rect 35526 32756 35532 32768
rect 35483 32728 35532 32756
rect 35483 32725 35495 32728
rect 35437 32719 35495 32725
rect 35526 32716 35532 32728
rect 35584 32716 35590 32768
rect 37826 32716 37832 32768
rect 37884 32756 37890 32768
rect 38933 32759 38991 32765
rect 38933 32756 38945 32759
rect 37884 32728 38945 32756
rect 37884 32716 37890 32728
rect 38933 32725 38945 32728
rect 38979 32725 38991 32759
rect 38933 32719 38991 32725
rect 40037 32759 40095 32765
rect 40037 32725 40049 32759
rect 40083 32756 40095 32759
rect 40126 32756 40132 32768
rect 40083 32728 40132 32756
rect 40083 32725 40095 32728
rect 40037 32719 40095 32725
rect 40126 32716 40132 32728
rect 40184 32716 40190 32768
rect 45554 32716 45560 32768
rect 45612 32756 45618 32768
rect 45649 32759 45707 32765
rect 45649 32756 45661 32759
rect 45612 32728 45661 32756
rect 45612 32716 45618 32728
rect 45649 32725 45661 32728
rect 45695 32725 45707 32759
rect 45649 32719 45707 32725
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 1765 32555 1823 32561
rect 1765 32521 1777 32555
rect 1811 32552 1823 32555
rect 5442 32552 5448 32564
rect 1811 32524 5448 32552
rect 1811 32521 1823 32524
rect 1765 32515 1823 32521
rect 5442 32512 5448 32524
rect 5500 32512 5506 32564
rect 5994 32512 6000 32564
rect 6052 32552 6058 32564
rect 6641 32555 6699 32561
rect 6641 32552 6653 32555
rect 6052 32524 6653 32552
rect 6052 32512 6058 32524
rect 6641 32521 6653 32524
rect 6687 32521 6699 32555
rect 10318 32552 10324 32564
rect 10279 32524 10324 32552
rect 6641 32515 6699 32521
rect 10318 32512 10324 32524
rect 10376 32512 10382 32564
rect 10781 32555 10839 32561
rect 10781 32521 10793 32555
rect 10827 32521 10839 32555
rect 10781 32515 10839 32521
rect 9208 32487 9266 32493
rect 9208 32453 9220 32487
rect 9254 32484 9266 32487
rect 10796 32484 10824 32515
rect 12066 32512 12072 32564
rect 12124 32552 12130 32564
rect 12253 32555 12311 32561
rect 12253 32552 12265 32555
rect 12124 32524 12265 32552
rect 12124 32512 12130 32524
rect 12253 32521 12265 32524
rect 12299 32521 12311 32555
rect 14550 32552 14556 32564
rect 14463 32524 14556 32552
rect 12253 32515 12311 32521
rect 14550 32512 14556 32524
rect 14608 32552 14614 32564
rect 15381 32555 15439 32561
rect 15381 32552 15393 32555
rect 14608 32524 15393 32552
rect 14608 32512 14614 32524
rect 15381 32521 15393 32524
rect 15427 32521 15439 32555
rect 15381 32515 15439 32521
rect 15473 32555 15531 32561
rect 15473 32521 15485 32555
rect 15519 32552 15531 32555
rect 17402 32552 17408 32564
rect 15519 32524 17408 32552
rect 15519 32521 15531 32524
rect 15473 32515 15531 32521
rect 17402 32512 17408 32524
rect 17460 32512 17466 32564
rect 18046 32552 18052 32564
rect 18007 32524 18052 32552
rect 18046 32512 18052 32524
rect 18104 32512 18110 32564
rect 24026 32512 24032 32564
rect 24084 32552 24090 32564
rect 24673 32555 24731 32561
rect 24673 32552 24685 32555
rect 24084 32524 24685 32552
rect 24084 32512 24090 32524
rect 24673 32521 24685 32524
rect 24719 32521 24731 32555
rect 24673 32515 24731 32521
rect 26234 32512 26240 32564
rect 26292 32552 26298 32564
rect 28537 32555 28595 32561
rect 26292 32524 26337 32552
rect 26292 32512 26298 32524
rect 28537 32521 28549 32555
rect 28583 32552 28595 32555
rect 28718 32552 28724 32564
rect 28583 32524 28724 32552
rect 28583 32521 28595 32524
rect 28537 32515 28595 32521
rect 28718 32512 28724 32524
rect 28776 32512 28782 32564
rect 33134 32552 33140 32564
rect 33095 32524 33140 32552
rect 33134 32512 33140 32524
rect 33192 32512 33198 32564
rect 33594 32552 33600 32564
rect 33555 32524 33600 32552
rect 33594 32512 33600 32524
rect 33652 32512 33658 32564
rect 34057 32555 34115 32561
rect 34057 32521 34069 32555
rect 34103 32552 34115 32555
rect 34606 32552 34612 32564
rect 34103 32524 34612 32552
rect 34103 32521 34115 32524
rect 34057 32515 34115 32521
rect 34606 32512 34612 32524
rect 34664 32512 34670 32564
rect 37918 32552 37924 32564
rect 35544 32524 37924 32552
rect 9254 32456 10824 32484
rect 13440 32487 13498 32493
rect 9254 32453 9266 32456
rect 9208 32447 9266 32453
rect 13440 32453 13452 32487
rect 13486 32484 13498 32487
rect 13538 32484 13544 32496
rect 13486 32456 13544 32484
rect 13486 32453 13498 32456
rect 13440 32447 13498 32453
rect 13538 32444 13544 32456
rect 13596 32444 13602 32496
rect 17420 32484 17448 32512
rect 20254 32484 20260 32496
rect 17420 32456 20260 32484
rect 20254 32444 20260 32456
rect 20312 32444 20318 32496
rect 23842 32484 23848 32496
rect 20732 32456 21588 32484
rect 1578 32416 1584 32428
rect 1539 32388 1584 32416
rect 1578 32376 1584 32388
rect 1636 32376 1642 32428
rect 3786 32416 3792 32428
rect 3747 32388 3792 32416
rect 3786 32376 3792 32388
rect 3844 32376 3850 32428
rect 6825 32419 6883 32425
rect 6825 32385 6837 32419
rect 6871 32416 6883 32419
rect 6914 32416 6920 32428
rect 6871 32388 6920 32416
rect 6871 32385 6883 32388
rect 6825 32379 6883 32385
rect 6914 32376 6920 32388
rect 6972 32376 6978 32428
rect 10965 32419 11023 32425
rect 10965 32385 10977 32419
rect 11011 32416 11023 32419
rect 11054 32416 11060 32428
rect 11011 32388 11060 32416
rect 11011 32385 11023 32388
rect 10965 32379 11023 32385
rect 11054 32376 11060 32388
rect 11112 32376 11118 32428
rect 13170 32416 13176 32428
rect 13131 32388 13176 32416
rect 13170 32376 13176 32388
rect 13228 32376 13234 32428
rect 17218 32376 17224 32428
rect 17276 32416 17282 32428
rect 17957 32419 18015 32425
rect 17957 32416 17969 32419
rect 17276 32388 17969 32416
rect 17276 32376 17282 32388
rect 17957 32385 17969 32388
rect 18003 32385 18015 32419
rect 18138 32416 18144 32428
rect 18099 32388 18144 32416
rect 17957 32379 18015 32385
rect 18138 32376 18144 32388
rect 18196 32376 18202 32428
rect 18969 32419 19027 32425
rect 18969 32385 18981 32419
rect 19015 32416 19027 32419
rect 19242 32416 19248 32428
rect 19015 32388 19248 32416
rect 19015 32385 19027 32388
rect 18969 32379 19027 32385
rect 19242 32376 19248 32388
rect 19300 32376 19306 32428
rect 20732 32425 20760 32456
rect 20717 32419 20775 32425
rect 20717 32416 20729 32419
rect 20456 32388 20729 32416
rect 3970 32348 3976 32360
rect 3931 32320 3976 32348
rect 3970 32308 3976 32320
rect 4028 32308 4034 32360
rect 4062 32308 4068 32360
rect 4120 32348 4126 32360
rect 4249 32351 4307 32357
rect 4249 32348 4261 32351
rect 4120 32320 4261 32348
rect 4120 32308 4126 32320
rect 4249 32317 4261 32320
rect 4295 32317 4307 32351
rect 8938 32348 8944 32360
rect 8899 32320 8944 32348
rect 4249 32311 4307 32317
rect 8938 32308 8944 32320
rect 8996 32308 9002 32360
rect 11793 32351 11851 32357
rect 11793 32317 11805 32351
rect 11839 32348 11851 32351
rect 11882 32348 11888 32360
rect 11839 32320 11888 32348
rect 11839 32317 11851 32320
rect 11793 32311 11851 32317
rect 11882 32308 11888 32320
rect 11940 32308 11946 32360
rect 15562 32308 15568 32360
rect 15620 32348 15626 32360
rect 17586 32348 17592 32360
rect 15620 32320 17592 32348
rect 15620 32308 15626 32320
rect 17586 32308 17592 32320
rect 17644 32308 17650 32360
rect 19061 32351 19119 32357
rect 19061 32317 19073 32351
rect 19107 32348 19119 32351
rect 19334 32348 19340 32360
rect 19107 32320 19340 32348
rect 19107 32317 19119 32320
rect 19061 32311 19119 32317
rect 19334 32308 19340 32320
rect 19392 32308 19398 32360
rect 12158 32280 12164 32292
rect 12119 32252 12164 32280
rect 12158 32240 12164 32252
rect 12216 32240 12222 32292
rect 20162 32280 20168 32292
rect 19352 32252 20168 32280
rect 15010 32212 15016 32224
rect 14971 32184 15016 32212
rect 15010 32172 15016 32184
rect 15068 32172 15074 32224
rect 19352 32221 19380 32252
rect 20162 32240 20168 32252
rect 20220 32280 20226 32292
rect 20456 32280 20484 32388
rect 20717 32385 20729 32388
rect 20763 32385 20775 32419
rect 21266 32416 21272 32428
rect 20717 32379 20775 32385
rect 21100 32388 21272 32416
rect 20625 32351 20683 32357
rect 20625 32317 20637 32351
rect 20671 32348 20683 32351
rect 21100 32348 21128 32388
rect 21266 32376 21272 32388
rect 21324 32416 21330 32428
rect 21453 32419 21511 32425
rect 21453 32416 21465 32419
rect 21324 32388 21465 32416
rect 21324 32376 21330 32388
rect 21453 32385 21465 32388
rect 21499 32385 21511 32419
rect 21453 32379 21511 32385
rect 20671 32320 21128 32348
rect 21177 32351 21235 32357
rect 20671 32317 20683 32320
rect 20625 32311 20683 32317
rect 21177 32317 21189 32351
rect 21223 32348 21235 32351
rect 21560 32348 21588 32456
rect 22020 32456 23848 32484
rect 22020 32360 22048 32456
rect 23842 32444 23848 32456
rect 23900 32484 23906 32496
rect 28350 32484 28356 32496
rect 23900 32456 28356 32484
rect 23900 32444 23906 32456
rect 22094 32376 22100 32428
rect 22152 32416 22158 32428
rect 22261 32419 22319 32425
rect 22261 32416 22273 32419
rect 22152 32388 22273 32416
rect 22152 32376 22158 32388
rect 22261 32385 22273 32388
rect 22307 32385 22319 32419
rect 22261 32379 22319 32385
rect 24765 32419 24823 32425
rect 24765 32385 24777 32419
rect 24811 32385 24823 32419
rect 25038 32416 25044 32428
rect 24999 32388 25044 32416
rect 24765 32379 24823 32385
rect 22002 32348 22008 32360
rect 21223 32320 21588 32348
rect 21963 32320 22008 32348
rect 21223 32317 21235 32320
rect 21177 32311 21235 32317
rect 22002 32308 22008 32320
rect 22060 32308 22066 32360
rect 24780 32348 24808 32379
rect 25038 32376 25044 32388
rect 25096 32376 25102 32428
rect 26142 32416 26148 32428
rect 26103 32388 26148 32416
rect 26142 32376 26148 32388
rect 26200 32376 26206 32428
rect 26421 32419 26479 32425
rect 26421 32385 26433 32419
rect 26467 32416 26479 32419
rect 26510 32416 26516 32428
rect 26467 32388 26516 32416
rect 26467 32385 26479 32388
rect 26421 32379 26479 32385
rect 26510 32376 26516 32388
rect 26568 32376 26574 32428
rect 27172 32425 27200 32456
rect 28350 32444 28356 32456
rect 28408 32444 28414 32496
rect 31018 32444 31024 32496
rect 31076 32484 31082 32496
rect 31076 32456 32720 32484
rect 31076 32444 31082 32456
rect 27157 32419 27215 32425
rect 27157 32385 27169 32419
rect 27203 32385 27215 32419
rect 27413 32419 27471 32425
rect 27413 32416 27425 32419
rect 27157 32379 27215 32385
rect 27264 32388 27425 32416
rect 25866 32348 25872 32360
rect 24780 32320 25872 32348
rect 25866 32308 25872 32320
rect 25924 32308 25930 32360
rect 26605 32351 26663 32357
rect 26605 32317 26617 32351
rect 26651 32348 26663 32351
rect 27264 32348 27292 32388
rect 27413 32385 27425 32388
rect 27459 32385 27471 32419
rect 31386 32416 31392 32428
rect 31347 32388 31392 32416
rect 27413 32379 27471 32385
rect 31386 32376 31392 32388
rect 31444 32376 31450 32428
rect 31662 32376 31668 32428
rect 31720 32416 31726 32428
rect 32692 32425 32720 32456
rect 32858 32444 32864 32496
rect 32916 32484 32922 32496
rect 33965 32487 34023 32493
rect 33965 32484 33977 32487
rect 32916 32456 33977 32484
rect 32916 32444 32922 32456
rect 33965 32453 33977 32456
rect 34011 32453 34023 32487
rect 33965 32447 34023 32453
rect 32493 32419 32551 32425
rect 32493 32416 32505 32419
rect 31720 32388 32505 32416
rect 31720 32376 31726 32388
rect 32493 32385 32505 32388
rect 32539 32385 32551 32419
rect 32493 32379 32551 32385
rect 32677 32419 32735 32425
rect 32677 32385 32689 32419
rect 32723 32385 32735 32419
rect 33042 32416 33048 32428
rect 33003 32388 33048 32416
rect 32677 32379 32735 32385
rect 33042 32376 33048 32388
rect 33100 32376 33106 32428
rect 34790 32376 34796 32428
rect 34848 32416 34854 32428
rect 35161 32419 35219 32425
rect 35161 32416 35173 32419
rect 34848 32388 35173 32416
rect 34848 32376 34854 32388
rect 35161 32385 35173 32388
rect 35207 32385 35219 32419
rect 35161 32379 35219 32385
rect 35250 32376 35256 32428
rect 35308 32416 35314 32428
rect 35544 32425 35572 32524
rect 37918 32512 37924 32524
rect 37976 32512 37982 32564
rect 40218 32512 40224 32564
rect 40276 32552 40282 32564
rect 40497 32555 40555 32561
rect 40497 32552 40509 32555
rect 40276 32524 40509 32552
rect 40276 32512 40282 32524
rect 40497 32521 40509 32524
rect 40543 32521 40555 32555
rect 47762 32552 47768 32564
rect 40497 32515 40555 32521
rect 40604 32524 47768 32552
rect 36354 32484 36360 32496
rect 36315 32456 36360 32484
rect 36354 32444 36360 32456
rect 36412 32444 36418 32496
rect 40604 32484 40632 32524
rect 47762 32512 47768 32524
rect 47820 32512 47826 32564
rect 39868 32456 40632 32484
rect 39868 32428 39896 32456
rect 45554 32444 45560 32496
rect 45612 32484 45618 32496
rect 45612 32456 45657 32484
rect 45612 32444 45618 32456
rect 46474 32444 46480 32496
rect 46532 32484 46538 32496
rect 47213 32487 47271 32493
rect 46532 32456 47164 32484
rect 46532 32444 46538 32456
rect 35529 32419 35587 32425
rect 35529 32416 35541 32419
rect 35308 32388 35541 32416
rect 35308 32376 35314 32388
rect 35529 32385 35541 32388
rect 35575 32385 35587 32419
rect 35529 32379 35587 32385
rect 35713 32419 35771 32425
rect 35713 32385 35725 32419
rect 35759 32416 35771 32419
rect 35986 32416 35992 32428
rect 35759 32388 35992 32416
rect 35759 32385 35771 32388
rect 35713 32379 35771 32385
rect 35986 32376 35992 32388
rect 36044 32376 36050 32428
rect 36170 32376 36176 32428
rect 36228 32416 36234 32428
rect 36541 32419 36599 32425
rect 36541 32416 36553 32419
rect 36228 32388 36553 32416
rect 36228 32376 36234 32388
rect 36541 32385 36553 32388
rect 36587 32385 36599 32419
rect 38010 32416 38016 32428
rect 37971 32388 38016 32416
rect 36541 32379 36599 32385
rect 38010 32376 38016 32388
rect 38068 32376 38074 32428
rect 38286 32425 38292 32428
rect 38280 32379 38292 32425
rect 38344 32416 38350 32428
rect 39850 32416 39856 32428
rect 38344 32388 38380 32416
rect 39811 32388 39856 32416
rect 38286 32376 38292 32379
rect 38344 32376 38350 32388
rect 39850 32376 39856 32388
rect 39908 32376 39914 32428
rect 40034 32416 40040 32428
rect 39995 32388 40040 32416
rect 40034 32376 40040 32388
rect 40092 32376 40098 32428
rect 40310 32416 40316 32428
rect 40271 32388 40316 32416
rect 40310 32376 40316 32388
rect 40368 32376 40374 32428
rect 44634 32376 44640 32428
rect 44692 32416 44698 32428
rect 44729 32419 44787 32425
rect 44729 32416 44741 32419
rect 44692 32388 44741 32416
rect 44692 32376 44698 32388
rect 44729 32385 44741 32388
rect 44775 32385 44787 32419
rect 47136 32416 47164 32456
rect 47213 32453 47225 32487
rect 47259 32484 47271 32487
rect 47302 32484 47308 32496
rect 47259 32456 47308 32484
rect 47259 32453 47271 32456
rect 47213 32447 47271 32453
rect 47302 32444 47308 32456
rect 47360 32444 47366 32496
rect 47765 32419 47823 32425
rect 47765 32416 47777 32419
rect 47136 32388 47777 32416
rect 44729 32379 44787 32385
rect 47765 32385 47777 32388
rect 47811 32385 47823 32419
rect 47765 32379 47823 32385
rect 26651 32320 27292 32348
rect 31481 32351 31539 32357
rect 26651 32317 26663 32320
rect 26605 32311 26663 32317
rect 31481 32317 31493 32351
rect 31527 32348 31539 32351
rect 31570 32348 31576 32360
rect 31527 32320 31576 32348
rect 31527 32317 31539 32320
rect 31481 32311 31539 32317
rect 31570 32308 31576 32320
rect 31628 32308 31634 32360
rect 31754 32308 31760 32360
rect 31812 32348 31818 32360
rect 32309 32351 32367 32357
rect 32309 32348 32321 32351
rect 31812 32320 32321 32348
rect 31812 32308 31818 32320
rect 32309 32317 32321 32320
rect 32355 32317 32367 32351
rect 32309 32311 32367 32317
rect 34241 32351 34299 32357
rect 34241 32317 34253 32351
rect 34287 32317 34299 32351
rect 34241 32311 34299 32317
rect 21361 32283 21419 32289
rect 21361 32280 21373 32283
rect 20220 32252 20484 32280
rect 20548 32252 21373 32280
rect 20220 32240 20226 32252
rect 19337 32215 19395 32221
rect 19337 32181 19349 32215
rect 19383 32181 19395 32215
rect 19337 32175 19395 32181
rect 19978 32172 19984 32224
rect 20036 32212 20042 32224
rect 20349 32215 20407 32221
rect 20349 32212 20361 32215
rect 20036 32184 20361 32212
rect 20036 32172 20042 32184
rect 20349 32181 20361 32184
rect 20395 32181 20407 32215
rect 20349 32175 20407 32181
rect 20438 32172 20444 32224
rect 20496 32212 20502 32224
rect 20548 32221 20576 32252
rect 21361 32249 21373 32252
rect 21407 32249 21419 32283
rect 21361 32243 21419 32249
rect 31021 32283 31079 32289
rect 31021 32249 31033 32283
rect 31067 32280 31079 32283
rect 31772 32280 31800 32308
rect 31067 32252 31800 32280
rect 34256 32280 34284 32311
rect 34698 32308 34704 32360
rect 34756 32348 34762 32360
rect 35345 32351 35403 32357
rect 35345 32348 35357 32351
rect 34756 32320 35357 32348
rect 34756 32308 34762 32320
rect 35345 32317 35357 32320
rect 35391 32317 35403 32351
rect 35345 32311 35403 32317
rect 35437 32351 35495 32357
rect 35437 32317 35449 32351
rect 35483 32348 35495 32351
rect 35618 32348 35624 32360
rect 35483 32320 35624 32348
rect 35483 32317 35495 32320
rect 35437 32311 35495 32317
rect 35618 32308 35624 32320
rect 35676 32308 35682 32360
rect 45370 32348 45376 32360
rect 45331 32320 45376 32348
rect 45370 32308 45376 32320
rect 45428 32308 45434 32360
rect 36906 32280 36912 32292
rect 34256 32252 36912 32280
rect 31067 32249 31079 32252
rect 31021 32243 31079 32249
rect 36906 32240 36912 32252
rect 36964 32240 36970 32292
rect 20533 32215 20591 32221
rect 20533 32212 20545 32215
rect 20496 32184 20545 32212
rect 20496 32172 20502 32184
rect 20533 32181 20545 32184
rect 20579 32181 20591 32215
rect 21266 32212 21272 32224
rect 21227 32184 21272 32212
rect 20533 32175 20591 32181
rect 21266 32172 21272 32184
rect 21324 32172 21330 32224
rect 23382 32212 23388 32224
rect 23343 32184 23388 32212
rect 23382 32172 23388 32184
rect 23440 32172 23446 32224
rect 34977 32215 35035 32221
rect 34977 32181 34989 32215
rect 35023 32212 35035 32215
rect 35434 32212 35440 32224
rect 35023 32184 35440 32212
rect 35023 32181 35035 32184
rect 34977 32175 35035 32181
rect 35434 32172 35440 32184
rect 35492 32172 35498 32224
rect 36170 32212 36176 32224
rect 36131 32184 36176 32212
rect 36170 32172 36176 32184
rect 36228 32172 36234 32224
rect 39390 32212 39396 32224
rect 39351 32184 39396 32212
rect 39390 32172 39396 32184
rect 39448 32172 39454 32224
rect 44821 32215 44879 32221
rect 44821 32181 44833 32215
rect 44867 32212 44879 32215
rect 46014 32212 46020 32224
rect 44867 32184 46020 32212
rect 44867 32181 44879 32184
rect 44821 32175 44879 32181
rect 46014 32172 46020 32184
rect 46072 32172 46078 32224
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 3970 31968 3976 32020
rect 4028 32008 4034 32020
rect 4525 32011 4583 32017
rect 4525 32008 4537 32011
rect 4028 31980 4537 32008
rect 4028 31968 4034 31980
rect 4525 31977 4537 31980
rect 4571 31977 4583 32011
rect 4525 31971 4583 31977
rect 8938 31968 8944 32020
rect 8996 32008 9002 32020
rect 9217 32011 9275 32017
rect 9217 32008 9229 32011
rect 8996 31980 9229 32008
rect 8996 31968 9002 31980
rect 9217 31977 9229 31980
rect 9263 31977 9275 32011
rect 11054 32008 11060 32020
rect 11015 31980 11060 32008
rect 9217 31971 9275 31977
rect 11054 31968 11060 31980
rect 11112 31968 11118 32020
rect 14274 32008 14280 32020
rect 14235 31980 14280 32008
rect 14274 31968 14280 31980
rect 14332 31968 14338 32020
rect 15378 32008 15384 32020
rect 15212 31980 15384 32008
rect 6181 31943 6239 31949
rect 6181 31909 6193 31943
rect 6227 31940 6239 31943
rect 9398 31940 9404 31952
rect 6227 31912 9404 31940
rect 6227 31909 6239 31912
rect 6181 31903 6239 31909
rect 9398 31900 9404 31912
rect 9456 31940 9462 31952
rect 14461 31943 14519 31949
rect 9456 31912 10456 31940
rect 9456 31900 9462 31912
rect 6730 31872 6736 31884
rect 4632 31844 6736 31872
rect 4632 31813 4660 31844
rect 6730 31832 6736 31844
rect 6788 31832 6794 31884
rect 7006 31872 7012 31884
rect 6967 31844 7012 31872
rect 7006 31832 7012 31844
rect 7064 31832 7070 31884
rect 10428 31881 10456 31912
rect 14461 31909 14473 31943
rect 14507 31940 14519 31943
rect 15010 31940 15016 31952
rect 14507 31912 15016 31940
rect 14507 31909 14519 31912
rect 14461 31903 14519 31909
rect 15010 31900 15016 31912
rect 15068 31900 15074 31952
rect 15212 31881 15240 31980
rect 15378 31968 15384 31980
rect 15436 31968 15442 32020
rect 19334 31968 19340 32020
rect 19392 32008 19398 32020
rect 19429 32011 19487 32017
rect 19429 32008 19441 32011
rect 19392 31980 19441 32008
rect 19392 31968 19398 31980
rect 19429 31977 19441 31980
rect 19475 31977 19487 32011
rect 19429 31971 19487 31977
rect 20438 31968 20444 32020
rect 20496 32008 20502 32020
rect 21913 32011 21971 32017
rect 20496 31980 21220 32008
rect 20496 31968 20502 31980
rect 21192 31940 21220 31980
rect 21913 31977 21925 32011
rect 21959 32008 21971 32011
rect 22094 32008 22100 32020
rect 21959 31980 22100 32008
rect 21959 31977 21971 31980
rect 21913 31971 21971 31977
rect 22094 31968 22100 31980
rect 22152 31968 22158 32020
rect 31018 31968 31024 32020
rect 31076 32008 31082 32020
rect 31076 31980 31984 32008
rect 31076 31968 31082 31980
rect 23845 31943 23903 31949
rect 23845 31940 23857 31943
rect 21192 31912 22140 31940
rect 10413 31875 10471 31881
rect 10413 31841 10425 31875
rect 10459 31841 10471 31875
rect 10413 31835 10471 31841
rect 15197 31875 15255 31881
rect 15197 31841 15209 31875
rect 15243 31841 15255 31875
rect 17586 31872 17592 31884
rect 17547 31844 17592 31872
rect 15197 31835 15255 31841
rect 17586 31832 17592 31844
rect 17644 31832 17650 31884
rect 20809 31875 20867 31881
rect 20809 31841 20821 31875
rect 20855 31872 20867 31875
rect 22002 31872 22008 31884
rect 20855 31844 22008 31872
rect 20855 31841 20867 31844
rect 20809 31835 20867 31841
rect 22002 31832 22008 31844
rect 22060 31832 22066 31884
rect 22112 31881 22140 31912
rect 22480 31912 23857 31940
rect 22480 31884 22508 31912
rect 23845 31909 23857 31912
rect 23891 31909 23903 31943
rect 23845 31903 23903 31909
rect 31113 31943 31171 31949
rect 31113 31909 31125 31943
rect 31159 31940 31171 31943
rect 31294 31940 31300 31952
rect 31159 31912 31300 31940
rect 31159 31909 31171 31912
rect 31113 31903 31171 31909
rect 31294 31900 31300 31912
rect 31352 31900 31358 31952
rect 22097 31875 22155 31881
rect 22097 31841 22109 31875
rect 22143 31841 22155 31875
rect 22462 31872 22468 31884
rect 22423 31844 22468 31872
rect 22097 31835 22155 31841
rect 22462 31832 22468 31844
rect 22520 31832 22526 31884
rect 22557 31875 22615 31881
rect 22557 31841 22569 31875
rect 22603 31872 22615 31875
rect 23382 31872 23388 31884
rect 22603 31844 23388 31872
rect 22603 31841 22615 31844
rect 22557 31835 22615 31841
rect 23382 31832 23388 31844
rect 23440 31832 23446 31884
rect 31754 31872 31760 31884
rect 31128 31844 31760 31872
rect 4617 31807 4675 31813
rect 4617 31773 4629 31807
rect 4663 31773 4675 31807
rect 4617 31767 4675 31773
rect 5442 31764 5448 31816
rect 5500 31804 5506 31816
rect 5905 31807 5963 31813
rect 5905 31804 5917 31807
rect 5500 31776 5917 31804
rect 5500 31764 5506 31776
rect 5905 31773 5917 31776
rect 5951 31773 5963 31807
rect 7098 31804 7104 31816
rect 7059 31776 7104 31804
rect 5905 31767 5963 31773
rect 7098 31764 7104 31776
rect 7156 31764 7162 31816
rect 9214 31804 9220 31816
rect 9175 31776 9220 31804
rect 9214 31764 9220 31776
rect 9272 31764 9278 31816
rect 10594 31804 10600 31816
rect 10555 31776 10600 31804
rect 10594 31764 10600 31776
rect 10652 31764 10658 31816
rect 11882 31764 11888 31816
rect 11940 31804 11946 31816
rect 14737 31807 14795 31813
rect 14737 31804 14749 31807
rect 11940 31776 14749 31804
rect 11940 31764 11946 31776
rect 14737 31773 14749 31776
rect 14783 31804 14795 31807
rect 15286 31804 15292 31816
rect 14783 31776 15292 31804
rect 14783 31773 14795 31776
rect 14737 31767 14795 31773
rect 15286 31764 15292 31776
rect 15344 31764 15350 31816
rect 17512 31776 22140 31804
rect 10689 31739 10747 31745
rect 10689 31705 10701 31739
rect 10735 31736 10747 31739
rect 14550 31736 14556 31748
rect 10735 31708 14556 31736
rect 10735 31705 10747 31708
rect 10689 31699 10747 31705
rect 14550 31696 14556 31708
rect 14608 31696 14614 31748
rect 15464 31739 15522 31745
rect 15464 31705 15476 31739
rect 15510 31736 15522 31739
rect 15654 31736 15660 31748
rect 15510 31708 15660 31736
rect 15510 31705 15522 31708
rect 15464 31699 15522 31705
rect 15654 31696 15660 31708
rect 15712 31696 15718 31748
rect 17512 31745 17540 31776
rect 17405 31739 17463 31745
rect 17405 31736 17417 31739
rect 16592 31708 17417 31736
rect 16592 31680 16620 31708
rect 17405 31705 17417 31708
rect 17451 31705 17463 31739
rect 17405 31699 17463 31705
rect 17497 31739 17555 31745
rect 17497 31705 17509 31739
rect 17543 31705 17555 31739
rect 17497 31699 17555 31705
rect 20162 31696 20168 31748
rect 20220 31736 20226 31748
rect 20542 31739 20600 31745
rect 20542 31736 20554 31739
rect 20220 31708 20554 31736
rect 20220 31696 20226 31708
rect 20542 31705 20554 31708
rect 20588 31705 20600 31739
rect 22112 31736 22140 31776
rect 22186 31764 22192 31816
rect 22244 31804 22250 31816
rect 23661 31807 23719 31813
rect 22244 31776 22289 31804
rect 22244 31764 22250 31776
rect 23661 31773 23673 31807
rect 23707 31804 23719 31807
rect 23934 31804 23940 31816
rect 23707 31776 23940 31804
rect 23707 31773 23719 31776
rect 23661 31767 23719 31773
rect 23934 31764 23940 31776
rect 23992 31804 23998 31816
rect 24765 31807 24823 31813
rect 24765 31804 24777 31807
rect 23992 31776 24777 31804
rect 23992 31764 23998 31776
rect 24765 31773 24777 31776
rect 24811 31773 24823 31807
rect 25038 31804 25044 31816
rect 24999 31776 25044 31804
rect 24765 31767 24823 31773
rect 25038 31764 25044 31776
rect 25096 31804 25102 31816
rect 25593 31807 25651 31813
rect 25593 31804 25605 31807
rect 25096 31776 25605 31804
rect 25096 31764 25102 31776
rect 25593 31773 25605 31776
rect 25639 31804 25651 31807
rect 25774 31804 25780 31816
rect 25639 31776 25780 31804
rect 25639 31773 25651 31776
rect 25593 31767 25651 31773
rect 25774 31764 25780 31776
rect 25832 31764 25838 31816
rect 30837 31807 30895 31813
rect 30837 31804 30849 31807
rect 30760 31776 30849 31804
rect 22370 31736 22376 31748
rect 22112 31708 22376 31736
rect 20542 31699 20600 31705
rect 22370 31696 22376 31708
rect 22428 31696 22434 31748
rect 24136 31708 25912 31736
rect 6546 31628 6552 31680
rect 6604 31668 6610 31680
rect 6733 31671 6791 31677
rect 6733 31668 6745 31671
rect 6604 31640 6745 31668
rect 6604 31628 6610 31640
rect 6733 31637 6745 31640
rect 6779 31637 6791 31671
rect 6733 31631 6791 31637
rect 16574 31628 16580 31680
rect 16632 31668 16638 31680
rect 17034 31668 17040 31680
rect 16632 31640 16725 31668
rect 16995 31640 17040 31668
rect 16632 31628 16638 31640
rect 17034 31628 17040 31640
rect 17092 31628 17098 31680
rect 17954 31628 17960 31680
rect 18012 31668 18018 31680
rect 24136 31668 24164 31708
rect 25884 31680 25912 31708
rect 29730 31696 29736 31748
rect 29788 31736 29794 31748
rect 30760 31736 30788 31776
rect 30837 31773 30849 31776
rect 30883 31773 30895 31807
rect 30837 31767 30895 31773
rect 30929 31807 30987 31813
rect 30929 31773 30941 31807
rect 30975 31804 30987 31807
rect 31018 31804 31024 31816
rect 30975 31776 31024 31804
rect 30975 31773 30987 31776
rect 30929 31767 30987 31773
rect 31018 31764 31024 31776
rect 31076 31764 31082 31816
rect 31128 31813 31156 31844
rect 31754 31832 31760 31844
rect 31812 31832 31818 31884
rect 31956 31881 31984 31980
rect 35618 31968 35624 32020
rect 35676 32008 35682 32020
rect 36725 32011 36783 32017
rect 36725 32008 36737 32011
rect 35676 31980 36737 32008
rect 35676 31968 35682 31980
rect 36725 31977 36737 31980
rect 36771 31977 36783 32011
rect 38286 32008 38292 32020
rect 38247 31980 38292 32008
rect 36725 31971 36783 31977
rect 38286 31968 38292 31980
rect 38344 31968 38350 32020
rect 38933 32011 38991 32017
rect 38933 31977 38945 32011
rect 38979 32008 38991 32011
rect 39114 32008 39120 32020
rect 38979 31980 39120 32008
rect 38979 31977 38991 31980
rect 38933 31971 38991 31977
rect 39114 31968 39120 31980
rect 39172 31968 39178 32020
rect 41322 31968 41328 32020
rect 41380 32008 41386 32020
rect 41417 32011 41475 32017
rect 41417 32008 41429 32011
rect 41380 31980 41429 32008
rect 41380 31968 41386 31980
rect 41417 31977 41429 31980
rect 41463 31977 41475 32011
rect 41417 31971 41475 31977
rect 31941 31875 31999 31881
rect 31941 31841 31953 31875
rect 31987 31841 31999 31875
rect 35342 31872 35348 31884
rect 35303 31844 35348 31872
rect 31941 31835 31999 31841
rect 35342 31832 35348 31844
rect 35400 31832 35406 31884
rect 37918 31872 37924 31884
rect 37879 31844 37924 31872
rect 37918 31832 37924 31844
rect 37976 31832 37982 31884
rect 38010 31832 38016 31884
rect 38068 31872 38074 31884
rect 40034 31872 40040 31884
rect 38068 31844 40040 31872
rect 38068 31832 38074 31844
rect 40034 31832 40040 31844
rect 40092 31832 40098 31884
rect 46014 31872 46020 31884
rect 45975 31844 46020 31872
rect 46014 31832 46020 31844
rect 46072 31832 46078 31884
rect 47673 31875 47731 31881
rect 47673 31841 47685 31875
rect 47719 31872 47731 31875
rect 47946 31872 47952 31884
rect 47719 31844 47952 31872
rect 47719 31841 47731 31844
rect 47673 31835 47731 31841
rect 47946 31832 47952 31844
rect 48004 31832 48010 31884
rect 31113 31807 31171 31813
rect 31113 31773 31125 31807
rect 31159 31773 31171 31807
rect 31113 31767 31171 31773
rect 31662 31764 31668 31816
rect 31720 31804 31726 31816
rect 31849 31807 31907 31813
rect 31849 31804 31861 31807
rect 31720 31776 31861 31804
rect 31720 31764 31726 31776
rect 31849 31773 31861 31776
rect 31895 31773 31907 31807
rect 31849 31767 31907 31773
rect 32033 31807 32091 31813
rect 32033 31773 32045 31807
rect 32079 31804 32091 31807
rect 32079 31776 34928 31804
rect 32079 31773 32091 31776
rect 32033 31767 32091 31773
rect 31680 31736 31708 31764
rect 29788 31708 31708 31736
rect 34900 31736 34928 31776
rect 35434 31764 35440 31816
rect 35492 31804 35498 31816
rect 35601 31807 35659 31813
rect 35601 31804 35613 31807
rect 35492 31776 35613 31804
rect 35492 31764 35498 31776
rect 35601 31773 35613 31776
rect 35647 31773 35659 31807
rect 37550 31804 37556 31816
rect 37511 31776 37556 31804
rect 35601 31767 35659 31773
rect 37550 31764 37556 31776
rect 37608 31764 37614 31816
rect 37642 31764 37648 31816
rect 37700 31804 37706 31816
rect 37737 31807 37795 31813
rect 37737 31804 37749 31807
rect 37700 31776 37749 31804
rect 37700 31764 37706 31776
rect 37737 31773 37749 31776
rect 37783 31773 37795 31807
rect 37737 31767 37795 31773
rect 37829 31807 37887 31813
rect 37829 31773 37841 31807
rect 37875 31773 37887 31807
rect 37829 31767 37887 31773
rect 35802 31736 35808 31748
rect 34900 31708 35808 31736
rect 29788 31696 29794 31708
rect 35802 31696 35808 31708
rect 35860 31696 35866 31748
rect 18012 31640 24164 31668
rect 18012 31628 18018 31640
rect 25130 31628 25136 31680
rect 25188 31668 25194 31680
rect 25682 31668 25688 31680
rect 25188 31640 25688 31668
rect 25188 31628 25194 31640
rect 25682 31628 25688 31640
rect 25740 31628 25746 31680
rect 25866 31628 25872 31680
rect 25924 31628 25930 31680
rect 31570 31668 31576 31680
rect 31531 31640 31576 31668
rect 31570 31628 31576 31640
rect 31628 31628 31634 31680
rect 34698 31628 34704 31680
rect 34756 31668 34762 31680
rect 36078 31668 36084 31680
rect 34756 31640 36084 31668
rect 34756 31628 34762 31640
rect 36078 31628 36084 31640
rect 36136 31628 36142 31680
rect 37844 31668 37872 31767
rect 37936 31736 37964 31832
rect 38105 31807 38163 31813
rect 38105 31773 38117 31807
rect 38151 31804 38163 31807
rect 39301 31807 39359 31813
rect 39301 31804 39313 31807
rect 38151 31776 39313 31804
rect 38151 31773 38163 31776
rect 38105 31767 38163 31773
rect 39301 31773 39313 31776
rect 39347 31804 39359 31807
rect 39390 31804 39396 31816
rect 39347 31776 39396 31804
rect 39347 31773 39359 31776
rect 39301 31767 39359 31773
rect 39390 31764 39396 31776
rect 39448 31764 39454 31816
rect 40126 31764 40132 31816
rect 40184 31804 40190 31816
rect 40293 31807 40351 31813
rect 40293 31804 40305 31807
rect 40184 31776 40305 31804
rect 40184 31764 40190 31776
rect 40293 31773 40305 31776
rect 40339 31773 40351 31807
rect 45830 31804 45836 31816
rect 45791 31776 45836 31804
rect 40293 31767 40351 31773
rect 45830 31764 45836 31776
rect 45888 31764 45894 31816
rect 38010 31736 38016 31748
rect 37936 31708 38016 31736
rect 38010 31696 38016 31708
rect 38068 31696 38074 31748
rect 39117 31739 39175 31745
rect 39117 31705 39129 31739
rect 39163 31736 39175 31739
rect 39206 31736 39212 31748
rect 39163 31708 39212 31736
rect 39163 31705 39175 31708
rect 39117 31699 39175 31705
rect 39206 31696 39212 31708
rect 39264 31696 39270 31748
rect 37918 31668 37924 31680
rect 37844 31640 37924 31668
rect 37918 31628 37924 31640
rect 37976 31628 37982 31680
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 13081 31467 13139 31473
rect 13081 31433 13093 31467
rect 13127 31433 13139 31467
rect 13081 31427 13139 31433
rect 13449 31467 13507 31473
rect 13449 31433 13461 31467
rect 13495 31464 13507 31467
rect 16574 31464 16580 31476
rect 13495 31436 16580 31464
rect 13495 31433 13507 31436
rect 13449 31427 13507 31433
rect 5905 31399 5963 31405
rect 5905 31365 5917 31399
rect 5951 31396 5963 31399
rect 6733 31399 6791 31405
rect 6733 31396 6745 31399
rect 5951 31368 6745 31396
rect 5951 31365 5963 31368
rect 5905 31359 5963 31365
rect 6733 31365 6745 31368
rect 6779 31365 6791 31399
rect 6733 31359 6791 31365
rect 6914 31356 6920 31408
rect 6972 31396 6978 31408
rect 8018 31396 8024 31408
rect 6972 31368 8024 31396
rect 6972 31356 6978 31368
rect 8018 31356 8024 31368
rect 8076 31396 8082 31408
rect 9214 31396 9220 31408
rect 8076 31368 9220 31396
rect 8076 31356 8082 31368
rect 5997 31331 6055 31337
rect 5997 31297 6009 31331
rect 6043 31297 6055 31331
rect 6546 31328 6552 31340
rect 6507 31300 6552 31328
rect 5997 31291 6055 31297
rect 6012 31260 6040 31291
rect 6546 31288 6552 31300
rect 6604 31288 6610 31340
rect 9048 31337 9076 31368
rect 9214 31356 9220 31368
rect 9272 31356 9278 31408
rect 9033 31331 9091 31337
rect 9033 31297 9045 31331
rect 9079 31297 9091 31331
rect 9033 31291 9091 31297
rect 10505 31331 10563 31337
rect 10505 31297 10517 31331
rect 10551 31328 10563 31331
rect 11698 31328 11704 31340
rect 10551 31300 11704 31328
rect 10551 31297 10563 31300
rect 10505 31291 10563 31297
rect 11698 31288 11704 31300
rect 11756 31288 11762 31340
rect 12621 31331 12679 31337
rect 12621 31297 12633 31331
rect 12667 31328 12679 31331
rect 13096 31328 13124 31427
rect 16574 31424 16580 31436
rect 16632 31424 16638 31476
rect 20162 31464 20168 31476
rect 20123 31436 20168 31464
rect 20162 31424 20168 31436
rect 20220 31424 20226 31476
rect 24857 31467 24915 31473
rect 24857 31433 24869 31467
rect 24903 31464 24915 31467
rect 24946 31464 24952 31476
rect 24903 31436 24952 31464
rect 24903 31433 24915 31436
rect 24857 31427 24915 31433
rect 24946 31424 24952 31436
rect 25004 31424 25010 31476
rect 25774 31464 25780 31476
rect 25735 31436 25780 31464
rect 25774 31424 25780 31436
rect 25832 31424 25838 31476
rect 34790 31424 34796 31476
rect 34848 31464 34854 31476
rect 35069 31467 35127 31473
rect 35069 31464 35081 31467
rect 34848 31436 35081 31464
rect 34848 31424 34854 31436
rect 35069 31433 35081 31436
rect 35115 31433 35127 31467
rect 35986 31464 35992 31476
rect 35947 31436 35992 31464
rect 35069 31427 35127 31433
rect 35986 31424 35992 31436
rect 36044 31424 36050 31476
rect 44269 31467 44327 31473
rect 44269 31433 44281 31467
rect 44315 31464 44327 31467
rect 44450 31464 44456 31476
rect 44315 31436 44456 31464
rect 44315 31433 44327 31436
rect 44269 31427 44327 31433
rect 44450 31424 44456 31436
rect 44508 31464 44514 31476
rect 45370 31464 45376 31476
rect 44508 31436 45376 31464
rect 44508 31424 44514 31436
rect 45370 31424 45376 31436
rect 45428 31424 45434 31476
rect 15286 31356 15292 31408
rect 15344 31396 15350 31408
rect 15473 31399 15531 31405
rect 15473 31396 15485 31399
rect 15344 31368 15485 31396
rect 15344 31356 15350 31368
rect 15473 31365 15485 31368
rect 15519 31396 15531 31399
rect 16945 31399 17003 31405
rect 16945 31396 16957 31399
rect 15519 31368 16957 31396
rect 15519 31365 15531 31368
rect 15473 31359 15531 31365
rect 16945 31365 16957 31368
rect 16991 31365 17003 31399
rect 16945 31359 17003 31365
rect 19889 31399 19947 31405
rect 19889 31365 19901 31399
rect 19935 31396 19947 31399
rect 21266 31396 21272 31408
rect 19935 31368 21272 31396
rect 19935 31365 19947 31368
rect 19889 31359 19947 31365
rect 21266 31356 21272 31368
rect 21324 31356 21330 31408
rect 31018 31396 31024 31408
rect 30208 31368 31024 31396
rect 12667 31300 13124 31328
rect 12667 31297 12679 31300
rect 12621 31291 12679 31297
rect 16482 31288 16488 31340
rect 16540 31328 16546 31340
rect 17954 31328 17960 31340
rect 16540 31300 17960 31328
rect 16540 31288 16546 31300
rect 17954 31288 17960 31300
rect 18012 31288 18018 31340
rect 18049 31331 18107 31337
rect 18049 31297 18061 31331
rect 18095 31297 18107 31331
rect 18049 31291 18107 31297
rect 6086 31260 6092 31272
rect 5999 31232 6092 31260
rect 6086 31220 6092 31232
rect 6144 31260 6150 31272
rect 6454 31260 6460 31272
rect 6144 31232 6460 31260
rect 6144 31220 6150 31232
rect 6454 31220 6460 31232
rect 6512 31220 6518 31272
rect 8202 31260 8208 31272
rect 8163 31232 8208 31260
rect 8202 31220 8208 31232
rect 8260 31220 8266 31272
rect 13538 31260 13544 31272
rect 13499 31232 13544 31260
rect 13538 31220 13544 31232
rect 13596 31220 13602 31272
rect 13633 31263 13691 31269
rect 13633 31229 13645 31263
rect 13679 31229 13691 31263
rect 13633 31223 13691 31229
rect 17405 31263 17463 31269
rect 17405 31229 17417 31263
rect 17451 31260 17463 31263
rect 18064 31260 18092 31291
rect 19334 31288 19340 31340
rect 19392 31328 19398 31340
rect 19521 31331 19579 31337
rect 19521 31328 19533 31331
rect 19392 31300 19533 31328
rect 19392 31288 19398 31300
rect 19521 31297 19533 31300
rect 19567 31297 19579 31331
rect 19521 31291 19579 31297
rect 19679 31331 19737 31337
rect 19679 31297 19691 31331
rect 19725 31328 19737 31331
rect 19797 31331 19855 31337
rect 19725 31297 19748 31328
rect 19679 31291 19748 31297
rect 19797 31297 19809 31331
rect 19843 31297 19855 31331
rect 19797 31291 19855 31297
rect 17451 31232 18092 31260
rect 17451 31229 17463 31232
rect 17405 31223 17463 31229
rect 12526 31152 12532 31204
rect 12584 31192 12590 31204
rect 13648 31192 13676 31223
rect 12584 31164 13676 31192
rect 15841 31195 15899 31201
rect 12584 31152 12590 31164
rect 15841 31161 15853 31195
rect 15887 31192 15899 31195
rect 17034 31192 17040 31204
rect 15887 31164 17040 31192
rect 15887 31161 15899 31164
rect 15841 31155 15899 31161
rect 17034 31152 17040 31164
rect 17092 31152 17098 31204
rect 17313 31195 17371 31201
rect 17313 31161 17325 31195
rect 17359 31192 17371 31195
rect 17494 31192 17500 31204
rect 17359 31164 17500 31192
rect 17359 31161 17371 31164
rect 17313 31155 17371 31161
rect 17494 31152 17500 31164
rect 17552 31152 17558 31204
rect 19720 31192 19748 31291
rect 19812 31260 19840 31291
rect 19978 31288 19984 31340
rect 20036 31328 20042 31340
rect 24673 31331 24731 31337
rect 20036 31300 20081 31328
rect 20036 31288 20042 31300
rect 24673 31297 24685 31331
rect 24719 31297 24731 31331
rect 24673 31291 24731 31297
rect 20346 31260 20352 31272
rect 19812 31232 20352 31260
rect 20346 31220 20352 31232
rect 20404 31220 20410 31272
rect 24688 31260 24716 31291
rect 24762 31288 24768 31340
rect 24820 31328 24826 31340
rect 25133 31331 25191 31337
rect 24820 31300 24865 31328
rect 24820 31288 24826 31300
rect 25133 31297 25145 31331
rect 25179 31328 25191 31331
rect 25590 31328 25596 31340
rect 25179 31300 25596 31328
rect 25179 31297 25191 31300
rect 25133 31291 25191 31297
rect 25590 31288 25596 31300
rect 25648 31288 25654 31340
rect 25682 31288 25688 31340
rect 25740 31328 25746 31340
rect 25740 31300 25785 31328
rect 25740 31288 25746 31300
rect 25866 31288 25872 31340
rect 25924 31328 25930 31340
rect 28350 31328 28356 31340
rect 25924 31300 25969 31328
rect 28311 31300 28356 31328
rect 25924 31288 25930 31300
rect 28350 31288 28356 31300
rect 28408 31288 28414 31340
rect 28620 31331 28678 31337
rect 28620 31297 28632 31331
rect 28666 31328 28678 31331
rect 28902 31328 28908 31340
rect 28666 31300 28908 31328
rect 28666 31297 28678 31300
rect 28620 31291 28678 31297
rect 28902 31288 28908 31300
rect 28960 31288 28966 31340
rect 30208 31337 30236 31368
rect 31018 31356 31024 31368
rect 31076 31356 31082 31408
rect 35342 31396 35348 31408
rect 33704 31368 35348 31396
rect 30193 31331 30251 31337
rect 30193 31297 30205 31331
rect 30239 31297 30251 31331
rect 30193 31291 30251 31297
rect 30377 31331 30435 31337
rect 30377 31297 30389 31331
rect 30423 31297 30435 31331
rect 31294 31328 31300 31340
rect 31255 31300 31300 31328
rect 30377 31291 30435 31297
rect 25498 31260 25504 31272
rect 24688 31232 25504 31260
rect 25498 31220 25504 31232
rect 25556 31220 25562 31272
rect 22462 31192 22468 31204
rect 19720 31164 22468 31192
rect 22462 31152 22468 31164
rect 22520 31152 22526 31204
rect 25222 31192 25228 31204
rect 25056 31164 25228 31192
rect 9214 31124 9220 31136
rect 9175 31096 9220 31124
rect 9214 31084 9220 31096
rect 9272 31084 9278 31136
rect 10318 31124 10324 31136
rect 10279 31096 10324 31124
rect 10318 31084 10324 31096
rect 10376 31084 10382 31136
rect 10778 31084 10784 31136
rect 10836 31124 10842 31136
rect 12437 31127 12495 31133
rect 12437 31124 12449 31127
rect 10836 31096 12449 31124
rect 10836 31084 10842 31096
rect 12437 31093 12449 31096
rect 12483 31093 12495 31127
rect 15930 31124 15936 31136
rect 15891 31096 15936 31124
rect 12437 31087 12495 31093
rect 15930 31084 15936 31096
rect 15988 31084 15994 31136
rect 17862 31124 17868 31136
rect 17823 31096 17868 31124
rect 17862 31084 17868 31096
rect 17920 31084 17926 31136
rect 25056 31133 25084 31164
rect 25222 31152 25228 31164
rect 25280 31152 25286 31204
rect 30392 31192 30420 31291
rect 31294 31288 31300 31300
rect 31352 31288 31358 31340
rect 31481 31331 31539 31337
rect 31481 31297 31493 31331
rect 31527 31328 31539 31331
rect 31570 31328 31576 31340
rect 31527 31300 31576 31328
rect 31527 31297 31539 31300
rect 31481 31291 31539 31297
rect 31570 31288 31576 31300
rect 31628 31288 31634 31340
rect 33704 31337 33732 31368
rect 35342 31356 35348 31368
rect 35400 31356 35406 31408
rect 35621 31399 35679 31405
rect 35621 31365 35633 31399
rect 35667 31396 35679 31399
rect 36170 31396 36176 31408
rect 35667 31368 36176 31396
rect 35667 31365 35679 31368
rect 35621 31359 35679 31365
rect 36170 31356 36176 31368
rect 36228 31356 36234 31408
rect 37918 31396 37924 31408
rect 37660 31368 37924 31396
rect 33962 31337 33968 31340
rect 33689 31331 33747 31337
rect 33689 31297 33701 31331
rect 33735 31297 33747 31331
rect 33689 31291 33747 31297
rect 33956 31291 33968 31337
rect 34020 31328 34026 31340
rect 35526 31328 35532 31340
rect 34020 31300 34056 31328
rect 35487 31300 35532 31328
rect 33962 31288 33968 31291
rect 34020 31288 34026 31300
rect 35526 31288 35532 31300
rect 35584 31288 35590 31340
rect 35802 31328 35808 31340
rect 35715 31300 35808 31328
rect 35802 31288 35808 31300
rect 35860 31328 35866 31340
rect 37660 31328 37688 31368
rect 37918 31356 37924 31368
rect 37976 31356 37982 31408
rect 39390 31396 39396 31408
rect 39040 31368 39396 31396
rect 37826 31328 37832 31340
rect 35860 31300 37688 31328
rect 37787 31300 37832 31328
rect 35860 31288 35866 31300
rect 37826 31288 37832 31300
rect 37884 31328 37890 31340
rect 38378 31328 38384 31340
rect 37884 31300 38384 31328
rect 37884 31288 37890 31300
rect 38378 31288 38384 31300
rect 38436 31288 38442 31340
rect 39040 31337 39068 31368
rect 39390 31356 39396 31368
rect 39448 31356 39454 31408
rect 39025 31331 39083 31337
rect 39025 31297 39037 31331
rect 39071 31297 39083 31331
rect 39206 31328 39212 31340
rect 39167 31300 39212 31328
rect 39025 31291 39083 31297
rect 39206 31288 39212 31300
rect 39264 31288 39270 31340
rect 42610 31288 42616 31340
rect 42668 31328 42674 31340
rect 43145 31331 43203 31337
rect 43145 31328 43157 31331
rect 42668 31300 43157 31328
rect 42668 31288 42674 31300
rect 43145 31297 43157 31300
rect 43191 31297 43203 31331
rect 44726 31328 44732 31340
rect 44687 31300 44732 31328
rect 43145 31291 43203 31297
rect 44726 31288 44732 31300
rect 44784 31288 44790 31340
rect 37461 31263 37519 31269
rect 37461 31229 37473 31263
rect 37507 31260 37519 31263
rect 37642 31260 37648 31272
rect 37507 31232 37648 31260
rect 37507 31229 37519 31232
rect 37461 31223 37519 31229
rect 37642 31220 37648 31232
rect 37700 31220 37706 31272
rect 37734 31220 37740 31272
rect 37792 31260 37798 31272
rect 42886 31260 42892 31272
rect 37792 31232 37837 31260
rect 42847 31232 42892 31260
rect 37792 31220 37798 31232
rect 42886 31220 42892 31232
rect 42944 31220 42950 31272
rect 30392 31164 33732 31192
rect 25041 31127 25099 31133
rect 25041 31093 25053 31127
rect 25087 31093 25099 31127
rect 25041 31087 25099 31093
rect 25133 31127 25191 31133
rect 25133 31093 25145 31127
rect 25179 31124 25191 31127
rect 25406 31124 25412 31136
rect 25179 31096 25412 31124
rect 25179 31093 25191 31096
rect 25133 31087 25191 31093
rect 25406 31084 25412 31096
rect 25464 31084 25470 31136
rect 29730 31124 29736 31136
rect 29691 31096 29736 31124
rect 29730 31084 29736 31096
rect 29788 31084 29794 31136
rect 30282 31124 30288 31136
rect 30243 31096 30288 31124
rect 30282 31084 30288 31096
rect 30340 31084 30346 31136
rect 31481 31127 31539 31133
rect 31481 31093 31493 31127
rect 31527 31124 31539 31127
rect 33042 31124 33048 31136
rect 31527 31096 33048 31124
rect 31527 31093 31539 31096
rect 31481 31087 31539 31093
rect 33042 31084 33048 31096
rect 33100 31084 33106 31136
rect 33704 31124 33732 31164
rect 37458 31124 37464 31136
rect 33704 31096 37464 31124
rect 37458 31084 37464 31096
rect 37516 31084 37522 31136
rect 39114 31124 39120 31136
rect 39075 31096 39120 31124
rect 39114 31084 39120 31096
rect 39172 31084 39178 31136
rect 44910 31124 44916 31136
rect 44871 31096 44916 31124
rect 44910 31084 44916 31096
rect 44968 31084 44974 31136
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 13538 30880 13544 30932
rect 13596 30920 13602 30932
rect 13725 30923 13783 30929
rect 13725 30920 13737 30923
rect 13596 30892 13737 30920
rect 13596 30880 13602 30892
rect 13725 30889 13737 30892
rect 13771 30889 13783 30923
rect 15654 30920 15660 30932
rect 15615 30892 15660 30920
rect 13725 30883 13783 30889
rect 15654 30880 15660 30892
rect 15712 30880 15718 30932
rect 28902 30920 28908 30932
rect 28863 30892 28908 30920
rect 28902 30880 28908 30892
rect 28960 30880 28966 30932
rect 36449 30923 36507 30929
rect 36449 30889 36461 30923
rect 36495 30920 36507 30923
rect 37550 30920 37556 30932
rect 36495 30892 37556 30920
rect 36495 30889 36507 30892
rect 36449 30883 36507 30889
rect 37550 30880 37556 30892
rect 37608 30880 37614 30932
rect 42610 30920 42616 30932
rect 42571 30892 42616 30920
rect 42610 30880 42616 30892
rect 42668 30880 42674 30932
rect 45830 30880 45836 30932
rect 45888 30920 45894 30932
rect 46569 30923 46627 30929
rect 46569 30920 46581 30923
rect 45888 30892 46581 30920
rect 45888 30880 45894 30892
rect 46569 30889 46581 30892
rect 46615 30889 46627 30923
rect 46569 30883 46627 30889
rect 42886 30812 42892 30864
rect 42944 30852 42950 30864
rect 44082 30852 44088 30864
rect 42944 30824 44088 30852
rect 42944 30812 42950 30824
rect 44082 30812 44088 30824
rect 44140 30852 44146 30864
rect 44140 30824 45232 30852
rect 44140 30812 44146 30824
rect 6825 30787 6883 30793
rect 6825 30753 6837 30787
rect 6871 30784 6883 30787
rect 6914 30784 6920 30796
rect 6871 30756 6920 30784
rect 6871 30753 6883 30756
rect 6825 30747 6883 30753
rect 6914 30744 6920 30756
rect 6972 30744 6978 30796
rect 9766 30784 9772 30796
rect 8588 30756 9772 30784
rect 6089 30719 6147 30725
rect 6089 30685 6101 30719
rect 6135 30716 6147 30719
rect 7098 30716 7104 30728
rect 6135 30688 7104 30716
rect 6135 30685 6147 30688
rect 6089 30679 6147 30685
rect 7098 30676 7104 30688
rect 7156 30676 7162 30728
rect 8588 30725 8616 30756
rect 9766 30744 9772 30756
rect 9824 30744 9830 30796
rect 12342 30784 12348 30796
rect 12303 30756 12348 30784
rect 12342 30744 12348 30756
rect 12400 30744 12406 30796
rect 27338 30784 27344 30796
rect 25792 30756 27344 30784
rect 8573 30719 8631 30725
rect 8573 30685 8585 30719
rect 8619 30685 8631 30719
rect 8573 30679 8631 30685
rect 9306 30676 9312 30728
rect 9364 30716 9370 30728
rect 10778 30725 10784 30728
rect 9585 30719 9643 30725
rect 9585 30716 9597 30719
rect 9364 30688 9597 30716
rect 9364 30676 9370 30688
rect 9585 30685 9597 30688
rect 9631 30685 9643 30719
rect 9585 30679 9643 30685
rect 9861 30719 9919 30725
rect 9861 30685 9873 30719
rect 9907 30716 9919 30719
rect 10505 30719 10563 30725
rect 10505 30716 10517 30719
rect 9907 30688 10517 30716
rect 9907 30685 9919 30688
rect 9861 30679 9919 30685
rect 10505 30685 10517 30688
rect 10551 30685 10563 30719
rect 10772 30716 10784 30725
rect 10739 30688 10784 30716
rect 10505 30679 10563 30685
rect 10772 30679 10784 30688
rect 10778 30676 10784 30679
rect 10836 30676 10842 30728
rect 15841 30719 15899 30725
rect 15841 30685 15853 30719
rect 15887 30716 15899 30719
rect 15930 30716 15936 30728
rect 15887 30688 15936 30716
rect 15887 30685 15899 30688
rect 15841 30679 15899 30685
rect 15930 30676 15936 30688
rect 15988 30676 15994 30728
rect 17701 30719 17759 30725
rect 17701 30685 17713 30719
rect 17747 30716 17759 30719
rect 17862 30716 17868 30728
rect 17747 30688 17868 30716
rect 17747 30685 17759 30688
rect 17701 30679 17759 30685
rect 17862 30676 17868 30688
rect 17920 30676 17926 30728
rect 17957 30719 18015 30725
rect 17957 30685 17969 30719
rect 18003 30716 18015 30719
rect 18414 30716 18420 30728
rect 18003 30688 18420 30716
rect 18003 30685 18015 30688
rect 17957 30679 18015 30685
rect 18414 30676 18420 30688
rect 18472 30676 18478 30728
rect 25406 30716 25412 30728
rect 25367 30688 25412 30716
rect 25406 30676 25412 30688
rect 25464 30676 25470 30728
rect 25557 30719 25615 30725
rect 25557 30685 25569 30719
rect 25603 30716 25615 30719
rect 25792 30716 25820 30756
rect 27338 30744 27344 30756
rect 27396 30744 27402 30796
rect 30285 30787 30343 30793
rect 30285 30753 30297 30787
rect 30331 30784 30343 30787
rect 34698 30784 34704 30796
rect 30331 30756 34704 30784
rect 30331 30753 30343 30756
rect 30285 30747 30343 30753
rect 34698 30744 34704 30756
rect 34756 30744 34762 30796
rect 45204 30793 45232 30824
rect 43717 30787 43775 30793
rect 43717 30753 43729 30787
rect 43763 30753 43775 30787
rect 43717 30747 43775 30753
rect 45189 30787 45247 30793
rect 45189 30753 45201 30787
rect 45235 30753 45247 30787
rect 45189 30747 45247 30753
rect 25958 30725 25964 30728
rect 25603 30688 25820 30716
rect 25915 30719 25964 30725
rect 25603 30685 25615 30688
rect 25557 30679 25615 30685
rect 25915 30685 25927 30719
rect 25961 30685 25964 30719
rect 25915 30679 25964 30685
rect 25958 30676 25964 30679
rect 26016 30676 26022 30728
rect 29089 30719 29147 30725
rect 29089 30685 29101 30719
rect 29135 30716 29147 30719
rect 29135 30688 29776 30716
rect 29135 30685 29147 30688
rect 29089 30679 29147 30685
rect 7116 30648 7144 30676
rect 12434 30648 12440 30660
rect 7116 30620 12440 30648
rect 12434 30608 12440 30620
rect 12492 30608 12498 30660
rect 12612 30651 12670 30657
rect 12612 30617 12624 30651
rect 12658 30648 12670 30651
rect 12894 30648 12900 30660
rect 12658 30620 12900 30648
rect 12658 30617 12670 30620
rect 12612 30611 12670 30617
rect 12894 30608 12900 30620
rect 12952 30608 12958 30660
rect 25130 30608 25136 30660
rect 25188 30648 25194 30660
rect 25685 30651 25743 30657
rect 25685 30648 25697 30651
rect 25188 30620 25697 30648
rect 25188 30608 25194 30620
rect 25685 30617 25697 30620
rect 25731 30617 25743 30651
rect 25685 30611 25743 30617
rect 25777 30651 25835 30657
rect 25777 30617 25789 30651
rect 25823 30617 25835 30651
rect 25777 30611 25835 30617
rect 8386 30580 8392 30592
rect 8347 30552 8392 30580
rect 8386 30540 8392 30552
rect 8444 30540 8450 30592
rect 11885 30583 11943 30589
rect 11885 30549 11897 30583
rect 11931 30580 11943 30583
rect 12158 30580 12164 30592
rect 11931 30552 12164 30580
rect 11931 30549 11943 30552
rect 11885 30543 11943 30549
rect 12158 30540 12164 30552
rect 12216 30540 12222 30592
rect 16574 30540 16580 30592
rect 16632 30580 16638 30592
rect 16632 30552 16677 30580
rect 16632 30540 16638 30552
rect 23566 30540 23572 30592
rect 23624 30580 23630 30592
rect 25792 30580 25820 30611
rect 23624 30552 25820 30580
rect 26053 30583 26111 30589
rect 23624 30540 23630 30552
rect 26053 30549 26065 30583
rect 26099 30580 26111 30583
rect 26234 30580 26240 30592
rect 26099 30552 26240 30580
rect 26099 30549 26111 30552
rect 26053 30543 26111 30549
rect 26234 30540 26240 30552
rect 26292 30540 26298 30592
rect 29748 30589 29776 30688
rect 36906 30676 36912 30728
rect 36964 30716 36970 30728
rect 37182 30716 37188 30728
rect 36964 30688 37188 30716
rect 36964 30676 36970 30688
rect 37182 30676 37188 30688
rect 37240 30676 37246 30728
rect 37277 30719 37335 30725
rect 37277 30685 37289 30719
rect 37323 30685 37335 30719
rect 37458 30716 37464 30728
rect 37419 30688 37464 30716
rect 37277 30679 37335 30685
rect 36078 30648 36084 30660
rect 35991 30620 36084 30648
rect 36078 30608 36084 30620
rect 36136 30608 36142 30660
rect 36262 30648 36268 30660
rect 36223 30620 36268 30648
rect 36262 30608 36268 30620
rect 36320 30608 36326 30660
rect 37292 30648 37320 30679
rect 37458 30676 37464 30688
rect 37516 30676 37522 30728
rect 42429 30719 42487 30725
rect 42429 30685 42441 30719
rect 42475 30716 42487 30719
rect 43732 30716 43760 30747
rect 44450 30716 44456 30728
rect 42475 30688 43116 30716
rect 43732 30688 44456 30716
rect 42475 30685 42487 30688
rect 42429 30679 42487 30685
rect 37918 30648 37924 30660
rect 37292 30620 37924 30648
rect 37918 30608 37924 30620
rect 37976 30648 37982 30660
rect 37976 30620 41276 30648
rect 37976 30608 37982 30620
rect 29733 30583 29791 30589
rect 29733 30549 29745 30583
rect 29779 30549 29791 30583
rect 29733 30543 29791 30549
rect 29822 30540 29828 30592
rect 29880 30580 29886 30592
rect 30101 30583 30159 30589
rect 30101 30580 30113 30583
rect 29880 30552 30113 30580
rect 29880 30540 29886 30552
rect 30101 30549 30113 30552
rect 30147 30549 30159 30583
rect 30101 30543 30159 30549
rect 30190 30540 30196 30592
rect 30248 30580 30254 30592
rect 36096 30580 36124 30608
rect 41248 30592 41276 30620
rect 37826 30580 37832 30592
rect 30248 30552 30293 30580
rect 36096 30552 37832 30580
rect 30248 30540 30254 30552
rect 37826 30540 37832 30552
rect 37884 30540 37890 30592
rect 41230 30540 41236 30592
rect 41288 30580 41294 30592
rect 42794 30580 42800 30592
rect 41288 30552 42800 30580
rect 41288 30540 41294 30552
rect 42794 30540 42800 30552
rect 42852 30540 42858 30592
rect 43088 30589 43116 30688
rect 44450 30676 44456 30688
rect 44508 30676 44514 30728
rect 44637 30719 44695 30725
rect 44637 30685 44649 30719
rect 44683 30685 44695 30719
rect 44637 30679 44695 30685
rect 43441 30651 43499 30657
rect 43441 30617 43453 30651
rect 43487 30648 43499 30651
rect 44174 30648 44180 30660
rect 43487 30620 44180 30648
rect 43487 30617 43499 30620
rect 43441 30611 43499 30617
rect 44174 30608 44180 30620
rect 44232 30608 44238 30660
rect 44542 30608 44548 30660
rect 44600 30648 44606 30660
rect 44652 30648 44680 30679
rect 44910 30676 44916 30728
rect 44968 30716 44974 30728
rect 45445 30719 45503 30725
rect 45445 30716 45457 30719
rect 44968 30688 45457 30716
rect 44968 30676 44974 30688
rect 45445 30685 45457 30688
rect 45491 30685 45503 30719
rect 45445 30679 45503 30685
rect 45830 30648 45836 30660
rect 44600 30620 45836 30648
rect 44600 30608 44606 30620
rect 45830 30608 45836 30620
rect 45888 30608 45894 30660
rect 43073 30583 43131 30589
rect 43073 30549 43085 30583
rect 43119 30549 43131 30583
rect 43530 30580 43536 30592
rect 43491 30552 43536 30580
rect 43073 30543 43131 30549
rect 43530 30540 43536 30552
rect 43588 30540 43594 30592
rect 43714 30540 43720 30592
rect 43772 30580 43778 30592
rect 44269 30583 44327 30589
rect 44269 30580 44281 30583
rect 43772 30552 44281 30580
rect 43772 30540 43778 30552
rect 44269 30549 44281 30552
rect 44315 30549 44327 30583
rect 44269 30543 44327 30549
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 11698 30376 11704 30388
rect 11659 30348 11704 30376
rect 11698 30336 11704 30348
rect 11756 30336 11762 30388
rect 12894 30376 12900 30388
rect 12855 30348 12900 30376
rect 12894 30336 12900 30348
rect 12952 30336 12958 30388
rect 29917 30379 29975 30385
rect 22940 30348 25176 30376
rect 9668 30311 9726 30317
rect 6932 30280 9628 30308
rect 6932 30249 6960 30280
rect 6917 30243 6975 30249
rect 6917 30209 6929 30243
rect 6963 30209 6975 30243
rect 6917 30203 6975 30209
rect 9214 30200 9220 30252
rect 9272 30240 9278 30252
rect 9401 30243 9459 30249
rect 9401 30240 9413 30243
rect 9272 30212 9413 30240
rect 9272 30200 9278 30212
rect 9401 30209 9413 30212
rect 9447 30209 9459 30243
rect 9600 30240 9628 30280
rect 9668 30277 9680 30311
rect 9714 30308 9726 30311
rect 10318 30308 10324 30320
rect 9714 30280 10324 30308
rect 9714 30277 9726 30280
rect 9668 30271 9726 30277
rect 10318 30268 10324 30280
rect 10376 30268 10382 30320
rect 17681 30311 17739 30317
rect 11900 30280 16574 30308
rect 11900 30240 11928 30280
rect 9600 30212 11928 30240
rect 12069 30243 12127 30249
rect 9401 30203 9459 30209
rect 12069 30209 12081 30243
rect 12115 30240 12127 30243
rect 13078 30240 13084 30252
rect 12115 30212 12940 30240
rect 13039 30212 13084 30240
rect 12115 30209 12127 30212
rect 12069 30203 12127 30209
rect 6546 30132 6552 30184
rect 6604 30172 6610 30184
rect 6825 30175 6883 30181
rect 6825 30172 6837 30175
rect 6604 30144 6837 30172
rect 6604 30132 6610 30144
rect 6825 30141 6837 30144
rect 6871 30141 6883 30175
rect 12158 30172 12164 30184
rect 12119 30144 12164 30172
rect 6825 30135 6883 30141
rect 12158 30132 12164 30144
rect 12216 30132 12222 30184
rect 12253 30175 12311 30181
rect 12253 30141 12265 30175
rect 12299 30141 12311 30175
rect 12912 30172 12940 30212
rect 13078 30200 13084 30212
rect 13136 30200 13142 30252
rect 15470 30200 15476 30252
rect 15528 30240 15534 30252
rect 15565 30243 15623 30249
rect 15565 30240 15577 30243
rect 15528 30212 15577 30240
rect 15528 30200 15534 30212
rect 15565 30209 15577 30212
rect 15611 30209 15623 30243
rect 16546 30240 16574 30280
rect 17681 30277 17693 30311
rect 17727 30308 17739 30311
rect 18322 30308 18328 30320
rect 17727 30280 18328 30308
rect 17727 30277 17739 30280
rect 17681 30271 17739 30277
rect 18322 30268 18328 30280
rect 18380 30268 18386 30320
rect 22940 30308 22968 30348
rect 25148 30308 25176 30348
rect 29917 30345 29929 30379
rect 29963 30376 29975 30379
rect 30190 30376 30196 30388
rect 29963 30348 30196 30376
rect 29963 30345 29975 30348
rect 29917 30339 29975 30345
rect 30190 30336 30196 30348
rect 30248 30336 30254 30388
rect 40126 30376 40132 30388
rect 40184 30385 40190 30388
rect 40093 30348 40132 30376
rect 40126 30336 40132 30348
rect 40184 30339 40193 30385
rect 44174 30376 44180 30388
rect 44135 30348 44180 30376
rect 40184 30336 40190 30339
rect 44174 30336 44180 30348
rect 44232 30336 44238 30388
rect 39114 30308 39120 30320
rect 18432 30280 22968 30308
rect 23032 30280 25084 30308
rect 25148 30280 34744 30308
rect 18432 30240 18460 30280
rect 16546 30212 18460 30240
rect 15565 30203 15623 30209
rect 22094 30200 22100 30252
rect 22152 30240 22158 30252
rect 23032 30249 23060 30280
rect 23290 30249 23296 30252
rect 22189 30243 22247 30249
rect 22189 30240 22201 30243
rect 22152 30212 22201 30240
rect 22152 30200 22158 30212
rect 22189 30209 22201 30212
rect 22235 30209 22247 30243
rect 23017 30243 23075 30249
rect 23017 30240 23029 30243
rect 22189 30203 22247 30209
rect 22388 30212 23029 30240
rect 16574 30172 16580 30184
rect 12912 30144 16580 30172
rect 12253 30135 12311 30141
rect 10594 30064 10600 30116
rect 10652 30104 10658 30116
rect 10781 30107 10839 30113
rect 10781 30104 10793 30107
rect 10652 30076 10793 30104
rect 10652 30064 10658 30076
rect 10781 30073 10793 30076
rect 10827 30073 10839 30107
rect 12268 30104 12296 30135
rect 16574 30132 16580 30144
rect 16632 30172 16638 30184
rect 17862 30172 17868 30184
rect 16632 30144 17868 30172
rect 16632 30132 16638 30144
rect 17862 30132 17868 30144
rect 17920 30132 17926 30184
rect 18414 30172 18420 30184
rect 18375 30144 18420 30172
rect 18414 30132 18420 30144
rect 18472 30132 18478 30184
rect 22002 30132 22008 30184
rect 22060 30172 22066 30184
rect 22388 30172 22416 30212
rect 23017 30209 23029 30212
rect 23063 30209 23075 30243
rect 23017 30203 23075 30209
rect 23284 30203 23296 30249
rect 23348 30240 23354 30252
rect 23348 30212 23384 30240
rect 23290 30200 23296 30203
rect 23348 30200 23354 30212
rect 22060 30144 22416 30172
rect 22060 30132 22066 30144
rect 22462 30132 22468 30184
rect 22520 30172 22526 30184
rect 25056 30181 25084 30280
rect 25774 30240 25780 30252
rect 25735 30212 25780 30240
rect 25774 30200 25780 30212
rect 25832 30200 25838 30252
rect 27338 30240 27344 30252
rect 27299 30212 27344 30240
rect 27338 30200 27344 30212
rect 27396 30200 27402 30252
rect 29549 30243 29607 30249
rect 29549 30209 29561 30243
rect 29595 30240 29607 30243
rect 29730 30240 29736 30252
rect 29595 30212 29736 30240
rect 29595 30209 29607 30212
rect 29549 30203 29607 30209
rect 29730 30200 29736 30212
rect 29788 30200 29794 30252
rect 32490 30240 32496 30252
rect 32451 30212 32496 30240
rect 32490 30200 32496 30212
rect 32548 30200 32554 30252
rect 32674 30200 32680 30252
rect 32732 30240 32738 30252
rect 34330 30240 34336 30252
rect 32732 30212 34336 30240
rect 32732 30200 32738 30212
rect 34330 30200 34336 30212
rect 34388 30200 34394 30252
rect 34606 30240 34612 30252
rect 34567 30212 34612 30240
rect 34606 30200 34612 30212
rect 34664 30200 34670 30252
rect 25041 30175 25099 30181
rect 22520 30144 22565 30172
rect 22520 30132 22526 30144
rect 25041 30141 25053 30175
rect 25087 30172 25099 30175
rect 25958 30172 25964 30184
rect 25087 30144 25964 30172
rect 25087 30141 25099 30144
rect 25041 30135 25099 30141
rect 25958 30132 25964 30144
rect 26016 30132 26022 30184
rect 27522 30172 27528 30184
rect 27483 30144 27528 30172
rect 27522 30132 27528 30144
rect 27580 30132 27586 30184
rect 29641 30175 29699 30181
rect 29641 30141 29653 30175
rect 29687 30172 29699 30175
rect 30282 30172 30288 30184
rect 29687 30144 30288 30172
rect 29687 30141 29699 30144
rect 29641 30135 29699 30141
rect 30282 30132 30288 30144
rect 30340 30132 30346 30184
rect 31938 30132 31944 30184
rect 31996 30172 32002 30184
rect 32766 30172 32772 30184
rect 31996 30144 32772 30172
rect 31996 30132 32002 30144
rect 32766 30132 32772 30144
rect 32824 30132 32830 30184
rect 34716 30172 34744 30280
rect 34992 30280 35848 30308
rect 34790 30200 34796 30252
rect 34848 30240 34854 30252
rect 34848 30212 34893 30240
rect 34848 30200 34854 30212
rect 34992 30172 35020 30280
rect 35434 30240 35440 30252
rect 35395 30212 35440 30240
rect 35434 30200 35440 30212
rect 35492 30200 35498 30252
rect 35713 30243 35771 30249
rect 35713 30209 35725 30243
rect 35759 30209 35771 30243
rect 35713 30203 35771 30209
rect 34716 30144 35020 30172
rect 12434 30104 12440 30116
rect 10781 30067 10839 30073
rect 12176 30076 12440 30104
rect 6549 30039 6607 30045
rect 6549 30005 6561 30039
rect 6595 30036 6607 30039
rect 6730 30036 6736 30048
rect 6595 30008 6736 30036
rect 6595 30005 6607 30008
rect 6549 29999 6607 30005
rect 6730 29996 6736 30008
rect 6788 29996 6794 30048
rect 9306 29996 9312 30048
rect 9364 30036 9370 30048
rect 12176 30036 12204 30076
rect 12434 30064 12440 30076
rect 12492 30064 12498 30116
rect 18322 30064 18328 30116
rect 18380 30104 18386 30116
rect 24854 30104 24860 30116
rect 18380 30076 23060 30104
rect 18380 30064 18386 30076
rect 15378 30036 15384 30048
rect 9364 30008 12204 30036
rect 15339 30008 15384 30036
rect 9364 29996 9370 30008
rect 15378 29996 15384 30008
rect 15436 29996 15442 30048
rect 21542 29996 21548 30048
rect 21600 30036 21606 30048
rect 22005 30039 22063 30045
rect 22005 30036 22017 30039
rect 21600 30008 22017 30036
rect 21600 29996 21606 30008
rect 22005 30005 22017 30008
rect 22051 30005 22063 30039
rect 22370 30036 22376 30048
rect 22331 30008 22376 30036
rect 22005 29999 22063 30005
rect 22370 29996 22376 30008
rect 22428 29996 22434 30048
rect 23032 30036 23060 30076
rect 24320 30076 24860 30104
rect 24320 30036 24348 30076
rect 24854 30064 24860 30076
rect 24912 30104 24918 30116
rect 25774 30104 25780 30116
rect 24912 30076 25780 30104
rect 24912 30064 24918 30076
rect 25774 30064 25780 30076
rect 25832 30104 25838 30116
rect 28994 30104 29000 30116
rect 25832 30076 29000 30104
rect 25832 30064 25838 30076
rect 28994 30064 29000 30076
rect 29052 30064 29058 30116
rect 31570 30064 31576 30116
rect 31628 30104 31634 30116
rect 32677 30107 32735 30113
rect 32677 30104 32689 30107
rect 31628 30076 32689 30104
rect 31628 30064 31634 30076
rect 32677 30073 32689 30076
rect 32723 30073 32735 30107
rect 32677 30067 32735 30073
rect 33226 30064 33232 30116
rect 33284 30104 33290 30116
rect 34606 30104 34612 30116
rect 33284 30076 34612 30104
rect 33284 30064 33290 30076
rect 34606 30064 34612 30076
rect 34664 30104 34670 30116
rect 35728 30104 35756 30203
rect 34664 30076 35756 30104
rect 35820 30104 35848 30280
rect 38672 30280 39120 30308
rect 35897 30243 35955 30249
rect 35897 30209 35909 30243
rect 35943 30240 35955 30243
rect 36446 30240 36452 30252
rect 35943 30212 36452 30240
rect 35943 30209 35955 30212
rect 35897 30203 35955 30209
rect 36446 30200 36452 30212
rect 36504 30200 36510 30252
rect 37734 30200 37740 30252
rect 37792 30240 37798 30252
rect 38286 30240 38292 30252
rect 37792 30212 38292 30240
rect 37792 30200 37798 30212
rect 38286 30200 38292 30212
rect 38344 30240 38350 30252
rect 38672 30249 38700 30280
rect 39114 30268 39120 30280
rect 39172 30308 39178 30320
rect 40221 30311 40279 30317
rect 40221 30308 40233 30311
rect 39172 30280 40233 30308
rect 39172 30268 39178 30280
rect 40221 30277 40233 30280
rect 40267 30277 40279 30311
rect 44329 30311 44387 30317
rect 44329 30308 44341 30311
rect 40221 30271 40279 30277
rect 43272 30280 44341 30308
rect 38473 30243 38531 30249
rect 38473 30240 38485 30243
rect 38344 30212 38485 30240
rect 38344 30200 38350 30212
rect 38473 30209 38485 30212
rect 38519 30209 38531 30243
rect 38473 30203 38531 30209
rect 38657 30243 38715 30249
rect 38657 30209 38669 30243
rect 38703 30209 38715 30243
rect 38657 30203 38715 30209
rect 38838 30200 38844 30252
rect 38896 30240 38902 30252
rect 39577 30243 39635 30249
rect 39577 30240 39589 30243
rect 38896 30212 39589 30240
rect 38896 30200 38902 30212
rect 39577 30209 39589 30212
rect 39623 30209 39635 30243
rect 39577 30203 39635 30209
rect 40037 30243 40095 30249
rect 40037 30209 40049 30243
rect 40083 30209 40095 30243
rect 40037 30203 40095 30209
rect 40313 30243 40371 30249
rect 40313 30209 40325 30243
rect 40359 30240 40371 30243
rect 40678 30240 40684 30252
rect 40359 30212 40684 30240
rect 40359 30209 40371 30212
rect 40313 30203 40371 30209
rect 38378 30172 38384 30184
rect 38339 30144 38384 30172
rect 38378 30132 38384 30144
rect 38436 30132 38442 30184
rect 39206 30132 39212 30184
rect 39264 30172 39270 30184
rect 39301 30175 39359 30181
rect 39301 30172 39313 30175
rect 39264 30144 39313 30172
rect 39264 30132 39270 30144
rect 39301 30141 39313 30144
rect 39347 30141 39359 30175
rect 39482 30172 39488 30184
rect 39443 30144 39488 30172
rect 39301 30135 39359 30141
rect 39482 30132 39488 30144
rect 39540 30132 39546 30184
rect 40052 30104 40080 30203
rect 40678 30200 40684 30212
rect 40736 30200 40742 30252
rect 40770 30200 40776 30252
rect 40828 30240 40834 30252
rect 40957 30243 41015 30249
rect 40828 30212 40873 30240
rect 40828 30200 40834 30212
rect 40957 30209 40969 30243
rect 41003 30240 41015 30243
rect 41322 30240 41328 30252
rect 41003 30212 41328 30240
rect 41003 30209 41015 30212
rect 40957 30203 41015 30209
rect 40586 30132 40592 30184
rect 40644 30172 40650 30184
rect 40972 30172 41000 30203
rect 41322 30200 41328 30212
rect 41380 30200 41386 30252
rect 43272 30249 43300 30280
rect 44329 30277 44341 30280
rect 44375 30277 44387 30311
rect 44542 30308 44548 30320
rect 44503 30280 44548 30308
rect 44329 30271 44387 30277
rect 44542 30268 44548 30280
rect 44600 30268 44606 30320
rect 43257 30243 43315 30249
rect 43257 30209 43269 30243
rect 43303 30209 43315 30243
rect 43257 30203 43315 30209
rect 40644 30144 41000 30172
rect 43272 30172 43300 30203
rect 43346 30200 43352 30252
rect 43404 30240 43410 30252
rect 43533 30243 43591 30249
rect 43404 30212 43449 30240
rect 43404 30200 43410 30212
rect 43533 30209 43545 30243
rect 43579 30240 43591 30243
rect 44174 30240 44180 30252
rect 43579 30212 44180 30240
rect 43579 30209 43591 30212
rect 43533 30203 43591 30209
rect 44174 30200 44180 30212
rect 44232 30240 44238 30252
rect 44560 30240 44588 30268
rect 47762 30240 47768 30252
rect 44232 30212 44588 30240
rect 47723 30212 47768 30240
rect 44232 30200 44238 30212
rect 47762 30200 47768 30212
rect 47820 30200 47826 30252
rect 43438 30172 43444 30184
rect 43272 30144 43444 30172
rect 40644 30132 40650 30144
rect 43438 30132 43444 30144
rect 43496 30132 43502 30184
rect 40218 30104 40224 30116
rect 35820 30076 39528 30104
rect 40052 30076 40224 30104
rect 34664 30064 34670 30076
rect 23032 30008 24348 30036
rect 24397 30039 24455 30045
rect 24397 30005 24409 30039
rect 24443 30036 24455 30039
rect 24762 30036 24768 30048
rect 24443 30008 24768 30036
rect 24443 30005 24455 30008
rect 24397 29999 24455 30005
rect 24762 29996 24768 30008
rect 24820 29996 24826 30048
rect 25406 29996 25412 30048
rect 25464 30036 25470 30048
rect 27157 30039 27215 30045
rect 27157 30036 27169 30039
rect 25464 30008 27169 30036
rect 25464 29996 25470 30008
rect 27157 30005 27169 30008
rect 27203 30005 27215 30039
rect 32306 30036 32312 30048
rect 32267 30008 32312 30036
rect 27157 29999 27215 30005
rect 32306 29996 32312 30008
rect 32364 29996 32370 30048
rect 34054 29996 34060 30048
rect 34112 30036 34118 30048
rect 34149 30039 34207 30045
rect 34149 30036 34161 30039
rect 34112 30008 34161 30036
rect 34112 29996 34118 30008
rect 34149 30005 34161 30008
rect 34195 30005 34207 30039
rect 34149 29999 34207 30005
rect 34698 29996 34704 30048
rect 34756 30036 34762 30048
rect 35253 30039 35311 30045
rect 35253 30036 35265 30039
rect 34756 30008 35265 30036
rect 34756 29996 34762 30008
rect 35253 30005 35265 30008
rect 35299 30005 35311 30039
rect 35728 30036 35756 30076
rect 36630 30036 36636 30048
rect 35728 30008 36636 30036
rect 35253 29999 35311 30005
rect 36630 29996 36636 30008
rect 36688 29996 36694 30048
rect 38838 30036 38844 30048
rect 38799 30008 38844 30036
rect 38838 29996 38844 30008
rect 38896 29996 38902 30048
rect 38930 29996 38936 30048
rect 38988 30036 38994 30048
rect 39393 30039 39451 30045
rect 39393 30036 39405 30039
rect 38988 30008 39405 30036
rect 38988 29996 38994 30008
rect 39393 30005 39405 30008
rect 39439 30005 39451 30039
rect 39500 30036 39528 30076
rect 40218 30064 40224 30076
rect 40276 30104 40282 30116
rect 40773 30107 40831 30113
rect 40773 30104 40785 30107
rect 40276 30076 40785 30104
rect 40276 30064 40282 30076
rect 40773 30073 40785 30076
rect 40819 30073 40831 30107
rect 40773 30067 40831 30073
rect 43162 30064 43168 30116
rect 43220 30104 43226 30116
rect 43346 30104 43352 30116
rect 43220 30076 43352 30104
rect 43220 30064 43226 30076
rect 43346 30064 43352 30076
rect 43404 30104 43410 30116
rect 43404 30076 44404 30104
rect 43404 30064 43410 30076
rect 43254 30036 43260 30048
rect 39500 30008 43260 30036
rect 39393 29999 39451 30005
rect 43254 29996 43260 30008
rect 43312 29996 43318 30048
rect 43717 30039 43775 30045
rect 43717 30005 43729 30039
rect 43763 30036 43775 30039
rect 43898 30036 43904 30048
rect 43763 30008 43904 30036
rect 43763 30005 43775 30008
rect 43717 29999 43775 30005
rect 43898 29996 43904 30008
rect 43956 29996 43962 30048
rect 44376 30045 44404 30076
rect 44361 30039 44419 30045
rect 44361 30005 44373 30039
rect 44407 30005 44419 30039
rect 44361 29999 44419 30005
rect 46474 29996 46480 30048
rect 46532 30036 46538 30048
rect 47029 30039 47087 30045
rect 47029 30036 47041 30039
rect 46532 30008 47041 30036
rect 46532 29996 46538 30008
rect 47029 30005 47041 30008
rect 47075 30005 47087 30039
rect 47854 30036 47860 30048
rect 47815 30008 47860 30036
rect 47029 29999 47087 30005
rect 47854 29996 47860 30008
rect 47912 29996 47918 30048
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 5166 29792 5172 29844
rect 5224 29832 5230 29844
rect 6822 29832 6828 29844
rect 5224 29804 6828 29832
rect 5224 29792 5230 29804
rect 6822 29792 6828 29804
rect 6880 29832 6886 29844
rect 44085 29835 44143 29841
rect 6880 29804 44036 29832
rect 6880 29792 6886 29804
rect 198 29724 204 29776
rect 256 29764 262 29776
rect 13078 29764 13084 29776
rect 256 29736 6914 29764
rect 13039 29736 13084 29764
rect 256 29724 262 29736
rect 6730 29696 6736 29708
rect 6691 29668 6736 29696
rect 6730 29656 6736 29668
rect 6788 29656 6794 29708
rect 6886 29696 6914 29736
rect 13078 29724 13084 29736
rect 13136 29724 13142 29776
rect 17494 29764 17500 29776
rect 17455 29736 17500 29764
rect 17494 29724 17500 29736
rect 17552 29724 17558 29776
rect 23290 29764 23296 29776
rect 23251 29736 23296 29764
rect 23290 29724 23296 29736
rect 23348 29724 23354 29776
rect 25498 29764 25504 29776
rect 25148 29736 25504 29764
rect 7193 29699 7251 29705
rect 7193 29696 7205 29699
rect 6886 29668 7205 29696
rect 7193 29665 7205 29668
rect 7239 29665 7251 29699
rect 7193 29659 7251 29665
rect 10965 29699 11023 29705
rect 10965 29665 10977 29699
rect 11011 29696 11023 29699
rect 12158 29696 12164 29708
rect 11011 29668 12164 29696
rect 11011 29665 11023 29668
rect 10965 29659 11023 29665
rect 12158 29656 12164 29668
rect 12216 29656 12222 29708
rect 12434 29696 12440 29708
rect 12395 29668 12440 29696
rect 12434 29656 12440 29668
rect 12492 29656 12498 29708
rect 17770 29656 17776 29708
rect 17828 29696 17834 29708
rect 18049 29699 18107 29705
rect 18049 29696 18061 29699
rect 17828 29668 18061 29696
rect 17828 29656 17834 29668
rect 18049 29665 18061 29668
rect 18095 29665 18107 29699
rect 19242 29696 19248 29708
rect 18049 29659 18107 29665
rect 18432 29668 19248 29696
rect 18432 29640 18460 29668
rect 19242 29656 19248 29668
rect 19300 29656 19306 29708
rect 20898 29696 20904 29708
rect 19628 29668 20904 29696
rect 10594 29588 10600 29640
rect 10652 29628 10658 29640
rect 10873 29631 10931 29637
rect 10873 29628 10885 29631
rect 10652 29600 10885 29628
rect 10652 29588 10658 29600
rect 10873 29597 10885 29600
rect 10919 29597 10931 29631
rect 14274 29628 14280 29640
rect 14235 29600 14280 29628
rect 10873 29591 10931 29597
rect 14274 29588 14280 29600
rect 14332 29588 14338 29640
rect 14734 29588 14740 29640
rect 14792 29628 14798 29640
rect 15013 29631 15071 29637
rect 15013 29628 15025 29631
rect 14792 29600 15025 29628
rect 14792 29588 14798 29600
rect 15013 29597 15025 29600
rect 15059 29628 15071 29631
rect 18414 29628 18420 29640
rect 15059 29600 18420 29628
rect 15059 29597 15071 29600
rect 15013 29591 15071 29597
rect 18414 29588 18420 29600
rect 18472 29588 18478 29640
rect 18598 29588 18604 29640
rect 18656 29628 18662 29640
rect 19628 29637 19656 29668
rect 20898 29656 20904 29668
rect 20956 29656 20962 29708
rect 22462 29656 22468 29708
rect 22520 29696 22526 29708
rect 24946 29696 24952 29708
rect 22520 29668 24952 29696
rect 22520 29656 22526 29668
rect 24946 29656 24952 29668
rect 25004 29656 25010 29708
rect 25148 29705 25176 29736
rect 25498 29724 25504 29736
rect 25556 29724 25562 29776
rect 27338 29764 27344 29776
rect 27299 29736 27344 29764
rect 27338 29724 27344 29736
rect 27396 29724 27402 29776
rect 32858 29764 32864 29776
rect 32819 29736 32864 29764
rect 32858 29724 32864 29736
rect 32916 29724 32922 29776
rect 33873 29767 33931 29773
rect 33873 29733 33885 29767
rect 33919 29764 33931 29767
rect 33962 29764 33968 29776
rect 33919 29736 33968 29764
rect 33919 29733 33931 29736
rect 33873 29727 33931 29733
rect 33962 29724 33968 29736
rect 34020 29724 34026 29776
rect 42889 29767 42947 29773
rect 42889 29733 42901 29767
rect 42935 29764 42947 29767
rect 44008 29764 44036 29804
rect 44085 29801 44097 29835
rect 44131 29832 44143 29835
rect 44726 29832 44732 29844
rect 44131 29804 44732 29832
rect 44131 29801 44143 29804
rect 44085 29795 44143 29801
rect 44726 29792 44732 29804
rect 44784 29792 44790 29844
rect 44634 29764 44640 29776
rect 42935 29736 43576 29764
rect 44008 29736 44640 29764
rect 42935 29733 42947 29736
rect 42889 29727 42947 29733
rect 43548 29708 43576 29736
rect 44634 29724 44640 29736
rect 44692 29724 44698 29776
rect 25133 29699 25191 29705
rect 25133 29665 25145 29699
rect 25179 29665 25191 29699
rect 25406 29696 25412 29708
rect 25367 29668 25412 29696
rect 25133 29659 25191 29665
rect 25406 29656 25412 29668
rect 25464 29656 25470 29708
rect 25958 29696 25964 29708
rect 25919 29668 25964 29696
rect 25958 29656 25964 29668
rect 26016 29656 26022 29708
rect 29638 29656 29644 29708
rect 29696 29696 29702 29708
rect 35342 29696 35348 29708
rect 29696 29668 30236 29696
rect 29696 29656 29702 29668
rect 19429 29631 19487 29637
rect 19429 29628 19441 29631
rect 18656 29600 19441 29628
rect 18656 29588 18662 29600
rect 19429 29597 19441 29600
rect 19475 29597 19487 29631
rect 19429 29591 19487 29597
rect 19613 29631 19671 29637
rect 19613 29597 19625 29631
rect 19659 29597 19671 29631
rect 19613 29591 19671 29597
rect 19889 29631 19947 29637
rect 19889 29597 19901 29631
rect 19935 29628 19947 29631
rect 20622 29628 20628 29640
rect 19935 29600 20628 29628
rect 19935 29597 19947 29600
rect 19889 29591 19947 29597
rect 20622 29588 20628 29600
rect 20680 29588 20686 29640
rect 21269 29631 21327 29637
rect 21269 29597 21281 29631
rect 21315 29628 21327 29631
rect 22002 29628 22008 29640
rect 21315 29600 22008 29628
rect 21315 29597 21327 29600
rect 21269 29591 21327 29597
rect 22002 29588 22008 29600
rect 22060 29588 22066 29640
rect 23474 29628 23480 29640
rect 23435 29600 23480 29628
rect 23474 29588 23480 29600
rect 23532 29588 23538 29640
rect 24762 29588 24768 29640
rect 24820 29628 24826 29640
rect 25225 29631 25283 29637
rect 25225 29628 25237 29631
rect 24820 29600 25237 29628
rect 24820 29588 24826 29600
rect 25225 29597 25237 29600
rect 25271 29597 25283 29631
rect 25225 29591 25283 29597
rect 25317 29631 25375 29637
rect 25317 29597 25329 29631
rect 25363 29628 25375 29631
rect 25774 29628 25780 29640
rect 25363 29600 25780 29628
rect 25363 29597 25375 29600
rect 25317 29591 25375 29597
rect 25774 29588 25780 29600
rect 25832 29588 25838 29640
rect 26234 29637 26240 29640
rect 26228 29628 26240 29637
rect 26195 29600 26240 29628
rect 26228 29591 26240 29600
rect 26234 29588 26240 29591
rect 26292 29588 26298 29640
rect 29733 29631 29791 29637
rect 29733 29597 29745 29631
rect 29779 29628 29791 29631
rect 29822 29628 29828 29640
rect 29779 29600 29828 29628
rect 29779 29597 29791 29600
rect 29733 29591 29791 29597
rect 29822 29588 29828 29600
rect 29880 29588 29886 29640
rect 29917 29631 29975 29637
rect 29917 29597 29929 29631
rect 29963 29628 29975 29631
rect 30098 29628 30104 29640
rect 29963 29600 30104 29628
rect 29963 29597 29975 29600
rect 29917 29591 29975 29597
rect 30098 29588 30104 29600
rect 30156 29588 30162 29640
rect 30208 29637 30236 29668
rect 33980 29668 35348 29696
rect 30193 29631 30251 29637
rect 30193 29597 30205 29631
rect 30239 29628 30251 29631
rect 31018 29628 31024 29640
rect 30239 29600 31024 29628
rect 30239 29597 30251 29600
rect 30193 29591 30251 29597
rect 31018 29588 31024 29600
rect 31076 29588 31082 29640
rect 31481 29631 31539 29637
rect 31481 29597 31493 29631
rect 31527 29628 31539 29631
rect 33980 29628 34008 29668
rect 35342 29656 35348 29668
rect 35400 29696 35406 29708
rect 35621 29699 35679 29705
rect 35621 29696 35633 29699
rect 35400 29668 35633 29696
rect 35400 29656 35406 29668
rect 35621 29665 35633 29668
rect 35667 29665 35679 29699
rect 37366 29696 37372 29708
rect 35621 29659 35679 29665
rect 35728 29668 37372 29696
rect 31527 29600 34008 29628
rect 31527 29597 31539 29600
rect 31481 29591 31539 29597
rect 34054 29588 34060 29640
rect 34112 29628 34118 29640
rect 34241 29631 34299 29637
rect 34112 29600 34157 29628
rect 34112 29588 34118 29600
rect 34241 29597 34253 29631
rect 34287 29597 34299 29631
rect 34241 29591 34299 29597
rect 6914 29520 6920 29572
rect 6972 29560 6978 29572
rect 12713 29563 12771 29569
rect 6972 29532 7017 29560
rect 6972 29520 6978 29532
rect 12713 29529 12725 29563
rect 12759 29560 12771 29563
rect 15280 29563 15338 29569
rect 12759 29532 15240 29560
rect 12759 29529 12771 29532
rect 12713 29523 12771 29529
rect 10226 29452 10232 29504
rect 10284 29492 10290 29504
rect 10505 29495 10563 29501
rect 10505 29492 10517 29495
rect 10284 29464 10517 29492
rect 10284 29452 10290 29464
rect 10505 29461 10517 29464
rect 10551 29461 10563 29495
rect 12618 29492 12624 29504
rect 12579 29464 12624 29492
rect 10505 29455 10563 29461
rect 12618 29452 12624 29464
rect 12676 29452 12682 29504
rect 14458 29492 14464 29504
rect 14419 29464 14464 29492
rect 14458 29452 14464 29464
rect 14516 29452 14522 29504
rect 15212 29492 15240 29532
rect 15280 29529 15292 29563
rect 15326 29560 15338 29563
rect 15378 29560 15384 29572
rect 15326 29532 15384 29560
rect 15326 29529 15338 29532
rect 15280 29523 15338 29529
rect 15378 29520 15384 29532
rect 15436 29520 15442 29572
rect 17862 29560 17868 29572
rect 17823 29532 17868 29560
rect 17862 29520 17868 29532
rect 17920 29520 17926 29572
rect 21542 29569 21548 29572
rect 17957 29563 18015 29569
rect 17957 29529 17969 29563
rect 18003 29560 18015 29563
rect 21536 29560 21548 29569
rect 18003 29532 21404 29560
rect 21503 29532 21548 29560
rect 18003 29529 18015 29532
rect 17957 29523 18015 29529
rect 16393 29495 16451 29501
rect 16393 29492 16405 29495
rect 15212 29464 16405 29492
rect 16393 29461 16405 29464
rect 16439 29492 16451 29495
rect 17218 29492 17224 29504
rect 16439 29464 17224 29492
rect 16439 29461 16451 29464
rect 16393 29455 16451 29461
rect 17218 29452 17224 29464
rect 17276 29452 17282 29504
rect 19978 29452 19984 29504
rect 20036 29492 20042 29504
rect 20073 29495 20131 29501
rect 20073 29492 20085 29495
rect 20036 29464 20085 29492
rect 20036 29452 20042 29464
rect 20073 29461 20085 29464
rect 20119 29461 20131 29495
rect 21376 29492 21404 29532
rect 21536 29523 21548 29532
rect 21542 29520 21548 29523
rect 21600 29520 21606 29572
rect 31748 29563 31806 29569
rect 22066 29532 30604 29560
rect 22066 29492 22094 29532
rect 21376 29464 22094 29492
rect 22649 29495 22707 29501
rect 20073 29455 20131 29461
rect 22649 29461 22661 29495
rect 22695 29492 22707 29495
rect 23566 29492 23572 29504
rect 22695 29464 23572 29492
rect 22695 29461 22707 29464
rect 22649 29455 22707 29461
rect 23566 29452 23572 29464
rect 23624 29452 23630 29504
rect 23842 29452 23848 29504
rect 23900 29492 23906 29504
rect 24949 29495 25007 29501
rect 24949 29492 24961 29495
rect 23900 29464 24961 29492
rect 23900 29452 23906 29464
rect 24949 29461 24961 29464
rect 24995 29461 25007 29495
rect 24949 29455 25007 29461
rect 25038 29452 25044 29504
rect 25096 29492 25102 29504
rect 27614 29492 27620 29504
rect 25096 29464 27620 29492
rect 25096 29452 25102 29464
rect 27614 29452 27620 29464
rect 27672 29492 27678 29504
rect 29086 29492 29092 29504
rect 27672 29464 29092 29492
rect 27672 29452 27678 29464
rect 29086 29452 29092 29464
rect 29144 29452 29150 29504
rect 30377 29495 30435 29501
rect 30377 29461 30389 29495
rect 30423 29492 30435 29495
rect 30466 29492 30472 29504
rect 30423 29464 30472 29492
rect 30423 29461 30435 29464
rect 30377 29455 30435 29461
rect 30466 29452 30472 29464
rect 30524 29452 30530 29504
rect 30576 29492 30604 29532
rect 31748 29529 31760 29563
rect 31794 29560 31806 29563
rect 32306 29560 32312 29572
rect 31794 29532 32312 29560
rect 31794 29529 31806 29532
rect 31748 29523 31806 29529
rect 32306 29520 32312 29532
rect 32364 29520 32370 29572
rect 33502 29520 33508 29572
rect 33560 29560 33566 29572
rect 34256 29560 34284 29591
rect 34330 29588 34336 29640
rect 34388 29628 34394 29640
rect 35728 29628 35756 29668
rect 37366 29656 37372 29668
rect 37424 29656 37430 29708
rect 37921 29699 37979 29705
rect 37921 29665 37933 29699
rect 37967 29696 37979 29699
rect 40034 29696 40040 29708
rect 37967 29668 39896 29696
rect 39995 29668 40040 29696
rect 37967 29665 37979 29668
rect 37921 29659 37979 29665
rect 34388 29600 35756 29628
rect 34388 29588 34394 29600
rect 36446 29588 36452 29640
rect 36504 29628 36510 29640
rect 37645 29631 37703 29637
rect 37645 29628 37657 29631
rect 36504 29600 37657 29628
rect 36504 29588 36510 29600
rect 37645 29597 37657 29600
rect 37691 29597 37703 29631
rect 37826 29628 37832 29640
rect 37787 29600 37832 29628
rect 37645 29591 37703 29597
rect 37826 29588 37832 29600
rect 37884 29588 37890 29640
rect 38010 29628 38016 29640
rect 37971 29600 38016 29628
rect 38010 29588 38016 29600
rect 38068 29588 38074 29640
rect 38197 29631 38255 29637
rect 38197 29597 38209 29631
rect 38243 29628 38255 29631
rect 38657 29631 38715 29637
rect 38657 29628 38669 29631
rect 38243 29600 38669 29628
rect 38243 29597 38255 29600
rect 38197 29591 38255 29597
rect 38657 29597 38669 29600
rect 38703 29597 38715 29631
rect 38657 29591 38715 29597
rect 38841 29631 38899 29637
rect 38841 29597 38853 29631
rect 38887 29628 38899 29631
rect 38930 29628 38936 29640
rect 38887 29600 38936 29628
rect 38887 29597 38899 29600
rect 38841 29591 38899 29597
rect 38930 29588 38936 29600
rect 38988 29588 38994 29640
rect 39114 29628 39120 29640
rect 39075 29600 39120 29628
rect 39114 29588 39120 29600
rect 39172 29628 39178 29640
rect 39482 29628 39488 29640
rect 39172 29600 39488 29628
rect 39172 29588 39178 29600
rect 39482 29588 39488 29600
rect 39540 29588 39546 29640
rect 39868 29628 39896 29668
rect 40034 29656 40040 29668
rect 40092 29656 40098 29708
rect 42978 29656 42984 29708
rect 43036 29696 43042 29708
rect 43073 29699 43131 29705
rect 43073 29696 43085 29699
rect 43036 29668 43085 29696
rect 43036 29656 43042 29668
rect 43073 29665 43085 29668
rect 43119 29665 43131 29699
rect 43073 29659 43131 29665
rect 43530 29656 43536 29708
rect 43588 29696 43594 29708
rect 43717 29699 43775 29705
rect 43717 29696 43729 29699
rect 43588 29668 43729 29696
rect 43588 29656 43594 29668
rect 43717 29665 43729 29668
rect 43763 29665 43775 29699
rect 46474 29696 46480 29708
rect 46435 29668 46480 29696
rect 43717 29659 43775 29665
rect 46474 29656 46480 29668
rect 46532 29656 46538 29708
rect 46661 29699 46719 29705
rect 46661 29665 46673 29699
rect 46707 29696 46719 29699
rect 47854 29696 47860 29708
rect 46707 29668 47860 29696
rect 46707 29665 46719 29668
rect 46661 29659 46719 29665
rect 47854 29656 47860 29668
rect 47912 29656 47918 29708
rect 40770 29628 40776 29640
rect 39868 29600 40776 29628
rect 40770 29588 40776 29600
rect 40828 29628 40834 29640
rect 42886 29628 42892 29640
rect 40828 29600 41460 29628
rect 42847 29600 42892 29628
rect 40828 29588 40834 29600
rect 33560 29532 34284 29560
rect 33560 29520 33566 29532
rect 34790 29520 34796 29572
rect 34848 29560 34854 29572
rect 34885 29563 34943 29569
rect 34885 29560 34897 29563
rect 34848 29532 34897 29560
rect 34848 29520 34854 29532
rect 34885 29529 34897 29532
rect 34931 29529 34943 29563
rect 34885 29523 34943 29529
rect 37461 29563 37519 29569
rect 37461 29529 37473 29563
rect 37507 29560 37519 29563
rect 40282 29563 40340 29569
rect 40282 29560 40294 29563
rect 37507 29532 40294 29560
rect 37507 29529 37519 29532
rect 37461 29523 37519 29529
rect 40282 29529 40294 29532
rect 40328 29529 40340 29563
rect 40282 29523 40340 29529
rect 33318 29492 33324 29504
rect 30576 29464 33324 29492
rect 33318 29452 33324 29464
rect 33376 29452 33382 29504
rect 33410 29452 33416 29504
rect 33468 29492 33474 29504
rect 38654 29492 38660 29504
rect 33468 29464 38660 29492
rect 33468 29452 33474 29464
rect 38654 29452 38660 29464
rect 38712 29452 38718 29504
rect 38838 29452 38844 29504
rect 38896 29492 38902 29504
rect 39025 29495 39083 29501
rect 39025 29492 39037 29495
rect 38896 29464 39037 29492
rect 38896 29452 38902 29464
rect 39025 29461 39037 29464
rect 39071 29492 39083 29495
rect 40494 29492 40500 29504
rect 39071 29464 40500 29492
rect 39071 29461 39083 29464
rect 39025 29455 39083 29461
rect 40494 29452 40500 29464
rect 40552 29452 40558 29504
rect 41432 29501 41460 29600
rect 42886 29588 42892 29600
rect 42944 29588 42950 29640
rect 43257 29631 43315 29637
rect 43257 29597 43269 29631
rect 43303 29628 43315 29631
rect 43438 29628 43444 29640
rect 43303 29600 43444 29628
rect 43303 29597 43315 29600
rect 43257 29591 43315 29597
rect 43438 29588 43444 29600
rect 43496 29588 43502 29640
rect 43898 29628 43904 29640
rect 43859 29600 43904 29628
rect 43898 29588 43904 29600
rect 43956 29588 43962 29640
rect 43165 29563 43223 29569
rect 43165 29529 43177 29563
rect 43211 29560 43223 29563
rect 44174 29560 44180 29572
rect 43211 29532 44180 29560
rect 43211 29529 43223 29532
rect 43165 29523 43223 29529
rect 44174 29520 44180 29532
rect 44232 29520 44238 29572
rect 48314 29560 48320 29572
rect 48275 29532 48320 29560
rect 48314 29520 48320 29532
rect 48372 29520 48378 29572
rect 41417 29495 41475 29501
rect 41417 29461 41429 29495
rect 41463 29461 41475 29495
rect 41417 29455 41475 29461
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 6825 29291 6883 29297
rect 6825 29257 6837 29291
rect 6871 29288 6883 29291
rect 6914 29288 6920 29300
rect 6871 29260 6920 29288
rect 6871 29257 6883 29260
rect 6825 29251 6883 29257
rect 6914 29248 6920 29260
rect 6972 29248 6978 29300
rect 13262 29248 13268 29300
rect 13320 29288 13326 29300
rect 15470 29288 15476 29300
rect 13320 29260 14688 29288
rect 15431 29260 15476 29288
rect 13320 29248 13326 29260
rect 8386 29229 8392 29232
rect 8380 29220 8392 29229
rect 8347 29192 8392 29220
rect 8380 29183 8392 29192
rect 8386 29180 8392 29183
rect 8444 29180 8450 29232
rect 14458 29180 14464 29232
rect 14516 29229 14522 29232
rect 14516 29220 14528 29229
rect 14660 29220 14688 29260
rect 15470 29248 15476 29260
rect 15528 29248 15534 29300
rect 15654 29248 15660 29300
rect 15712 29288 15718 29300
rect 29638 29288 29644 29300
rect 15712 29260 29644 29288
rect 15712 29248 15718 29260
rect 29638 29248 29644 29260
rect 29696 29248 29702 29300
rect 29822 29288 29828 29300
rect 29783 29260 29828 29288
rect 29822 29248 29828 29260
rect 29880 29248 29886 29300
rect 33318 29248 33324 29300
rect 33376 29288 33382 29300
rect 34146 29288 34152 29300
rect 33376 29260 34152 29288
rect 33376 29248 33382 29260
rect 34146 29248 34152 29260
rect 34204 29248 34210 29300
rect 34256 29260 47256 29288
rect 19092 29223 19150 29229
rect 14516 29192 14561 29220
rect 14660 29192 18368 29220
rect 14516 29183 14528 29192
rect 14516 29180 14522 29183
rect 5626 29152 5632 29164
rect 5587 29124 5632 29152
rect 5626 29112 5632 29124
rect 5684 29112 5690 29164
rect 6733 29155 6791 29161
rect 6733 29121 6745 29155
rect 6779 29152 6791 29155
rect 6822 29152 6828 29164
rect 6779 29124 6828 29152
rect 6779 29121 6791 29124
rect 6733 29115 6791 29121
rect 6822 29112 6828 29124
rect 6880 29112 6886 29164
rect 15654 29152 15660 29164
rect 15567 29124 15660 29152
rect 15654 29112 15660 29124
rect 15712 29112 15718 29164
rect 15841 29155 15899 29161
rect 15841 29121 15853 29155
rect 15887 29152 15899 29155
rect 16850 29152 16856 29164
rect 15887 29124 16856 29152
rect 15887 29121 15899 29124
rect 15841 29115 15899 29121
rect 16850 29112 16856 29124
rect 16908 29112 16914 29164
rect 18340 29152 18368 29192
rect 19092 29189 19104 29223
rect 19138 29220 19150 29223
rect 19426 29220 19432 29232
rect 19138 29192 19432 29220
rect 19138 29189 19150 29192
rect 19092 29183 19150 29189
rect 19426 29180 19432 29192
rect 19484 29180 19490 29232
rect 32030 29220 32036 29232
rect 19904 29192 32036 29220
rect 18340 29124 19288 29152
rect 8110 29084 8116 29096
rect 8071 29056 8116 29084
rect 8110 29044 8116 29056
rect 8168 29044 8174 29096
rect 14734 29084 14740 29096
rect 14695 29056 14740 29084
rect 14734 29044 14740 29056
rect 14792 29044 14798 29096
rect 5537 29019 5595 29025
rect 5537 28985 5549 29019
rect 5583 29016 5595 29019
rect 6914 29016 6920 29028
rect 5583 28988 6920 29016
rect 5583 28985 5595 28988
rect 5537 28979 5595 28985
rect 6914 28976 6920 28988
rect 6972 28976 6978 29028
rect 12710 28976 12716 29028
rect 12768 29016 12774 29028
rect 13357 29019 13415 29025
rect 13357 29016 13369 29019
rect 12768 28988 13369 29016
rect 12768 28976 12774 28988
rect 13357 28985 13369 28988
rect 13403 28985 13415 29019
rect 13357 28979 13415 28985
rect 9490 28948 9496 28960
rect 9451 28920 9496 28948
rect 9490 28908 9496 28920
rect 9548 28908 9554 28960
rect 13538 28908 13544 28960
rect 13596 28948 13602 28960
rect 15672 28948 15700 29112
rect 19260 29084 19288 29124
rect 19334 29112 19340 29164
rect 19392 29152 19398 29164
rect 19797 29155 19855 29161
rect 19797 29152 19809 29155
rect 19392 29124 19809 29152
rect 19392 29112 19398 29124
rect 19797 29121 19809 29124
rect 19843 29121 19855 29155
rect 19797 29115 19855 29121
rect 19904 29084 19932 29192
rect 32030 29180 32036 29192
rect 32088 29180 32094 29232
rect 32398 29180 32404 29232
rect 32456 29220 32462 29232
rect 34256 29220 34284 29260
rect 35342 29220 35348 29232
rect 32456 29192 34284 29220
rect 34348 29192 35348 29220
rect 32456 29180 32462 29192
rect 20070 29161 20076 29164
rect 20064 29115 20076 29161
rect 20128 29152 20134 29164
rect 20128 29124 20164 29152
rect 20070 29112 20076 29115
rect 20128 29112 20134 29124
rect 20622 29112 20628 29164
rect 20680 29152 20686 29164
rect 22005 29155 22063 29161
rect 20680 29124 20852 29152
rect 20680 29112 20686 29124
rect 19260 29056 19932 29084
rect 20824 29084 20852 29124
rect 22005 29121 22017 29155
rect 22051 29152 22063 29155
rect 22094 29152 22100 29164
rect 22051 29124 22100 29152
rect 22051 29121 22063 29124
rect 22005 29115 22063 29121
rect 22094 29112 22100 29124
rect 22152 29112 22158 29164
rect 22189 29155 22247 29161
rect 22189 29121 22201 29155
rect 22235 29121 22247 29155
rect 22189 29115 22247 29121
rect 22465 29155 22523 29161
rect 22465 29121 22477 29155
rect 22511 29152 22523 29155
rect 22554 29152 22560 29164
rect 22511 29124 22560 29152
rect 22511 29121 22523 29124
rect 22465 29115 22523 29121
rect 22204 29084 22232 29115
rect 22554 29112 22560 29124
rect 22612 29112 22618 29164
rect 22649 29155 22707 29161
rect 22649 29121 22661 29155
rect 22695 29152 22707 29155
rect 23566 29152 23572 29164
rect 22695 29124 23572 29152
rect 22695 29121 22707 29124
rect 22649 29115 22707 29121
rect 23566 29112 23572 29124
rect 23624 29112 23630 29164
rect 24305 29155 24363 29161
rect 24305 29121 24317 29155
rect 24351 29152 24363 29155
rect 24762 29152 24768 29164
rect 24351 29124 24768 29152
rect 24351 29121 24363 29124
rect 24305 29115 24363 29121
rect 24762 29112 24768 29124
rect 24820 29152 24826 29164
rect 25317 29155 25375 29161
rect 25317 29152 25329 29155
rect 24820 29124 25329 29152
rect 24820 29112 24826 29124
rect 25317 29121 25329 29124
rect 25363 29121 25375 29155
rect 25317 29115 25375 29121
rect 25409 29155 25467 29161
rect 25409 29121 25421 29155
rect 25455 29121 25467 29155
rect 25409 29115 25467 29121
rect 22922 29084 22928 29096
rect 20824 29056 22928 29084
rect 22922 29044 22928 29056
rect 22980 29044 22986 29096
rect 24394 29084 24400 29096
rect 24355 29056 24400 29084
rect 24394 29044 24400 29056
rect 24452 29044 24458 29096
rect 24854 29044 24860 29096
rect 24912 29084 24918 29096
rect 25424 29084 25452 29115
rect 25498 29112 25504 29164
rect 25556 29152 25562 29164
rect 25593 29155 25651 29161
rect 25593 29152 25605 29155
rect 25556 29124 25605 29152
rect 25556 29112 25562 29124
rect 25593 29121 25605 29124
rect 25639 29152 25651 29155
rect 27522 29152 27528 29164
rect 25639 29124 27200 29152
rect 27483 29124 27528 29152
rect 25639 29121 25651 29124
rect 25593 29115 25651 29121
rect 25774 29084 25780 29096
rect 24912 29056 25780 29084
rect 24912 29044 24918 29056
rect 25774 29044 25780 29056
rect 25832 29044 25838 29096
rect 27172 29093 27200 29124
rect 27522 29112 27528 29124
rect 27580 29112 27586 29164
rect 28712 29155 28770 29161
rect 28712 29121 28724 29155
rect 28758 29152 28770 29155
rect 30285 29155 30343 29161
rect 30285 29152 30297 29155
rect 28758 29124 30297 29152
rect 28758 29121 28770 29124
rect 28712 29115 28770 29121
rect 30285 29121 30297 29124
rect 30331 29121 30343 29155
rect 30466 29152 30472 29164
rect 30427 29124 30472 29152
rect 30285 29115 30343 29121
rect 30466 29112 30472 29124
rect 30524 29112 30530 29164
rect 30745 29155 30803 29161
rect 30745 29121 30757 29155
rect 30791 29152 30803 29155
rect 30926 29152 30932 29164
rect 30791 29124 30932 29152
rect 30791 29121 30803 29124
rect 30745 29115 30803 29121
rect 30926 29112 30932 29124
rect 30984 29112 30990 29164
rect 31018 29112 31024 29164
rect 31076 29152 31082 29164
rect 32493 29155 32551 29161
rect 32493 29152 32505 29155
rect 31076 29124 32505 29152
rect 31076 29112 31082 29124
rect 32493 29121 32505 29124
rect 32539 29152 32551 29155
rect 32674 29152 32680 29164
rect 32539 29124 32680 29152
rect 32539 29121 32551 29124
rect 32493 29115 32551 29121
rect 32674 29112 32680 29124
rect 32732 29112 32738 29164
rect 32769 29155 32827 29161
rect 32769 29121 32781 29155
rect 32815 29121 32827 29155
rect 32769 29115 32827 29121
rect 27157 29087 27215 29093
rect 27157 29053 27169 29087
rect 27203 29053 27215 29087
rect 27157 29047 27215 29053
rect 27338 29044 27344 29096
rect 27396 29084 27402 29096
rect 27433 29087 27491 29093
rect 27433 29084 27445 29087
rect 27396 29056 27445 29084
rect 27396 29044 27402 29056
rect 27433 29053 27445 29056
rect 27479 29053 27491 29087
rect 27433 29047 27491 29053
rect 28445 29087 28503 29093
rect 28445 29053 28457 29087
rect 28491 29053 28503 29087
rect 30650 29084 30656 29096
rect 30611 29056 30656 29084
rect 28445 29047 28503 29053
rect 23750 28976 23756 29028
rect 23808 29016 23814 29028
rect 23937 29019 23995 29025
rect 23937 29016 23949 29019
rect 23808 28988 23949 29016
rect 23808 28976 23814 28988
rect 23937 28985 23949 28988
rect 23983 28985 23995 29019
rect 25590 29016 25596 29028
rect 25551 28988 25596 29016
rect 23937 28979 23995 28985
rect 25590 28976 25596 28988
rect 25648 28976 25654 29028
rect 13596 28920 15700 28948
rect 17957 28951 18015 28957
rect 13596 28908 13602 28920
rect 17957 28917 17969 28951
rect 18003 28948 18015 28951
rect 18322 28948 18328 28960
rect 18003 28920 18328 28948
rect 18003 28917 18015 28920
rect 17957 28911 18015 28917
rect 18322 28908 18328 28920
rect 18380 28948 18386 28960
rect 18598 28948 18604 28960
rect 18380 28920 18604 28948
rect 18380 28908 18386 28920
rect 18598 28908 18604 28920
rect 18656 28908 18662 28960
rect 21174 28948 21180 28960
rect 21135 28920 21180 28948
rect 21174 28908 21180 28920
rect 21232 28908 21238 28960
rect 28460 28948 28488 29047
rect 30650 29044 30656 29056
rect 30708 29044 30714 29096
rect 32784 29084 32812 29115
rect 32950 29112 32956 29164
rect 33008 29152 33014 29164
rect 33502 29152 33508 29164
rect 33008 29124 33053 29152
rect 33463 29124 33508 29152
rect 33008 29112 33014 29124
rect 33502 29112 33508 29124
rect 33560 29112 33566 29164
rect 34348 29161 34376 29192
rect 35342 29180 35348 29192
rect 35400 29180 35406 29232
rect 37274 29180 37280 29232
rect 37332 29220 37338 29232
rect 38010 29220 38016 29232
rect 37332 29192 38016 29220
rect 37332 29180 37338 29192
rect 38010 29180 38016 29192
rect 38068 29180 38074 29232
rect 40129 29223 40187 29229
rect 40129 29189 40141 29223
rect 40175 29220 40187 29223
rect 40218 29220 40224 29232
rect 40175 29192 40224 29220
rect 40175 29189 40187 29192
rect 40129 29183 40187 29189
rect 40218 29180 40224 29192
rect 40276 29180 40282 29232
rect 40678 29220 40684 29232
rect 40639 29192 40684 29220
rect 40678 29180 40684 29192
rect 40736 29180 40742 29232
rect 43530 29180 43536 29232
rect 43588 29220 43594 29232
rect 43625 29223 43683 29229
rect 43625 29220 43637 29223
rect 43588 29192 43637 29220
rect 43588 29180 43594 29192
rect 43625 29189 43637 29192
rect 43671 29189 43683 29223
rect 43625 29183 43683 29189
rect 33689 29155 33747 29161
rect 33689 29121 33701 29155
rect 33735 29121 33747 29155
rect 33689 29115 33747 29121
rect 34333 29155 34391 29161
rect 34333 29121 34345 29155
rect 34379 29121 34391 29155
rect 34589 29155 34647 29161
rect 34589 29152 34601 29155
rect 34333 29115 34391 29121
rect 34440 29124 34601 29152
rect 33226 29084 33232 29096
rect 31496 29056 33232 29084
rect 30098 28976 30104 29028
rect 30156 29016 30162 29028
rect 31496 29016 31524 29056
rect 33226 29044 33232 29056
rect 33284 29044 33290 29096
rect 33410 29084 33416 29096
rect 33371 29056 33416 29084
rect 33410 29044 33416 29056
rect 33468 29044 33474 29096
rect 30156 28988 31524 29016
rect 30156 28976 30162 28988
rect 31570 28976 31576 29028
rect 31628 29016 31634 29028
rect 33520 29016 33548 29112
rect 31628 28988 33548 29016
rect 33704 29016 33732 29115
rect 33873 29087 33931 29093
rect 33873 29053 33885 29087
rect 33919 29084 33931 29087
rect 34440 29084 34468 29124
rect 34589 29121 34601 29124
rect 34635 29121 34647 29155
rect 34589 29115 34647 29121
rect 35434 29112 35440 29164
rect 35492 29152 35498 29164
rect 36357 29155 36415 29161
rect 36357 29152 36369 29155
rect 35492 29124 36369 29152
rect 35492 29112 35498 29124
rect 36357 29121 36369 29124
rect 36403 29121 36415 29155
rect 36630 29152 36636 29164
rect 36591 29124 36636 29152
rect 36357 29115 36415 29121
rect 36630 29112 36636 29124
rect 36688 29112 36694 29164
rect 36817 29155 36875 29161
rect 36817 29121 36829 29155
rect 36863 29121 36875 29155
rect 36817 29115 36875 29121
rect 36262 29084 36268 29096
rect 33919 29056 34468 29084
rect 36175 29056 36268 29084
rect 33919 29053 33931 29056
rect 33873 29047 33931 29053
rect 36262 29044 36268 29056
rect 36320 29084 36326 29096
rect 36832 29084 36860 29115
rect 38286 29112 38292 29164
rect 38344 29152 38350 29164
rect 38381 29155 38439 29161
rect 38381 29152 38393 29155
rect 38344 29124 38393 29152
rect 38344 29112 38350 29124
rect 38381 29121 38393 29124
rect 38427 29121 38439 29155
rect 38381 29115 38439 29121
rect 38473 29155 38531 29161
rect 38473 29121 38485 29155
rect 38519 29121 38531 29155
rect 38473 29115 38531 29121
rect 38565 29155 38623 29161
rect 38565 29121 38577 29155
rect 38611 29152 38623 29155
rect 38654 29152 38660 29164
rect 38611 29124 38660 29152
rect 38611 29121 38623 29124
rect 38565 29115 38623 29121
rect 38488 29084 38516 29115
rect 38654 29112 38660 29124
rect 38712 29112 38718 29164
rect 38749 29155 38807 29161
rect 38749 29121 38761 29155
rect 38795 29121 38807 29155
rect 40586 29152 40592 29164
rect 40547 29124 40592 29152
rect 38749 29115 38807 29121
rect 36320 29056 36860 29084
rect 38304 29056 38516 29084
rect 36320 29044 36326 29056
rect 36173 29019 36231 29025
rect 36173 29016 36185 29019
rect 33704 28988 34376 29016
rect 31628 28976 31634 28988
rect 28810 28948 28816 28960
rect 28460 28920 28816 28948
rect 28810 28908 28816 28920
rect 28868 28908 28874 28960
rect 32309 28951 32367 28957
rect 32309 28917 32321 28951
rect 32355 28948 32367 28951
rect 32490 28948 32496 28960
rect 32355 28920 32496 28948
rect 32355 28917 32367 28920
rect 32309 28911 32367 28917
rect 32490 28908 32496 28920
rect 32548 28908 32554 28960
rect 34348 28948 34376 28988
rect 35268 28988 36185 29016
rect 35268 28948 35296 28988
rect 36173 28985 36185 28988
rect 36219 28985 36231 29019
rect 36173 28979 36231 28985
rect 34348 28920 35296 28948
rect 35713 28951 35771 28957
rect 35713 28917 35725 28951
rect 35759 28948 35771 28951
rect 36280 28948 36308 29044
rect 38304 29028 38332 29056
rect 37918 28976 37924 29028
rect 37976 29016 37982 29028
rect 38105 29019 38163 29025
rect 38105 29016 38117 29019
rect 37976 28988 38117 29016
rect 37976 28976 37982 28988
rect 38105 28985 38117 28988
rect 38151 28985 38163 29019
rect 38105 28979 38163 28985
rect 38286 28976 38292 29028
rect 38344 28976 38350 29028
rect 38378 28976 38384 29028
rect 38436 29016 38442 29028
rect 38764 29016 38792 29115
rect 40586 29112 40592 29124
rect 40644 29112 40650 29164
rect 40770 29152 40776 29164
rect 40731 29124 40776 29152
rect 40770 29112 40776 29124
rect 40828 29112 40834 29164
rect 42794 29112 42800 29164
rect 42852 29152 42858 29164
rect 43349 29155 43407 29161
rect 43349 29152 43361 29155
rect 42852 29124 43361 29152
rect 42852 29112 42858 29124
rect 43349 29121 43361 29124
rect 43395 29121 43407 29155
rect 43349 29115 43407 29121
rect 43714 29112 43720 29164
rect 43772 29152 43778 29164
rect 47228 29161 47256 29260
rect 47213 29155 47271 29161
rect 43772 29124 43817 29152
rect 43772 29112 43778 29124
rect 47213 29121 47225 29155
rect 47259 29152 47271 29155
rect 47302 29152 47308 29164
rect 47259 29124 47308 29152
rect 47259 29121 47271 29124
rect 47213 29115 47271 29121
rect 47302 29112 47308 29124
rect 47360 29112 47366 29164
rect 39206 29044 39212 29096
rect 39264 29084 39270 29096
rect 43162 29084 43168 29096
rect 39264 29056 43168 29084
rect 39264 29044 39270 29056
rect 43162 29044 43168 29056
rect 43220 29044 43226 29096
rect 43254 29044 43260 29096
rect 43312 29084 43318 29096
rect 43533 29087 43591 29093
rect 43533 29084 43545 29087
rect 43312 29056 43545 29084
rect 43312 29044 43318 29056
rect 43533 29053 43545 29056
rect 43579 29084 43591 29087
rect 43898 29084 43904 29096
rect 43579 29056 43904 29084
rect 43579 29053 43591 29056
rect 43533 29047 43591 29053
rect 43898 29044 43904 29056
rect 43956 29044 43962 29096
rect 38436 28988 38792 29016
rect 39853 29019 39911 29025
rect 38436 28976 38442 28988
rect 39853 28985 39865 29019
rect 39899 29016 39911 29019
rect 40218 29016 40224 29028
rect 39899 28988 40224 29016
rect 39899 28985 39911 28988
rect 39853 28979 39911 28985
rect 40218 28976 40224 28988
rect 40276 29016 40282 29028
rect 40678 29016 40684 29028
rect 40276 28988 40684 29016
rect 40276 28976 40282 28988
rect 40678 28976 40684 28988
rect 40736 28976 40742 29028
rect 43346 29016 43352 29028
rect 43307 28988 43352 29016
rect 43346 28976 43352 28988
rect 43404 28976 43410 29028
rect 44634 28976 44640 29028
rect 44692 29016 44698 29028
rect 46198 29016 46204 29028
rect 44692 28988 46204 29016
rect 44692 28976 44698 28988
rect 46198 28976 46204 28988
rect 46256 28976 46262 29028
rect 47949 29019 48007 29025
rect 47949 28985 47961 29019
rect 47995 29016 48007 29019
rect 48314 29016 48320 29028
rect 47995 28988 48320 29016
rect 47995 28985 48007 28988
rect 47949 28979 48007 28985
rect 48314 28976 48320 28988
rect 48372 28976 48378 29028
rect 35759 28920 36308 28948
rect 35759 28917 35771 28920
rect 35713 28911 35771 28917
rect 38470 28908 38476 28960
rect 38528 28948 38534 28960
rect 39114 28948 39120 28960
rect 38528 28920 39120 28948
rect 38528 28908 38534 28920
rect 39114 28908 39120 28920
rect 39172 28948 39178 28960
rect 39669 28951 39727 28957
rect 39669 28948 39681 28951
rect 39172 28920 39681 28948
rect 39172 28908 39178 28920
rect 39669 28917 39681 28920
rect 39715 28917 39727 28951
rect 39669 28911 39727 28917
rect 46474 28908 46480 28960
rect 46532 28948 46538 28960
rect 46569 28951 46627 28957
rect 46569 28948 46581 28951
rect 46532 28920 46581 28948
rect 46532 28908 46538 28920
rect 46569 28917 46581 28920
rect 46615 28917 46627 28951
rect 47118 28948 47124 28960
rect 47079 28920 47124 28948
rect 46569 28911 46627 28917
rect 47118 28908 47124 28920
rect 47176 28908 47182 28960
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 8110 28744 8116 28756
rect 8071 28716 8116 28744
rect 8110 28704 8116 28716
rect 8168 28704 8174 28756
rect 13357 28747 13415 28753
rect 13357 28713 13369 28747
rect 13403 28744 13415 28747
rect 14274 28744 14280 28756
rect 13403 28716 14280 28744
rect 13403 28713 13415 28716
rect 13357 28707 13415 28713
rect 14274 28704 14280 28716
rect 14332 28704 14338 28756
rect 16850 28744 16856 28756
rect 16811 28716 16856 28744
rect 16850 28704 16856 28716
rect 16908 28704 16914 28756
rect 17770 28744 17776 28756
rect 17236 28716 17776 28744
rect 12158 28676 12164 28688
rect 12119 28648 12164 28676
rect 12158 28636 12164 28648
rect 12216 28636 12222 28688
rect 5534 28608 5540 28620
rect 5495 28580 5540 28608
rect 5534 28568 5540 28580
rect 5592 28568 5598 28620
rect 6914 28568 6920 28620
rect 6972 28608 6978 28620
rect 6972 28580 7017 28608
rect 6972 28568 6978 28580
rect 7098 28568 7104 28620
rect 7156 28608 7162 28620
rect 7156 28580 7201 28608
rect 7156 28568 7162 28580
rect 9490 28568 9496 28620
rect 9548 28608 9554 28620
rect 9585 28611 9643 28617
rect 9585 28608 9597 28611
rect 9548 28580 9597 28608
rect 9548 28568 9554 28580
rect 9585 28577 9597 28580
rect 9631 28577 9643 28611
rect 9585 28571 9643 28577
rect 9677 28611 9735 28617
rect 9677 28577 9689 28611
rect 9723 28577 9735 28611
rect 9677 28571 9735 28577
rect 12253 28611 12311 28617
rect 12253 28577 12265 28611
rect 12299 28608 12311 28611
rect 12299 28580 12756 28608
rect 12299 28577 12311 28580
rect 12253 28571 12311 28577
rect 8018 28500 8024 28552
rect 8076 28540 8082 28552
rect 8113 28543 8171 28549
rect 8113 28540 8125 28543
rect 8076 28512 8125 28540
rect 8076 28500 8082 28512
rect 8113 28509 8125 28512
rect 8159 28509 8171 28543
rect 8113 28503 8171 28509
rect 9306 28500 9312 28552
rect 9364 28540 9370 28552
rect 9692 28540 9720 28571
rect 12728 28549 12756 28580
rect 13722 28568 13728 28620
rect 13780 28608 13786 28620
rect 14829 28611 14887 28617
rect 14829 28608 14841 28611
rect 13780 28580 14841 28608
rect 13780 28568 13786 28580
rect 14829 28577 14841 28580
rect 14875 28608 14887 28611
rect 17236 28608 17264 28716
rect 17770 28704 17776 28716
rect 17828 28704 17834 28756
rect 19426 28744 19432 28756
rect 19387 28716 19432 28744
rect 19426 28704 19432 28716
rect 19484 28704 19490 28756
rect 19797 28747 19855 28753
rect 19797 28713 19809 28747
rect 19843 28744 19855 28747
rect 20438 28744 20444 28756
rect 19843 28716 20444 28744
rect 19843 28713 19855 28716
rect 19797 28707 19855 28713
rect 20438 28704 20444 28716
rect 20496 28744 20502 28756
rect 22370 28744 22376 28756
rect 20496 28716 22376 28744
rect 20496 28704 20502 28716
rect 22370 28704 22376 28716
rect 22428 28744 22434 28756
rect 22557 28747 22615 28753
rect 22557 28744 22569 28747
rect 22428 28716 22569 28744
rect 22428 28704 22434 28716
rect 22557 28713 22569 28716
rect 22603 28713 22615 28747
rect 22557 28707 22615 28713
rect 23293 28747 23351 28753
rect 23293 28713 23305 28747
rect 23339 28744 23351 28747
rect 23474 28744 23480 28756
rect 23339 28716 23480 28744
rect 23339 28713 23351 28716
rect 23293 28707 23351 28713
rect 23474 28704 23480 28716
rect 23532 28704 23538 28756
rect 24394 28704 24400 28756
rect 24452 28744 24458 28756
rect 24673 28747 24731 28753
rect 24673 28744 24685 28747
rect 24452 28716 24685 28744
rect 24452 28704 24458 28716
rect 24673 28713 24685 28716
rect 24719 28713 24731 28747
rect 24673 28707 24731 28713
rect 31205 28747 31263 28753
rect 31205 28713 31217 28747
rect 31251 28744 31263 28747
rect 31478 28744 31484 28756
rect 31251 28716 31484 28744
rect 31251 28713 31263 28716
rect 31205 28707 31263 28713
rect 31478 28704 31484 28716
rect 31536 28704 31542 28756
rect 32214 28704 32220 28756
rect 32272 28744 32278 28756
rect 33410 28744 33416 28756
rect 32272 28716 33416 28744
rect 32272 28704 32278 28716
rect 33410 28704 33416 28716
rect 33468 28704 33474 28756
rect 35342 28744 35348 28756
rect 35084 28716 35348 28744
rect 17328 28648 22692 28676
rect 17328 28617 17356 28648
rect 14875 28580 17264 28608
rect 17313 28611 17371 28617
rect 14875 28577 14887 28580
rect 14829 28571 14887 28577
rect 17313 28577 17325 28611
rect 17359 28577 17371 28611
rect 17313 28571 17371 28577
rect 17497 28611 17555 28617
rect 17497 28577 17509 28611
rect 17543 28608 17555 28611
rect 17770 28608 17776 28620
rect 17543 28580 17776 28608
rect 17543 28577 17555 28580
rect 17497 28571 17555 28577
rect 17770 28568 17776 28580
rect 17828 28568 17834 28620
rect 19978 28608 19984 28620
rect 19628 28580 19984 28608
rect 9364 28512 9720 28540
rect 12713 28543 12771 28549
rect 9364 28500 9370 28512
rect 12713 28509 12725 28543
rect 12759 28509 12771 28543
rect 12713 28503 12771 28509
rect 12820 28512 13860 28540
rect 11793 28475 11851 28481
rect 11793 28441 11805 28475
rect 11839 28472 11851 28475
rect 11882 28472 11888 28484
rect 11839 28444 11888 28472
rect 11839 28441 11851 28444
rect 11793 28435 11851 28441
rect 11882 28432 11888 28444
rect 11940 28432 11946 28484
rect 12820 28472 12848 28512
rect 13538 28472 13544 28484
rect 12728 28444 12848 28472
rect 13499 28444 13544 28472
rect 12728 28416 12756 28444
rect 13538 28432 13544 28444
rect 13596 28432 13602 28484
rect 13725 28475 13783 28481
rect 13725 28441 13737 28475
rect 13771 28441 13783 28475
rect 13832 28472 13860 28512
rect 14642 28500 14648 28552
rect 14700 28540 14706 28552
rect 14737 28543 14795 28549
rect 14737 28540 14749 28543
rect 14700 28512 14749 28540
rect 14700 28500 14706 28512
rect 14737 28509 14749 28512
rect 14783 28509 14795 28543
rect 17218 28540 17224 28552
rect 17179 28512 17224 28540
rect 14737 28503 14795 28509
rect 17218 28500 17224 28512
rect 17276 28500 17282 28552
rect 18230 28540 18236 28552
rect 18191 28512 18236 28540
rect 18230 28500 18236 28512
rect 18288 28500 18294 28552
rect 18322 28500 18328 28552
rect 18380 28540 18386 28552
rect 18598 28540 18604 28552
rect 18380 28512 18425 28540
rect 18559 28512 18604 28540
rect 18380 28500 18386 28512
rect 18598 28500 18604 28512
rect 18656 28500 18662 28552
rect 19628 28549 19656 28580
rect 19978 28568 19984 28580
rect 20036 28568 20042 28620
rect 20898 28568 20904 28620
rect 20956 28608 20962 28620
rect 22554 28608 22560 28620
rect 20956 28580 22560 28608
rect 20956 28568 20962 28580
rect 22554 28568 22560 28580
rect 22612 28568 22618 28620
rect 19613 28543 19671 28549
rect 19613 28509 19625 28543
rect 19659 28509 19671 28543
rect 19613 28503 19671 28509
rect 19889 28543 19947 28549
rect 19889 28509 19901 28543
rect 19935 28509 19947 28543
rect 19889 28503 19947 28509
rect 20533 28543 20591 28549
rect 20533 28509 20545 28543
rect 20579 28540 20591 28543
rect 20622 28540 20628 28552
rect 20579 28512 20628 28540
rect 20579 28509 20591 28512
rect 20533 28503 20591 28509
rect 18414 28472 18420 28484
rect 13832 28444 14688 28472
rect 18375 28444 18420 28472
rect 13725 28435 13783 28441
rect 9122 28404 9128 28416
rect 9083 28376 9128 28404
rect 9122 28364 9128 28376
rect 9180 28364 9186 28416
rect 9493 28407 9551 28413
rect 9493 28373 9505 28407
rect 9539 28404 9551 28407
rect 12710 28404 12716 28416
rect 9539 28376 12716 28404
rect 9539 28373 9551 28376
rect 9493 28367 9551 28373
rect 12710 28364 12716 28376
rect 12768 28364 12774 28416
rect 12894 28404 12900 28416
rect 12855 28376 12900 28404
rect 12894 28364 12900 28376
rect 12952 28364 12958 28416
rect 13740 28404 13768 28435
rect 14660 28413 14688 28444
rect 18414 28432 18420 28444
rect 18472 28432 18478 28484
rect 19426 28432 19432 28484
rect 19484 28472 19490 28484
rect 19904 28472 19932 28503
rect 20622 28500 20628 28512
rect 20680 28500 20686 28552
rect 20809 28543 20867 28549
rect 20809 28509 20821 28543
rect 20855 28540 20867 28543
rect 20916 28540 20944 28568
rect 22664 28552 22692 28648
rect 23750 28608 23756 28620
rect 23711 28580 23756 28608
rect 23750 28568 23756 28580
rect 23808 28568 23814 28620
rect 23845 28611 23903 28617
rect 23845 28577 23857 28611
rect 23891 28577 23903 28611
rect 25866 28608 25872 28620
rect 23845 28571 23903 28577
rect 24596 28580 25872 28608
rect 20855 28512 20944 28540
rect 20993 28543 21051 28549
rect 20855 28509 20867 28512
rect 20809 28503 20867 28509
rect 20993 28509 21005 28543
rect 21039 28540 21051 28543
rect 21174 28540 21180 28552
rect 21039 28512 21180 28540
rect 21039 28509 21051 28512
rect 20993 28503 21051 28509
rect 21174 28500 21180 28512
rect 21232 28500 21238 28552
rect 22370 28540 22376 28552
rect 22331 28512 22376 28540
rect 22370 28500 22376 28512
rect 22428 28500 22434 28552
rect 22646 28540 22652 28552
rect 22607 28512 22652 28540
rect 22646 28500 22652 28512
rect 22704 28500 22710 28552
rect 23566 28500 23572 28552
rect 23624 28540 23630 28552
rect 23860 28540 23888 28571
rect 23624 28512 23888 28540
rect 23624 28500 23630 28512
rect 24118 28500 24124 28552
rect 24176 28540 24182 28552
rect 24596 28549 24624 28580
rect 25866 28568 25872 28580
rect 25924 28568 25930 28620
rect 29086 28568 29092 28620
rect 29144 28608 29150 28620
rect 30101 28611 30159 28617
rect 29144 28580 30052 28608
rect 29144 28568 29150 28580
rect 24581 28543 24639 28549
rect 24581 28540 24593 28543
rect 24176 28512 24593 28540
rect 24176 28500 24182 28512
rect 24581 28509 24593 28512
rect 24627 28509 24639 28543
rect 24581 28503 24639 28509
rect 24765 28543 24823 28549
rect 24765 28509 24777 28543
rect 24811 28540 24823 28543
rect 24854 28540 24860 28552
rect 24811 28512 24860 28540
rect 24811 28509 24823 28512
rect 24765 28503 24823 28509
rect 24854 28500 24860 28512
rect 24912 28500 24918 28552
rect 29914 28540 29920 28552
rect 29875 28512 29920 28540
rect 29914 28500 29920 28512
rect 29972 28500 29978 28552
rect 30024 28540 30052 28580
rect 30101 28577 30113 28611
rect 30147 28608 30159 28611
rect 30650 28608 30656 28620
rect 30147 28580 30656 28608
rect 30147 28577 30159 28580
rect 30101 28571 30159 28577
rect 30650 28568 30656 28580
rect 30708 28608 30714 28620
rect 31570 28608 31576 28620
rect 30708 28580 31576 28608
rect 30708 28568 30714 28580
rect 31570 28568 31576 28580
rect 31628 28568 31634 28620
rect 35084 28617 35112 28716
rect 35342 28704 35348 28716
rect 35400 28704 35406 28756
rect 36446 28744 36452 28756
rect 36407 28716 36452 28744
rect 36446 28704 36452 28716
rect 36504 28704 36510 28756
rect 38286 28744 38292 28756
rect 38247 28716 38292 28744
rect 38286 28704 38292 28716
rect 38344 28704 38350 28756
rect 38654 28704 38660 28756
rect 38712 28744 38718 28756
rect 39301 28747 39359 28753
rect 39301 28744 39313 28747
rect 38712 28716 39313 28744
rect 38712 28704 38718 28716
rect 39301 28713 39313 28716
rect 39347 28713 39359 28747
rect 39301 28707 39359 28713
rect 37182 28636 37188 28688
rect 37240 28676 37246 28688
rect 40310 28676 40316 28688
rect 37240 28648 37412 28676
rect 40271 28648 40316 28676
rect 37240 28636 37246 28648
rect 32585 28611 32643 28617
rect 32585 28577 32597 28611
rect 32631 28608 32643 28611
rect 35069 28611 35127 28617
rect 35069 28608 35081 28611
rect 32631 28580 35081 28608
rect 32631 28577 32643 28580
rect 32585 28571 32643 28577
rect 35069 28577 35081 28580
rect 35115 28577 35127 28611
rect 35069 28571 35127 28577
rect 37384 28552 37412 28648
rect 40310 28636 40316 28648
rect 40368 28636 40374 28688
rect 40126 28608 40132 28620
rect 38580 28580 39160 28608
rect 30193 28543 30251 28549
rect 30193 28540 30205 28543
rect 30024 28512 30205 28540
rect 30193 28509 30205 28512
rect 30239 28509 30251 28543
rect 30193 28503 30251 28509
rect 31478 28500 31484 28552
rect 31536 28540 31542 28552
rect 33042 28540 33048 28552
rect 31536 28512 32444 28540
rect 33003 28512 33048 28540
rect 31536 28500 31542 28512
rect 32214 28472 32220 28484
rect 19484 28444 32220 28472
rect 19484 28432 19490 28444
rect 32214 28432 32220 28444
rect 32272 28432 32278 28484
rect 32318 28475 32376 28481
rect 32318 28441 32330 28475
rect 32364 28441 32376 28475
rect 32416 28472 32444 28512
rect 33042 28500 33048 28512
rect 33100 28500 33106 28552
rect 33138 28543 33196 28549
rect 33138 28509 33150 28543
rect 33184 28509 33196 28543
rect 33138 28503 33196 28509
rect 33152 28472 33180 28503
rect 33226 28500 33232 28552
rect 33284 28540 33290 28552
rect 33510 28543 33568 28549
rect 33510 28540 33522 28543
rect 33284 28512 33522 28540
rect 33284 28500 33290 28512
rect 33510 28509 33522 28512
rect 33556 28509 33568 28543
rect 33510 28503 33568 28509
rect 37185 28543 37243 28549
rect 37185 28509 37197 28543
rect 37231 28509 37243 28543
rect 37366 28540 37372 28552
rect 37327 28512 37372 28540
rect 37185 28503 37243 28509
rect 33318 28472 33324 28484
rect 32416 28444 33180 28472
rect 33279 28444 33324 28472
rect 32318 28435 32376 28441
rect 14277 28407 14335 28413
rect 14277 28404 14289 28407
rect 13740 28376 14289 28404
rect 14277 28373 14289 28376
rect 14323 28373 14335 28407
rect 14277 28367 14335 28373
rect 14645 28407 14703 28413
rect 14645 28373 14657 28407
rect 14691 28373 14703 28407
rect 18046 28404 18052 28416
rect 18007 28376 18052 28404
rect 14645 28367 14703 28373
rect 18046 28364 18052 28376
rect 18104 28364 18110 28416
rect 20254 28364 20260 28416
rect 20312 28404 20318 28416
rect 20349 28407 20407 28413
rect 20349 28404 20361 28407
rect 20312 28376 20361 28404
rect 20312 28364 20318 28376
rect 20349 28373 20361 28376
rect 20395 28373 20407 28407
rect 20349 28367 20407 28373
rect 22189 28407 22247 28413
rect 22189 28373 22201 28407
rect 22235 28404 22247 28407
rect 22278 28404 22284 28416
rect 22235 28376 22284 28404
rect 22235 28373 22247 28376
rect 22189 28367 22247 28373
rect 22278 28364 22284 28376
rect 22336 28364 22342 28416
rect 23382 28364 23388 28416
rect 23440 28404 23446 28416
rect 23661 28407 23719 28413
rect 23661 28404 23673 28407
rect 23440 28376 23673 28404
rect 23440 28364 23446 28376
rect 23661 28373 23673 28376
rect 23707 28373 23719 28407
rect 29730 28404 29736 28416
rect 29691 28376 29736 28404
rect 23661 28367 23719 28373
rect 29730 28364 29736 28376
rect 29788 28364 29794 28416
rect 32324 28404 32352 28435
rect 33318 28432 33324 28444
rect 33376 28432 33382 28484
rect 33410 28432 33416 28484
rect 33468 28472 33474 28484
rect 33468 28444 33513 28472
rect 33468 28432 33474 28444
rect 34974 28432 34980 28484
rect 35032 28472 35038 28484
rect 35314 28475 35372 28481
rect 35314 28472 35326 28475
rect 35032 28444 35326 28472
rect 35032 28432 35038 28444
rect 35314 28441 35326 28444
rect 35360 28441 35372 28475
rect 37200 28472 37228 28503
rect 37366 28500 37372 28512
rect 37424 28500 37430 28552
rect 38470 28540 38476 28552
rect 38528 28549 38534 28552
rect 38580 28549 38608 28580
rect 39132 28552 39160 28580
rect 39408 28580 40132 28608
rect 38435 28512 38476 28540
rect 38470 28500 38476 28512
rect 38528 28503 38535 28549
rect 38565 28543 38623 28549
rect 38565 28509 38577 28543
rect 38611 28509 38623 28543
rect 38657 28543 38715 28549
rect 38657 28530 38669 28543
rect 38703 28530 38715 28543
rect 38565 28503 38623 28509
rect 38528 28500 38534 28503
rect 37458 28472 37464 28484
rect 37200 28444 37464 28472
rect 35314 28435 35372 28441
rect 37458 28432 37464 28444
rect 37516 28432 37522 28484
rect 38654 28478 38660 28530
rect 38712 28478 38718 28530
rect 39114 28500 39120 28552
rect 39172 28540 39178 28552
rect 39408 28549 39436 28580
rect 40126 28568 40132 28580
rect 40184 28568 40190 28620
rect 42058 28568 42064 28620
rect 42116 28608 42122 28620
rect 42429 28611 42487 28617
rect 42429 28608 42441 28611
rect 42116 28580 42441 28608
rect 42116 28568 42122 28580
rect 42429 28577 42441 28580
rect 42475 28577 42487 28611
rect 42429 28571 42487 28577
rect 42521 28611 42579 28617
rect 42521 28577 42533 28611
rect 42567 28608 42579 28611
rect 43346 28608 43352 28620
rect 42567 28580 43352 28608
rect 42567 28577 42579 28580
rect 42521 28571 42579 28577
rect 43346 28568 43352 28580
rect 43404 28568 43410 28620
rect 46474 28608 46480 28620
rect 46435 28580 46480 28608
rect 46474 28568 46480 28580
rect 46532 28568 46538 28620
rect 46661 28611 46719 28617
rect 46661 28577 46673 28611
rect 46707 28608 46719 28611
rect 47118 28608 47124 28620
rect 46707 28580 47124 28608
rect 46707 28577 46719 28580
rect 46661 28571 46719 28577
rect 47118 28568 47124 28580
rect 47176 28568 47182 28620
rect 48222 28608 48228 28620
rect 48183 28580 48228 28608
rect 48222 28568 48228 28580
rect 48280 28568 48286 28620
rect 39209 28543 39267 28549
rect 39209 28540 39221 28543
rect 39172 28512 39221 28540
rect 39172 28500 39178 28512
rect 39209 28509 39221 28512
rect 39255 28509 39267 28543
rect 39209 28503 39267 28509
rect 39393 28543 39451 28549
rect 39393 28509 39405 28543
rect 39439 28509 39451 28543
rect 39393 28503 39451 28509
rect 40037 28543 40095 28549
rect 40037 28509 40049 28543
rect 40083 28540 40095 28543
rect 40218 28540 40224 28552
rect 40083 28512 40224 28540
rect 40083 28509 40095 28512
rect 40037 28503 40095 28509
rect 40218 28500 40224 28512
rect 40276 28500 40282 28552
rect 40313 28543 40371 28549
rect 40313 28509 40325 28543
rect 40359 28540 40371 28543
rect 40402 28540 40408 28552
rect 40359 28512 40408 28540
rect 40359 28509 40371 28512
rect 40313 28503 40371 28509
rect 40402 28500 40408 28512
rect 40460 28500 40466 28552
rect 42337 28543 42395 28549
rect 42337 28509 42349 28543
rect 42383 28509 42395 28543
rect 42337 28503 42395 28509
rect 42613 28543 42671 28549
rect 42613 28509 42625 28543
rect 42659 28540 42671 28543
rect 42794 28540 42800 28552
rect 42659 28512 42800 28540
rect 42659 28509 42671 28512
rect 42613 28503 42671 28509
rect 40129 28475 40187 28481
rect 40129 28441 40141 28475
rect 40175 28472 40187 28475
rect 40494 28472 40500 28484
rect 40175 28444 40500 28472
rect 40175 28441 40187 28444
rect 40129 28435 40187 28441
rect 40494 28432 40500 28444
rect 40552 28432 40558 28484
rect 42352 28472 42380 28503
rect 42794 28500 42800 28512
rect 42852 28500 42858 28552
rect 43625 28543 43683 28549
rect 43625 28509 43637 28543
rect 43671 28540 43683 28543
rect 43714 28540 43720 28552
rect 43671 28512 43720 28540
rect 43671 28509 43683 28512
rect 43625 28503 43683 28509
rect 43714 28500 43720 28512
rect 43772 28500 43778 28552
rect 43898 28540 43904 28552
rect 43859 28512 43904 28540
rect 43898 28500 43904 28512
rect 43956 28500 43962 28552
rect 43806 28472 43812 28484
rect 42352 28444 43812 28472
rect 43806 28432 43812 28444
rect 43864 28432 43870 28484
rect 33689 28407 33747 28413
rect 33689 28404 33701 28407
rect 32324 28376 33701 28404
rect 33689 28373 33701 28376
rect 33735 28373 33747 28407
rect 37550 28404 37556 28416
rect 37511 28376 37556 28404
rect 33689 28367 33747 28373
rect 37550 28364 37556 28376
rect 37608 28364 37614 28416
rect 41782 28364 41788 28416
rect 41840 28404 41846 28416
rect 42153 28407 42211 28413
rect 42153 28404 42165 28407
rect 41840 28376 42165 28404
rect 41840 28364 41846 28376
rect 42153 28373 42165 28376
rect 42199 28373 42211 28407
rect 42153 28367 42211 28373
rect 43530 28364 43536 28416
rect 43588 28404 43594 28416
rect 43717 28407 43775 28413
rect 43717 28404 43729 28407
rect 43588 28376 43729 28404
rect 43588 28364 43594 28376
rect 43717 28373 43729 28376
rect 43763 28373 43775 28407
rect 43717 28367 43775 28373
rect 43990 28364 43996 28416
rect 44048 28404 44054 28416
rect 44085 28407 44143 28413
rect 44085 28404 44097 28407
rect 44048 28376 44097 28404
rect 44048 28364 44054 28376
rect 44085 28373 44097 28376
rect 44131 28373 44143 28407
rect 44085 28367 44143 28373
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 11057 28203 11115 28209
rect 11057 28169 11069 28203
rect 11103 28200 11115 28203
rect 12618 28200 12624 28212
rect 11103 28172 12624 28200
rect 11103 28169 11115 28172
rect 11057 28163 11115 28169
rect 12618 28160 12624 28172
rect 12676 28160 12682 28212
rect 17126 28160 17132 28212
rect 17184 28200 17190 28212
rect 18233 28203 18291 28209
rect 18233 28200 18245 28203
rect 17184 28172 18245 28200
rect 17184 28160 17190 28172
rect 18233 28169 18245 28172
rect 18279 28200 18291 28203
rect 18598 28200 18604 28212
rect 18279 28172 18604 28200
rect 18279 28169 18291 28172
rect 18233 28163 18291 28169
rect 18598 28160 18604 28172
rect 18656 28160 18662 28212
rect 20070 28200 20076 28212
rect 20031 28172 20076 28200
rect 20070 28160 20076 28172
rect 20128 28160 20134 28212
rect 23382 28200 23388 28212
rect 23343 28172 23388 28200
rect 23382 28160 23388 28172
rect 23440 28160 23446 28212
rect 30193 28203 30251 28209
rect 30193 28169 30205 28203
rect 30239 28200 30251 28203
rect 30374 28200 30380 28212
rect 30239 28172 30380 28200
rect 30239 28169 30251 28172
rect 30193 28163 30251 28169
rect 30374 28160 30380 28172
rect 30432 28200 30438 28212
rect 33410 28200 33416 28212
rect 30432 28172 33416 28200
rect 30432 28160 30438 28172
rect 33410 28160 33416 28172
rect 33468 28160 33474 28212
rect 34974 28200 34980 28212
rect 34935 28172 34980 28200
rect 34974 28160 34980 28172
rect 35032 28160 35038 28212
rect 42794 28200 42800 28212
rect 42755 28172 42800 28200
rect 42794 28160 42800 28172
rect 42852 28160 42858 28212
rect 43162 28200 43168 28212
rect 43123 28172 43168 28200
rect 43162 28160 43168 28172
rect 43220 28160 43226 28212
rect 43806 28160 43812 28212
rect 43864 28200 43870 28212
rect 43993 28203 44051 28209
rect 43993 28200 44005 28203
rect 43864 28172 44005 28200
rect 43864 28160 43870 28172
rect 43993 28169 44005 28172
rect 44039 28169 44051 28203
rect 43993 28163 44051 28169
rect 12894 28092 12900 28144
rect 12952 28141 12958 28144
rect 12952 28132 12964 28141
rect 12952 28104 12997 28132
rect 12952 28095 12964 28104
rect 12952 28092 12958 28095
rect 18414 28092 18420 28144
rect 18472 28132 18478 28144
rect 18472 28104 22416 28132
rect 18472 28092 18478 28104
rect 6733 28067 6791 28073
rect 6733 28033 6745 28067
rect 6779 28064 6791 28067
rect 7190 28064 7196 28076
rect 6779 28036 7196 28064
rect 6779 28033 6791 28036
rect 6733 28027 6791 28033
rect 7190 28024 7196 28036
rect 7248 28024 7254 28076
rect 9122 28064 9128 28076
rect 9083 28036 9128 28064
rect 9122 28024 9128 28036
rect 9180 28024 9186 28076
rect 9214 28024 9220 28076
rect 9272 28064 9278 28076
rect 10689 28067 10747 28073
rect 10689 28064 10701 28067
rect 9272 28036 10701 28064
rect 9272 28024 9278 28036
rect 10689 28033 10701 28036
rect 10735 28033 10747 28067
rect 10689 28027 10747 28033
rect 13173 28067 13231 28073
rect 13173 28033 13185 28067
rect 13219 28064 13231 28067
rect 14734 28064 14740 28076
rect 13219 28036 14740 28064
rect 13219 28033 13231 28036
rect 13173 28027 13231 28033
rect 14734 28024 14740 28036
rect 14792 28064 14798 28076
rect 16853 28067 16911 28073
rect 16853 28064 16865 28067
rect 14792 28036 16865 28064
rect 14792 28024 14798 28036
rect 16853 28033 16865 28036
rect 16899 28033 16911 28067
rect 16853 28027 16911 28033
rect 17120 28067 17178 28073
rect 17120 28033 17132 28067
rect 17166 28064 17178 28067
rect 17402 28064 17408 28076
rect 17166 28036 17408 28064
rect 17166 28033 17178 28036
rect 17120 28027 17178 28033
rect 17402 28024 17408 28036
rect 17460 28024 17466 28076
rect 20254 28064 20260 28076
rect 20215 28036 20260 28064
rect 20254 28024 20260 28036
rect 20312 28024 20318 28076
rect 20438 28064 20444 28076
rect 20399 28036 20444 28064
rect 20438 28024 20444 28036
rect 20496 28024 20502 28076
rect 22278 28073 22284 28076
rect 22272 28064 22284 28073
rect 22239 28036 22284 28064
rect 22272 28027 22284 28036
rect 22278 28024 22284 28027
rect 22336 28024 22342 28076
rect 22388 28064 22416 28104
rect 22646 28092 22652 28144
rect 22704 28132 22710 28144
rect 29080 28135 29138 28141
rect 22704 28104 27936 28132
rect 22704 28092 22710 28104
rect 25038 28064 25044 28076
rect 22388 28036 25044 28064
rect 25038 28024 25044 28036
rect 25096 28024 25102 28076
rect 25406 28064 25412 28076
rect 25367 28036 25412 28064
rect 25406 28024 25412 28036
rect 25464 28024 25470 28076
rect 25700 28073 25728 28104
rect 25685 28067 25743 28073
rect 25685 28033 25697 28067
rect 25731 28033 25743 28067
rect 25685 28027 25743 28033
rect 27341 28067 27399 28073
rect 27341 28033 27353 28067
rect 27387 28064 27399 28067
rect 27798 28064 27804 28076
rect 27387 28036 27804 28064
rect 27387 28033 27399 28036
rect 27341 28027 27399 28033
rect 27798 28024 27804 28036
rect 27856 28024 27862 28076
rect 27908 28064 27936 28104
rect 29080 28101 29092 28135
rect 29126 28132 29138 28135
rect 29730 28132 29736 28144
rect 29126 28104 29736 28132
rect 29126 28101 29138 28104
rect 29080 28095 29138 28101
rect 29730 28092 29736 28104
rect 29788 28092 29794 28144
rect 37550 28092 37556 28144
rect 37608 28132 37614 28144
rect 38289 28135 38347 28141
rect 38289 28132 38301 28135
rect 37608 28104 38301 28132
rect 37608 28092 37614 28104
rect 38289 28101 38301 28104
rect 38335 28101 38347 28135
rect 38289 28095 38347 28101
rect 38473 28135 38531 28141
rect 38473 28101 38485 28135
rect 38519 28132 38531 28135
rect 39206 28132 39212 28144
rect 38519 28104 39212 28132
rect 38519 28101 38531 28104
rect 38473 28095 38531 28101
rect 39206 28092 39212 28104
rect 39264 28092 39270 28144
rect 40034 28092 40040 28144
rect 40092 28132 40098 28144
rect 40678 28132 40684 28144
rect 40092 28104 40684 28132
rect 40092 28092 40098 28104
rect 40678 28092 40684 28104
rect 40736 28092 40742 28144
rect 42996 28104 43944 28132
rect 30926 28064 30932 28076
rect 27908 28036 30932 28064
rect 30926 28024 30932 28036
rect 30984 28024 30990 28076
rect 34698 28024 34704 28076
rect 34756 28064 34762 28076
rect 34793 28067 34851 28073
rect 34793 28064 34805 28067
rect 34756 28036 34805 28064
rect 34756 28024 34762 28036
rect 34793 28033 34805 28036
rect 34839 28033 34851 28067
rect 34793 28027 34851 28033
rect 39945 28067 40003 28073
rect 39945 28033 39957 28067
rect 39991 28064 40003 28067
rect 40126 28064 40132 28076
rect 39991 28036 40132 28064
rect 39991 28033 40003 28036
rect 39945 28027 40003 28033
rect 40126 28024 40132 28036
rect 40184 28024 40190 28076
rect 41877 28067 41935 28073
rect 41877 28033 41889 28067
rect 41923 28064 41935 28067
rect 42058 28064 42064 28076
rect 41923 28036 42064 28064
rect 41923 28033 41935 28036
rect 41877 28027 41935 28033
rect 42058 28024 42064 28036
rect 42116 28024 42122 28076
rect 6825 27999 6883 28005
rect 6825 27965 6837 27999
rect 6871 27965 6883 27999
rect 6825 27959 6883 27965
rect 6840 27928 6868 27959
rect 7006 27956 7012 28008
rect 7064 27996 7070 28008
rect 7101 27999 7159 28005
rect 7101 27996 7113 27999
rect 7064 27968 7113 27996
rect 7064 27956 7070 27968
rect 7101 27965 7113 27968
rect 7147 27965 7159 27999
rect 10594 27996 10600 28008
rect 10555 27968 10600 27996
rect 7101 27959 7159 27965
rect 10594 27956 10600 27968
rect 10652 27956 10658 28008
rect 20346 27956 20352 28008
rect 20404 27996 20410 28008
rect 20533 27999 20591 28005
rect 20533 27996 20545 27999
rect 20404 27968 20545 27996
rect 20404 27956 20410 27968
rect 20533 27965 20545 27968
rect 20579 27965 20591 27999
rect 22002 27996 22008 28008
rect 21963 27968 22008 27996
rect 20533 27959 20591 27965
rect 8202 27928 8208 27940
rect 6840 27900 8208 27928
rect 8202 27888 8208 27900
rect 8260 27888 8266 27940
rect 8941 27863 8999 27869
rect 8941 27829 8953 27863
rect 8987 27860 8999 27863
rect 9030 27860 9036 27872
rect 8987 27832 9036 27860
rect 8987 27829 8999 27832
rect 8941 27823 8999 27829
rect 9030 27820 9036 27832
rect 9088 27820 9094 27872
rect 11790 27860 11796 27872
rect 11751 27832 11796 27860
rect 11790 27820 11796 27832
rect 11848 27820 11854 27872
rect 20548 27860 20576 27959
rect 22002 27956 22008 27968
rect 22060 27956 22066 28008
rect 27614 27996 27620 28008
rect 27575 27968 27620 27996
rect 27614 27956 27620 27968
rect 27672 27956 27678 28008
rect 28810 27996 28816 28008
rect 28771 27968 28816 27996
rect 28810 27956 28816 27968
rect 28868 27956 28874 28008
rect 34514 27996 34520 28008
rect 34427 27968 34520 27996
rect 34514 27956 34520 27968
rect 34572 27996 34578 28008
rect 39850 27996 39856 28008
rect 34572 27968 39856 27996
rect 34572 27956 34578 27968
rect 39850 27956 39856 27968
rect 39908 27956 39914 28008
rect 41601 27999 41659 28005
rect 41601 27965 41613 27999
rect 41647 27996 41659 27999
rect 41647 27968 42748 27996
rect 41647 27965 41659 27968
rect 41601 27959 41659 27965
rect 25593 27931 25651 27937
rect 25593 27897 25605 27931
rect 25639 27928 25651 27931
rect 26234 27928 26240 27940
rect 25639 27900 26240 27928
rect 25639 27897 25651 27900
rect 25593 27891 25651 27897
rect 26234 27888 26240 27900
rect 26292 27928 26298 27940
rect 27525 27931 27583 27937
rect 27525 27928 27537 27931
rect 26292 27900 27537 27928
rect 26292 27888 26298 27900
rect 27525 27897 27537 27900
rect 27571 27897 27583 27931
rect 27525 27891 27583 27897
rect 31662 27888 31668 27940
rect 31720 27928 31726 27940
rect 34609 27931 34667 27937
rect 34609 27928 34621 27931
rect 31720 27900 34621 27928
rect 31720 27888 31726 27900
rect 34609 27897 34621 27900
rect 34655 27897 34667 27931
rect 34609 27891 34667 27897
rect 37090 27888 37096 27940
rect 37148 27928 37154 27940
rect 37458 27928 37464 27940
rect 37148 27900 37464 27928
rect 37148 27888 37154 27900
rect 37458 27888 37464 27900
rect 37516 27928 37522 27940
rect 41414 27928 41420 27940
rect 37516 27900 41420 27928
rect 37516 27888 37522 27900
rect 41414 27888 41420 27900
rect 41472 27928 41478 27940
rect 42720 27928 42748 27968
rect 42794 27956 42800 28008
rect 42852 27996 42858 28008
rect 42996 28005 43024 28104
rect 43073 28067 43131 28073
rect 43073 28033 43085 28067
rect 43119 28064 43131 28067
rect 43254 28064 43260 28076
rect 43119 28036 43260 28064
rect 43119 28033 43131 28036
rect 43073 28027 43131 28033
rect 43254 28024 43260 28036
rect 43312 28024 43318 28076
rect 43441 28067 43499 28073
rect 43441 28033 43453 28067
rect 43487 28064 43499 28067
rect 43714 28064 43720 28076
rect 43487 28036 43720 28064
rect 43487 28033 43499 28036
rect 43441 28027 43499 28033
rect 43714 28024 43720 28036
rect 43772 28024 43778 28076
rect 43916 28073 43944 28104
rect 43901 28067 43959 28073
rect 43901 28033 43913 28067
rect 43947 28033 43959 28067
rect 43901 28027 43959 28033
rect 44082 28024 44088 28076
rect 44140 28064 44146 28076
rect 44637 28067 44695 28073
rect 44637 28064 44649 28067
rect 44140 28036 44649 28064
rect 44140 28024 44146 28036
rect 44637 28033 44649 28036
rect 44683 28033 44695 28067
rect 44637 28027 44695 28033
rect 44726 28024 44732 28076
rect 44784 28064 44790 28076
rect 44893 28067 44951 28073
rect 44893 28064 44905 28067
rect 44784 28036 44905 28064
rect 44784 28024 44790 28036
rect 44893 28033 44905 28036
rect 44939 28033 44951 28067
rect 47762 28064 47768 28076
rect 47723 28036 47768 28064
rect 44893 28027 44951 28033
rect 47762 28024 47768 28036
rect 47820 28024 47826 28076
rect 42981 27999 43039 28005
rect 42981 27996 42993 27999
rect 42852 27968 42993 27996
rect 42852 27956 42858 27968
rect 42981 27965 42993 27968
rect 43027 27965 43039 27999
rect 42981 27959 43039 27965
rect 43349 27999 43407 28005
rect 43349 27965 43361 27999
rect 43395 27996 43407 27999
rect 43530 27996 43536 28008
rect 43395 27968 43536 27996
rect 43395 27965 43407 27968
rect 43349 27959 43407 27965
rect 43530 27956 43536 27968
rect 43588 27956 43594 28008
rect 44358 27928 44364 27940
rect 41472 27900 42288 27928
rect 42720 27900 44364 27928
rect 41472 27888 41478 27900
rect 23934 27860 23940 27872
rect 20548 27832 23940 27860
rect 23934 27820 23940 27832
rect 23992 27820 23998 27872
rect 25222 27860 25228 27872
rect 25183 27832 25228 27860
rect 25222 27820 25228 27832
rect 25280 27820 25286 27872
rect 27154 27860 27160 27872
rect 27115 27832 27160 27860
rect 27154 27820 27160 27832
rect 27212 27820 27218 27872
rect 33318 27820 33324 27872
rect 33376 27860 33382 27872
rect 39022 27860 39028 27872
rect 33376 27832 39028 27860
rect 33376 27820 33382 27832
rect 39022 27820 39028 27832
rect 39080 27860 39086 27872
rect 42058 27860 42064 27872
rect 39080 27832 42064 27860
rect 39080 27820 39086 27832
rect 42058 27820 42064 27832
rect 42116 27820 42122 27872
rect 42260 27860 42288 27900
rect 44358 27888 44364 27900
rect 44416 27888 44422 27940
rect 42978 27860 42984 27872
rect 42260 27832 42984 27860
rect 42978 27820 42984 27832
rect 43036 27820 43042 27872
rect 43898 27820 43904 27872
rect 43956 27860 43962 27872
rect 46017 27863 46075 27869
rect 46017 27860 46029 27863
rect 43956 27832 46029 27860
rect 43956 27820 43962 27832
rect 46017 27829 46029 27832
rect 46063 27860 46075 27863
rect 46474 27860 46480 27872
rect 46063 27832 46480 27860
rect 46063 27829 46075 27832
rect 46017 27823 46075 27829
rect 46474 27820 46480 27832
rect 46532 27820 46538 27872
rect 47857 27863 47915 27869
rect 47857 27829 47869 27863
rect 47903 27860 47915 27863
rect 48130 27860 48136 27872
rect 47903 27832 48136 27860
rect 47903 27829 47915 27832
rect 47857 27823 47915 27829
rect 48130 27820 48136 27832
rect 48188 27820 48194 27872
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 12158 27656 12164 27668
rect 12119 27628 12164 27656
rect 12158 27616 12164 27628
rect 12216 27616 12222 27668
rect 17402 27656 17408 27668
rect 17363 27628 17408 27656
rect 17402 27616 17408 27628
rect 17460 27616 17466 27668
rect 17512 27628 17724 27656
rect 7190 27588 7196 27600
rect 7151 27560 7196 27588
rect 7190 27548 7196 27560
rect 7248 27548 7254 27600
rect 8205 27591 8263 27597
rect 8205 27557 8217 27591
rect 8251 27588 8263 27591
rect 9214 27588 9220 27600
rect 8251 27560 9220 27588
rect 8251 27557 8263 27560
rect 8205 27551 8263 27557
rect 9214 27548 9220 27560
rect 9272 27548 9278 27600
rect 10594 27588 10600 27600
rect 10555 27560 10600 27588
rect 10594 27548 10600 27560
rect 10652 27548 10658 27600
rect 14826 27548 14832 27600
rect 14884 27588 14890 27600
rect 17512 27588 17540 27628
rect 14884 27560 17540 27588
rect 14884 27548 14890 27560
rect 17586 27548 17592 27600
rect 17644 27548 17650 27600
rect 17696 27588 17724 27628
rect 22370 27616 22376 27668
rect 22428 27656 22434 27668
rect 22649 27659 22707 27665
rect 22649 27656 22661 27659
rect 22428 27628 22661 27656
rect 22428 27616 22434 27628
rect 22649 27625 22661 27628
rect 22695 27625 22707 27659
rect 22649 27619 22707 27625
rect 25774 27616 25780 27668
rect 25832 27616 25838 27668
rect 29733 27659 29791 27665
rect 29733 27625 29745 27659
rect 29779 27656 29791 27659
rect 29914 27656 29920 27668
rect 29779 27628 29920 27656
rect 29779 27625 29791 27628
rect 29733 27619 29791 27625
rect 29914 27616 29920 27628
rect 29972 27616 29978 27668
rect 38378 27656 38384 27668
rect 38339 27628 38384 27656
rect 38378 27616 38384 27628
rect 38436 27616 38442 27668
rect 38565 27659 38623 27665
rect 38565 27625 38577 27659
rect 38611 27656 38623 27659
rect 39114 27656 39120 27668
rect 38611 27628 39120 27656
rect 38611 27625 38623 27628
rect 38565 27619 38623 27625
rect 39114 27616 39120 27628
rect 39172 27616 39178 27668
rect 40678 27616 40684 27668
rect 40736 27656 40742 27668
rect 40736 27628 41414 27656
rect 40736 27616 40742 27628
rect 19426 27588 19432 27600
rect 17696 27560 19432 27588
rect 19426 27548 19432 27560
rect 19484 27548 19490 27600
rect 22554 27548 22560 27600
rect 22612 27588 22618 27600
rect 23014 27588 23020 27600
rect 22612 27560 23020 27588
rect 22612 27548 22618 27560
rect 23014 27548 23020 27560
rect 23072 27548 23078 27600
rect 25792 27588 25820 27616
rect 25958 27588 25964 27600
rect 25792 27560 25964 27588
rect 25958 27548 25964 27560
rect 26016 27588 26022 27600
rect 26237 27591 26295 27597
rect 26237 27588 26249 27591
rect 26016 27560 26249 27588
rect 26016 27548 26022 27560
rect 26237 27557 26249 27560
rect 26283 27557 26295 27591
rect 26237 27551 26295 27557
rect 36449 27591 36507 27597
rect 36449 27557 36461 27591
rect 36495 27588 36507 27591
rect 38396 27588 38424 27616
rect 40310 27588 40316 27600
rect 36495 27560 38424 27588
rect 40271 27560 40316 27588
rect 36495 27557 36507 27560
rect 36449 27551 36507 27557
rect 40310 27548 40316 27560
rect 40368 27548 40374 27600
rect 5368 27492 5948 27520
rect 5368 27461 5396 27492
rect 5353 27455 5411 27461
rect 5353 27421 5365 27455
rect 5399 27421 5411 27455
rect 5353 27415 5411 27421
rect 5813 27455 5871 27461
rect 5813 27421 5825 27455
rect 5859 27421 5871 27455
rect 5920 27452 5948 27492
rect 7208 27452 7236 27548
rect 7926 27520 7932 27532
rect 7887 27492 7932 27520
rect 7926 27480 7932 27492
rect 7984 27480 7990 27532
rect 9950 27480 9956 27532
rect 10008 27520 10014 27532
rect 10137 27523 10195 27529
rect 10137 27520 10149 27523
rect 10008 27492 10149 27520
rect 10008 27480 10014 27492
rect 10137 27489 10149 27492
rect 10183 27489 10195 27523
rect 10137 27483 10195 27489
rect 12526 27480 12532 27532
rect 12584 27520 12590 27532
rect 12713 27523 12771 27529
rect 12713 27520 12725 27523
rect 12584 27492 12725 27520
rect 12584 27480 12590 27492
rect 12713 27489 12725 27492
rect 12759 27520 12771 27523
rect 13722 27520 13728 27532
rect 12759 27492 13728 27520
rect 12759 27489 12771 27492
rect 12713 27483 12771 27489
rect 13722 27480 13728 27492
rect 13780 27480 13786 27532
rect 14645 27523 14703 27529
rect 14645 27489 14657 27523
rect 14691 27520 14703 27523
rect 15010 27520 15016 27532
rect 14691 27492 15016 27520
rect 14691 27489 14703 27492
rect 14645 27483 14703 27489
rect 15010 27480 15016 27492
rect 15068 27480 15074 27532
rect 17218 27480 17224 27532
rect 17276 27520 17282 27532
rect 17604 27520 17632 27548
rect 17681 27523 17739 27529
rect 17681 27520 17693 27523
rect 17276 27492 17693 27520
rect 17276 27480 17282 27492
rect 17681 27489 17693 27492
rect 17727 27489 17739 27523
rect 17681 27483 17739 27489
rect 17865 27523 17923 27529
rect 17865 27489 17877 27523
rect 17911 27520 17923 27523
rect 18046 27520 18052 27532
rect 17911 27492 18052 27520
rect 17911 27489 17923 27492
rect 17865 27483 17923 27489
rect 18046 27480 18052 27492
rect 18104 27480 18110 27532
rect 22002 27480 22008 27532
rect 22060 27520 22066 27532
rect 24857 27523 24915 27529
rect 24857 27520 24869 27523
rect 22060 27492 24869 27520
rect 22060 27480 22066 27492
rect 24857 27489 24869 27492
rect 24903 27489 24915 27523
rect 24857 27483 24915 27489
rect 7837 27455 7895 27461
rect 7837 27452 7849 27455
rect 5920 27424 6914 27452
rect 7208 27424 7849 27452
rect 5813 27415 5871 27421
rect 5077 27387 5135 27393
rect 5077 27353 5089 27387
rect 5123 27384 5135 27387
rect 5828 27384 5856 27415
rect 6086 27393 6092 27396
rect 5123 27356 5856 27384
rect 5123 27353 5135 27356
rect 5077 27347 5135 27353
rect 6080 27347 6092 27393
rect 6144 27384 6150 27396
rect 6886 27384 6914 27424
rect 7837 27421 7849 27424
rect 7883 27421 7895 27455
rect 10226 27452 10232 27464
rect 10187 27424 10232 27452
rect 7837 27415 7895 27421
rect 10226 27412 10232 27424
rect 10284 27412 10290 27464
rect 14461 27455 14519 27461
rect 14461 27421 14473 27455
rect 14507 27452 14519 27455
rect 14550 27452 14556 27464
rect 14507 27424 14556 27452
rect 14507 27421 14519 27424
rect 14461 27415 14519 27421
rect 14550 27412 14556 27424
rect 14608 27412 14614 27464
rect 14737 27455 14795 27461
rect 14737 27421 14749 27455
rect 14783 27452 14795 27455
rect 14826 27452 14832 27464
rect 14783 27424 14832 27452
rect 14783 27421 14795 27424
rect 14737 27415 14795 27421
rect 14826 27412 14832 27424
rect 14884 27412 14890 27464
rect 17586 27452 17592 27464
rect 17547 27424 17592 27452
rect 17586 27412 17592 27424
rect 17644 27412 17650 27464
rect 17770 27412 17776 27464
rect 17828 27452 17834 27464
rect 22833 27455 22891 27461
rect 17828 27424 17873 27452
rect 17828 27412 17834 27424
rect 22833 27421 22845 27455
rect 22879 27452 22891 27455
rect 22922 27452 22928 27464
rect 22879 27424 22928 27452
rect 22879 27421 22891 27424
rect 22833 27415 22891 27421
rect 22922 27412 22928 27424
rect 22980 27412 22986 27464
rect 23014 27412 23020 27464
rect 23072 27452 23078 27464
rect 23109 27455 23167 27461
rect 23109 27452 23121 27455
rect 23072 27424 23121 27452
rect 23072 27412 23078 27424
rect 23109 27421 23121 27424
rect 23155 27421 23167 27455
rect 23109 27415 23167 27421
rect 23293 27455 23351 27461
rect 23293 27421 23305 27455
rect 23339 27452 23351 27455
rect 23382 27452 23388 27464
rect 23339 27424 23388 27452
rect 23339 27421 23351 27424
rect 23293 27415 23351 27421
rect 23382 27412 23388 27424
rect 23440 27412 23446 27464
rect 24872 27452 24900 27483
rect 30006 27480 30012 27532
rect 30064 27520 30070 27532
rect 33045 27523 33103 27529
rect 33045 27520 33057 27523
rect 30064 27492 33057 27520
rect 30064 27480 30070 27492
rect 33045 27489 33057 27492
rect 33091 27489 33103 27523
rect 41386 27520 41414 27628
rect 43898 27616 43904 27668
rect 43956 27656 43962 27668
rect 44453 27659 44511 27665
rect 43956 27628 44220 27656
rect 43956 27616 43962 27628
rect 41509 27523 41567 27529
rect 41509 27520 41521 27523
rect 41386 27492 41521 27520
rect 33045 27483 33103 27489
rect 41509 27489 41521 27492
rect 41555 27520 41567 27523
rect 44082 27520 44088 27532
rect 41555 27492 44088 27520
rect 41555 27489 41567 27492
rect 41509 27483 41567 27489
rect 44082 27480 44088 27492
rect 44140 27480 44146 27532
rect 26789 27455 26847 27461
rect 26789 27452 26801 27455
rect 24872 27424 26801 27452
rect 26789 27421 26801 27424
rect 26835 27452 26847 27455
rect 28810 27452 28816 27464
rect 26835 27424 28816 27452
rect 26835 27421 26847 27424
rect 26789 27415 26847 27421
rect 28810 27412 28816 27424
rect 28868 27412 28874 27464
rect 29638 27412 29644 27464
rect 29696 27452 29702 27464
rect 29917 27455 29975 27461
rect 29917 27452 29929 27455
rect 29696 27424 29929 27452
rect 29696 27412 29702 27424
rect 29917 27421 29929 27424
rect 29963 27421 29975 27455
rect 29917 27415 29975 27421
rect 30098 27412 30104 27464
rect 30156 27452 30162 27464
rect 30193 27455 30251 27461
rect 30193 27452 30205 27455
rect 30156 27424 30205 27452
rect 30156 27412 30162 27424
rect 30193 27421 30205 27424
rect 30239 27421 30251 27455
rect 30374 27452 30380 27464
rect 30335 27424 30380 27452
rect 30193 27415 30251 27421
rect 30374 27412 30380 27424
rect 30432 27412 30438 27464
rect 32858 27452 32864 27464
rect 32819 27424 32864 27452
rect 32858 27412 32864 27424
rect 32916 27412 32922 27464
rect 33134 27452 33140 27464
rect 33095 27424 33140 27452
rect 33134 27412 33140 27424
rect 33192 27412 33198 27464
rect 36354 27452 36360 27464
rect 36315 27424 36360 27452
rect 36354 27412 36360 27424
rect 36412 27412 36418 27464
rect 36538 27452 36544 27464
rect 36499 27424 36544 27452
rect 36538 27412 36544 27424
rect 36596 27412 36602 27464
rect 38010 27452 38016 27464
rect 37971 27424 38016 27452
rect 38010 27412 38016 27424
rect 38068 27412 38074 27464
rect 40037 27455 40095 27461
rect 40037 27421 40049 27455
rect 40083 27452 40095 27455
rect 40218 27452 40224 27464
rect 40083 27424 40224 27452
rect 40083 27421 40095 27424
rect 40037 27415 40095 27421
rect 40218 27412 40224 27424
rect 40276 27412 40282 27464
rect 41782 27452 41788 27464
rect 41743 27424 41788 27452
rect 41782 27412 41788 27424
rect 41840 27412 41846 27464
rect 43346 27412 43352 27464
rect 43404 27452 43410 27464
rect 44192 27461 44220 27628
rect 44453 27625 44465 27659
rect 44499 27656 44511 27659
rect 44726 27656 44732 27668
rect 44499 27628 44732 27656
rect 44499 27625 44511 27628
rect 44453 27619 44511 27625
rect 44726 27616 44732 27628
rect 44784 27616 44790 27668
rect 46842 27520 46848 27532
rect 46803 27492 46848 27520
rect 46842 27480 46848 27492
rect 46900 27480 46906 27532
rect 48130 27520 48136 27532
rect 48091 27492 48136 27520
rect 48130 27480 48136 27492
rect 48188 27480 48194 27532
rect 48314 27520 48320 27532
rect 48275 27492 48320 27520
rect 48314 27480 48320 27492
rect 48372 27480 48378 27532
rect 43901 27455 43959 27461
rect 43901 27452 43913 27455
rect 43404 27424 43913 27452
rect 43404 27412 43410 27424
rect 43901 27421 43913 27424
rect 43947 27421 43959 27455
rect 43901 27415 43959 27421
rect 44177 27455 44235 27461
rect 44177 27421 44189 27455
rect 44223 27421 44235 27455
rect 44177 27415 44235 27421
rect 44269 27455 44327 27461
rect 44269 27421 44281 27455
rect 44315 27452 44327 27455
rect 44358 27452 44364 27464
rect 44315 27424 44364 27452
rect 44315 27421 44327 27424
rect 44269 27415 44327 27421
rect 44358 27412 44364 27424
rect 44416 27412 44422 27464
rect 8018 27384 8024 27396
rect 6144 27356 6180 27384
rect 6886 27356 8024 27384
rect 6086 27344 6092 27347
rect 6144 27344 6150 27356
rect 8018 27344 8024 27356
rect 8076 27344 8082 27396
rect 11790 27344 11796 27396
rect 11848 27384 11854 27396
rect 12529 27387 12587 27393
rect 12529 27384 12541 27387
rect 11848 27356 12541 27384
rect 11848 27344 11854 27356
rect 12529 27353 12541 27356
rect 12575 27353 12587 27387
rect 12529 27347 12587 27353
rect 15010 27344 15016 27396
rect 15068 27384 15074 27396
rect 23750 27384 23756 27396
rect 15068 27356 23756 27384
rect 15068 27344 15074 27356
rect 23750 27344 23756 27356
rect 23808 27344 23814 27396
rect 25124 27387 25182 27393
rect 25124 27353 25136 27387
rect 25170 27384 25182 27387
rect 25222 27384 25228 27396
rect 25170 27356 25228 27384
rect 25170 27353 25182 27356
rect 25124 27347 25182 27353
rect 25222 27344 25228 27356
rect 25280 27344 25286 27396
rect 27056 27387 27114 27393
rect 27056 27353 27068 27387
rect 27102 27384 27114 27387
rect 27154 27384 27160 27396
rect 27102 27356 27160 27384
rect 27102 27353 27114 27356
rect 27056 27347 27114 27353
rect 27154 27344 27160 27356
rect 27212 27344 27218 27396
rect 40313 27387 40371 27393
rect 40313 27353 40325 27387
rect 40359 27384 40371 27387
rect 41230 27384 41236 27396
rect 40359 27356 41236 27384
rect 40359 27353 40371 27356
rect 40313 27347 40371 27353
rect 41230 27344 41236 27356
rect 41288 27384 41294 27396
rect 41506 27384 41512 27396
rect 41288 27356 41512 27384
rect 41288 27344 41294 27356
rect 41506 27344 41512 27356
rect 41564 27344 41570 27396
rect 43990 27344 43996 27396
rect 44048 27384 44054 27396
rect 44085 27387 44143 27393
rect 44085 27384 44097 27387
rect 44048 27356 44097 27384
rect 44048 27344 44054 27356
rect 44085 27353 44097 27356
rect 44131 27353 44143 27387
rect 44085 27347 44143 27353
rect 1854 27276 1860 27328
rect 1912 27316 1918 27328
rect 12621 27319 12679 27325
rect 12621 27316 12633 27319
rect 1912 27288 12633 27316
rect 1912 27276 1918 27288
rect 12621 27285 12633 27288
rect 12667 27316 12679 27319
rect 12894 27316 12900 27328
rect 12667 27288 12900 27316
rect 12667 27285 12679 27288
rect 12621 27279 12679 27285
rect 12894 27276 12900 27288
rect 12952 27276 12958 27328
rect 14277 27319 14335 27325
rect 14277 27285 14289 27319
rect 14323 27316 14335 27319
rect 14366 27316 14372 27328
rect 14323 27288 14372 27316
rect 14323 27285 14335 27288
rect 14277 27279 14335 27285
rect 14366 27276 14372 27288
rect 14424 27276 14430 27328
rect 27522 27276 27528 27328
rect 27580 27316 27586 27328
rect 28169 27319 28227 27325
rect 28169 27316 28181 27319
rect 27580 27288 28181 27316
rect 27580 27276 27586 27288
rect 28169 27285 28181 27288
rect 28215 27285 28227 27319
rect 32674 27316 32680 27328
rect 32635 27288 32680 27316
rect 28169 27279 28227 27285
rect 32674 27276 32680 27288
rect 32732 27276 32738 27328
rect 38381 27319 38439 27325
rect 38381 27285 38393 27319
rect 38427 27316 38439 27319
rect 39666 27316 39672 27328
rect 38427 27288 39672 27316
rect 38427 27285 38439 27288
rect 38381 27279 38439 27285
rect 39666 27276 39672 27288
rect 39724 27316 39730 27328
rect 40129 27319 40187 27325
rect 40129 27316 40141 27319
rect 39724 27288 40141 27316
rect 39724 27276 39730 27288
rect 40129 27285 40141 27288
rect 40175 27285 40187 27319
rect 40129 27279 40187 27285
rect 42794 27276 42800 27328
rect 42852 27316 42858 27328
rect 42889 27319 42947 27325
rect 42889 27316 42901 27319
rect 42852 27288 42901 27316
rect 42852 27276 42858 27288
rect 42889 27285 42901 27288
rect 42935 27285 42947 27319
rect 42889 27279 42947 27285
rect 47486 27276 47492 27328
rect 47544 27316 47550 27328
rect 47670 27316 47676 27328
rect 47544 27288 47676 27316
rect 47544 27276 47550 27288
rect 47670 27276 47676 27288
rect 47728 27276 47734 27328
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 5997 27115 6055 27121
rect 5997 27081 6009 27115
rect 6043 27112 6055 27115
rect 6086 27112 6092 27124
rect 6043 27084 6092 27112
rect 6043 27081 6055 27084
rect 5997 27075 6055 27081
rect 6086 27072 6092 27084
rect 6144 27072 6150 27124
rect 6733 27115 6791 27121
rect 6733 27081 6745 27115
rect 6779 27081 6791 27115
rect 6733 27075 6791 27081
rect 7101 27115 7159 27121
rect 7101 27081 7113 27115
rect 7147 27112 7159 27115
rect 11790 27112 11796 27124
rect 7147 27084 11796 27112
rect 7147 27081 7159 27084
rect 7101 27075 7159 27081
rect 5813 26979 5871 26985
rect 5813 26945 5825 26979
rect 5859 26976 5871 26979
rect 6748 26976 6776 27075
rect 11790 27072 11796 27084
rect 11848 27072 11854 27124
rect 17586 27072 17592 27124
rect 17644 27112 17650 27124
rect 17865 27115 17923 27121
rect 17865 27112 17877 27115
rect 17644 27084 17877 27112
rect 17644 27072 17650 27084
rect 17865 27081 17877 27084
rect 17911 27081 17923 27115
rect 17865 27075 17923 27081
rect 21085 27115 21143 27121
rect 21085 27081 21097 27115
rect 21131 27112 21143 27115
rect 21174 27112 21180 27124
rect 21131 27084 21180 27112
rect 21131 27081 21143 27084
rect 21085 27075 21143 27081
rect 21174 27072 21180 27084
rect 21232 27072 21238 27124
rect 25317 27115 25375 27121
rect 25317 27081 25329 27115
rect 25363 27112 25375 27115
rect 25406 27112 25412 27124
rect 25363 27084 25412 27112
rect 25363 27081 25375 27084
rect 25317 27075 25375 27081
rect 25406 27072 25412 27084
rect 25464 27072 25470 27124
rect 27798 27112 27804 27124
rect 25516 27084 27660 27112
rect 27759 27084 27804 27112
rect 9306 27044 9312 27056
rect 8220 27016 9312 27044
rect 5859 26948 6776 26976
rect 7193 26979 7251 26985
rect 5859 26945 5871 26948
rect 5813 26939 5871 26945
rect 7193 26945 7205 26979
rect 7239 26976 7251 26979
rect 7926 26976 7932 26988
rect 7239 26948 7932 26976
rect 7239 26945 7251 26948
rect 7193 26939 7251 26945
rect 7926 26936 7932 26948
rect 7984 26936 7990 26988
rect 8018 26936 8024 26988
rect 8076 26976 8082 26988
rect 8076 26948 8121 26976
rect 8076 26936 8082 26948
rect 7377 26911 7435 26917
rect 7377 26877 7389 26911
rect 7423 26908 7435 26911
rect 8220 26908 8248 27016
rect 9306 27004 9312 27016
rect 9364 27004 9370 27056
rect 9030 26985 9036 26988
rect 9024 26976 9036 26985
rect 8991 26948 9036 26976
rect 9024 26939 9036 26948
rect 9030 26936 9036 26939
rect 9088 26936 9094 26988
rect 14366 26985 14372 26988
rect 14360 26976 14372 26985
rect 14327 26948 14372 26976
rect 14360 26939 14372 26948
rect 14366 26936 14372 26939
rect 14424 26936 14430 26988
rect 16206 26936 16212 26988
rect 16264 26976 16270 26988
rect 17037 26979 17095 26985
rect 17037 26976 17049 26979
rect 16264 26948 17049 26976
rect 16264 26936 16270 26948
rect 17037 26945 17049 26948
rect 17083 26945 17095 26979
rect 17037 26939 17095 26945
rect 18049 26979 18107 26985
rect 18049 26945 18061 26979
rect 18095 26976 18107 26979
rect 18138 26976 18144 26988
rect 18095 26948 18144 26976
rect 18095 26945 18107 26948
rect 18049 26939 18107 26945
rect 18138 26936 18144 26948
rect 18196 26936 18202 26988
rect 18233 26979 18291 26985
rect 18233 26945 18245 26979
rect 18279 26945 18291 26979
rect 18233 26939 18291 26945
rect 7423 26880 8248 26908
rect 8297 26911 8355 26917
rect 7423 26877 7435 26880
rect 7377 26871 7435 26877
rect 8297 26877 8309 26911
rect 8343 26908 8355 26911
rect 8757 26911 8815 26917
rect 8757 26908 8769 26911
rect 8343 26880 8769 26908
rect 8343 26877 8355 26880
rect 8297 26871 8355 26877
rect 8757 26877 8769 26880
rect 8803 26877 8815 26911
rect 8757 26871 8815 26877
rect 13630 26868 13636 26920
rect 13688 26908 13694 26920
rect 14093 26911 14151 26917
rect 14093 26908 14105 26911
rect 13688 26880 14105 26908
rect 13688 26868 13694 26880
rect 14093 26877 14105 26880
rect 14139 26877 14151 26911
rect 17126 26908 17132 26920
rect 17087 26880 17132 26908
rect 14093 26871 14151 26877
rect 17126 26868 17132 26880
rect 17184 26868 17190 26920
rect 17405 26911 17463 26917
rect 17405 26877 17417 26911
rect 17451 26908 17463 26911
rect 17862 26908 17868 26920
rect 17451 26880 17868 26908
rect 17451 26877 17463 26880
rect 17405 26871 17463 26877
rect 17862 26868 17868 26880
rect 17920 26908 17926 26920
rect 18248 26908 18276 26939
rect 24670 26936 24676 26988
rect 24728 26976 24734 26988
rect 25516 26985 25544 27084
rect 27522 27044 27528 27056
rect 27172 27016 27528 27044
rect 25501 26979 25559 26985
rect 25501 26976 25513 26979
rect 24728 26948 25513 26976
rect 24728 26936 24734 26948
rect 25501 26945 25513 26948
rect 25547 26945 25559 26979
rect 25501 26939 25559 26945
rect 25777 26979 25835 26985
rect 25777 26945 25789 26979
rect 25823 26945 25835 26979
rect 25958 26976 25964 26988
rect 25919 26948 25964 26976
rect 25777 26939 25835 26945
rect 17920 26880 18276 26908
rect 17920 26868 17926 26880
rect 20990 26868 20996 26920
rect 21048 26908 21054 26920
rect 21177 26911 21235 26917
rect 21177 26908 21189 26911
rect 21048 26880 21189 26908
rect 21048 26868 21054 26880
rect 21177 26877 21189 26880
rect 21223 26877 21235 26911
rect 21358 26908 21364 26920
rect 21319 26880 21364 26908
rect 21177 26871 21235 26877
rect 21358 26868 21364 26880
rect 21416 26868 21422 26920
rect 25792 26908 25820 26939
rect 25958 26936 25964 26948
rect 26016 26936 26022 26988
rect 27172 26985 27200 27016
rect 27522 27004 27528 27016
rect 27580 27004 27586 27056
rect 27632 26985 27660 27084
rect 27798 27072 27804 27084
rect 27856 27072 27862 27124
rect 33134 27072 33140 27124
rect 33192 27112 33198 27124
rect 33689 27115 33747 27121
rect 33689 27112 33701 27115
rect 33192 27084 33701 27112
rect 33192 27072 33198 27084
rect 33689 27081 33701 27084
rect 33735 27112 33747 27115
rect 36538 27112 36544 27124
rect 33735 27084 36544 27112
rect 33735 27081 33747 27084
rect 33689 27075 33747 27081
rect 36538 27072 36544 27084
rect 36596 27072 36602 27124
rect 37553 27115 37611 27121
rect 37553 27081 37565 27115
rect 37599 27112 37611 27115
rect 38010 27112 38016 27124
rect 37599 27084 38016 27112
rect 37599 27081 37611 27084
rect 37553 27075 37611 27081
rect 38010 27072 38016 27084
rect 38068 27072 38074 27124
rect 32576 27047 32634 27053
rect 32576 27013 32588 27047
rect 32622 27044 32634 27047
rect 32674 27044 32680 27056
rect 32622 27016 32680 27044
rect 32622 27013 32634 27016
rect 32576 27007 32634 27013
rect 32674 27004 32680 27016
rect 32732 27004 32738 27056
rect 33410 27004 33416 27056
rect 33468 27044 33474 27056
rect 34146 27044 34152 27056
rect 33468 27016 34152 27044
rect 33468 27004 33474 27016
rect 34146 27004 34152 27016
rect 34204 27044 34210 27056
rect 36173 27047 36231 27053
rect 36173 27044 36185 27047
rect 34204 27016 36185 27044
rect 34204 27004 34210 27016
rect 36173 27013 36185 27016
rect 36219 27013 36231 27047
rect 36173 27007 36231 27013
rect 36354 27004 36360 27056
rect 36412 27044 36418 27056
rect 40129 27047 40187 27053
rect 36412 27016 37688 27044
rect 36412 27004 36418 27016
rect 27157 26979 27215 26985
rect 27157 26945 27169 26979
rect 27203 26945 27215 26979
rect 27157 26939 27215 26945
rect 27341 26979 27399 26985
rect 27341 26945 27353 26979
rect 27387 26945 27399 26979
rect 27341 26939 27399 26945
rect 27617 26979 27675 26985
rect 27617 26945 27629 26979
rect 27663 26945 27675 26979
rect 27617 26939 27675 26945
rect 35345 26979 35403 26985
rect 35345 26945 35357 26979
rect 35391 26976 35403 26979
rect 35434 26976 35440 26988
rect 35391 26948 35440 26976
rect 35391 26945 35403 26948
rect 35345 26939 35403 26945
rect 26878 26908 26884 26920
rect 25792 26880 26884 26908
rect 26878 26868 26884 26880
rect 26936 26908 26942 26920
rect 27356 26908 27384 26939
rect 35434 26936 35440 26948
rect 35492 26936 35498 26988
rect 36538 26936 36544 26988
rect 36596 26976 36602 26988
rect 37660 26985 37688 27016
rect 40129 27013 40141 27047
rect 40175 27044 40187 27047
rect 40218 27044 40224 27056
rect 40175 27016 40224 27044
rect 40175 27013 40187 27016
rect 40129 27007 40187 27013
rect 40218 27004 40224 27016
rect 40276 27004 40282 27056
rect 37461 26979 37519 26985
rect 37461 26976 37473 26979
rect 36596 26948 37473 26976
rect 36596 26936 36602 26948
rect 37461 26945 37473 26948
rect 37507 26945 37519 26979
rect 37461 26939 37519 26945
rect 37645 26979 37703 26985
rect 37645 26945 37657 26979
rect 37691 26945 37703 26979
rect 37645 26939 37703 26945
rect 38562 26936 38568 26988
rect 38620 26976 38626 26988
rect 39301 26979 39359 26985
rect 39301 26976 39313 26979
rect 38620 26948 39313 26976
rect 38620 26936 38626 26948
rect 39301 26945 39313 26948
rect 39347 26945 39359 26979
rect 39301 26939 39359 26945
rect 40313 26979 40371 26985
rect 40313 26945 40325 26979
rect 40359 26945 40371 26979
rect 40313 26939 40371 26945
rect 26936 26880 27384 26908
rect 26936 26868 26942 26880
rect 32030 26868 32036 26920
rect 32088 26908 32094 26920
rect 32309 26911 32367 26917
rect 32309 26908 32321 26911
rect 32088 26880 32321 26908
rect 32088 26868 32094 26880
rect 32309 26877 32321 26880
rect 32355 26877 32367 26911
rect 36262 26908 36268 26920
rect 36223 26880 36268 26908
rect 32309 26871 32367 26877
rect 36262 26868 36268 26880
rect 36320 26868 36326 26920
rect 36446 26908 36452 26920
rect 36407 26880 36452 26908
rect 36446 26868 36452 26880
rect 36504 26908 36510 26920
rect 37366 26908 37372 26920
rect 36504 26880 37372 26908
rect 36504 26868 36510 26880
rect 37366 26868 37372 26880
rect 37424 26868 37430 26920
rect 38838 26868 38844 26920
rect 38896 26908 38902 26920
rect 39209 26911 39267 26917
rect 39209 26908 39221 26911
rect 38896 26880 39221 26908
rect 38896 26868 38902 26880
rect 39209 26877 39221 26880
rect 39255 26877 39267 26911
rect 39666 26908 39672 26920
rect 39627 26880 39672 26908
rect 39209 26871 39267 26877
rect 39666 26868 39672 26880
rect 39724 26908 39730 26920
rect 40328 26908 40356 26939
rect 41414 26936 41420 26988
rect 41472 26976 41478 26988
rect 41877 26979 41935 26985
rect 41472 26948 41517 26976
rect 41472 26936 41478 26948
rect 41877 26945 41889 26979
rect 41923 26976 41935 26979
rect 42886 26976 42892 26988
rect 41923 26948 42892 26976
rect 41923 26945 41935 26948
rect 41877 26939 41935 26945
rect 42886 26936 42892 26948
rect 42944 26936 42950 26988
rect 43901 26979 43959 26985
rect 43901 26945 43913 26979
rect 43947 26976 43959 26979
rect 43990 26976 43996 26988
rect 43947 26948 43996 26976
rect 43947 26945 43959 26948
rect 43901 26939 43959 26945
rect 43990 26936 43996 26948
rect 44048 26936 44054 26988
rect 44174 26985 44180 26988
rect 44168 26939 44180 26985
rect 44232 26976 44238 26988
rect 44232 26948 44268 26976
rect 44174 26936 44180 26939
rect 44232 26936 44238 26948
rect 46750 26936 46756 26988
rect 46808 26976 46814 26988
rect 46845 26979 46903 26985
rect 46845 26976 46857 26979
rect 46808 26948 46857 26976
rect 46808 26936 46814 26948
rect 46845 26945 46857 26948
rect 46891 26976 46903 26979
rect 47118 26976 47124 26988
rect 46891 26948 47124 26976
rect 46891 26945 46903 26948
rect 46845 26939 46903 26945
rect 47118 26936 47124 26948
rect 47176 26936 47182 26988
rect 47394 26936 47400 26988
rect 47452 26976 47458 26988
rect 47762 26976 47768 26988
rect 47452 26948 47768 26976
rect 47452 26936 47458 26948
rect 47762 26936 47768 26948
rect 47820 26936 47826 26988
rect 42058 26908 42064 26920
rect 39724 26880 40356 26908
rect 41971 26880 42064 26908
rect 39724 26868 39730 26880
rect 42058 26868 42064 26880
rect 42116 26908 42122 26920
rect 42978 26908 42984 26920
rect 42116 26880 42984 26908
rect 42116 26868 42122 26880
rect 42978 26868 42984 26880
rect 43036 26868 43042 26920
rect 10134 26772 10140 26784
rect 10095 26744 10140 26772
rect 10134 26732 10140 26744
rect 10192 26732 10198 26784
rect 15194 26732 15200 26784
rect 15252 26772 15258 26784
rect 15473 26775 15531 26781
rect 15473 26772 15485 26775
rect 15252 26744 15485 26772
rect 15252 26732 15258 26744
rect 15473 26741 15485 26744
rect 15519 26741 15531 26775
rect 15473 26735 15531 26741
rect 20717 26775 20775 26781
rect 20717 26741 20729 26775
rect 20763 26772 20775 26775
rect 20806 26772 20812 26784
rect 20763 26744 20812 26772
rect 20763 26741 20775 26744
rect 20717 26735 20775 26741
rect 20806 26732 20812 26744
rect 20864 26732 20870 26784
rect 23566 26732 23572 26784
rect 23624 26772 23630 26784
rect 24854 26772 24860 26784
rect 23624 26744 24860 26772
rect 23624 26732 23630 26744
rect 24854 26732 24860 26744
rect 24912 26732 24918 26784
rect 35161 26775 35219 26781
rect 35161 26741 35173 26775
rect 35207 26772 35219 26775
rect 35342 26772 35348 26784
rect 35207 26744 35348 26772
rect 35207 26741 35219 26744
rect 35161 26735 35219 26741
rect 35342 26732 35348 26744
rect 35400 26732 35406 26784
rect 35802 26772 35808 26784
rect 35763 26744 35808 26772
rect 35802 26732 35808 26744
rect 35860 26732 35866 26784
rect 40494 26772 40500 26784
rect 40455 26744 40500 26772
rect 40494 26732 40500 26744
rect 40552 26732 40558 26784
rect 45278 26772 45284 26784
rect 45239 26744 45284 26772
rect 45278 26732 45284 26744
rect 45336 26732 45342 26784
rect 46658 26732 46664 26784
rect 46716 26772 46722 26784
rect 46753 26775 46811 26781
rect 46753 26772 46765 26775
rect 46716 26744 46765 26772
rect 46716 26732 46722 26744
rect 46753 26741 46765 26744
rect 46799 26741 46811 26775
rect 46753 26735 46811 26741
rect 47857 26775 47915 26781
rect 47857 26741 47869 26775
rect 47903 26772 47915 26775
rect 48130 26772 48136 26784
rect 47903 26744 48136 26772
rect 47903 26741 47915 26744
rect 47857 26735 47915 26741
rect 48130 26732 48136 26744
rect 48188 26732 48194 26784
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 9950 26568 9956 26580
rect 9911 26540 9956 26568
rect 9950 26528 9956 26540
rect 10008 26528 10014 26580
rect 14550 26568 14556 26580
rect 14511 26540 14556 26568
rect 14550 26528 14556 26540
rect 14608 26528 14614 26580
rect 17770 26528 17776 26580
rect 17828 26568 17834 26580
rect 18141 26571 18199 26577
rect 18141 26568 18153 26571
rect 17828 26540 18153 26568
rect 17828 26528 17834 26540
rect 18141 26537 18153 26540
rect 18187 26537 18199 26571
rect 23566 26568 23572 26580
rect 18141 26531 18199 26537
rect 22066 26540 23572 26568
rect 20441 26503 20499 26509
rect 20441 26469 20453 26503
rect 20487 26469 20499 26503
rect 20441 26463 20499 26469
rect 9677 26435 9735 26441
rect 9677 26401 9689 26435
rect 9723 26432 9735 26435
rect 10134 26432 10140 26444
rect 9723 26404 10140 26432
rect 9723 26401 9735 26404
rect 9677 26395 9735 26401
rect 10134 26392 10140 26404
rect 10192 26392 10198 26444
rect 17221 26435 17279 26441
rect 17221 26432 17233 26435
rect 16546 26404 17233 26432
rect 9582 26364 9588 26376
rect 9543 26336 9588 26364
rect 9582 26324 9588 26336
rect 9640 26324 9646 26376
rect 12250 26364 12256 26376
rect 12211 26336 12256 26364
rect 12250 26324 12256 26336
rect 12308 26324 12314 26376
rect 14550 26324 14556 26376
rect 14608 26364 14614 26376
rect 14737 26367 14795 26373
rect 14737 26364 14749 26367
rect 14608 26336 14749 26364
rect 14608 26324 14614 26336
rect 14737 26333 14749 26336
rect 14783 26333 14795 26367
rect 14737 26327 14795 26333
rect 14918 26324 14924 26376
rect 14976 26364 14982 26376
rect 15013 26367 15071 26373
rect 15013 26364 15025 26367
rect 14976 26336 15025 26364
rect 14976 26324 14982 26336
rect 15013 26333 15025 26336
rect 15059 26333 15071 26367
rect 15194 26364 15200 26376
rect 15155 26336 15200 26364
rect 15013 26327 15071 26333
rect 15194 26324 15200 26336
rect 15252 26364 15258 26376
rect 16206 26364 16212 26376
rect 15252 26336 16212 26364
rect 15252 26324 15258 26336
rect 16206 26324 16212 26336
rect 16264 26364 16270 26376
rect 16546 26364 16574 26404
rect 17221 26401 17233 26404
rect 17267 26401 17279 26435
rect 17221 26395 17279 26401
rect 17589 26435 17647 26441
rect 17589 26401 17601 26435
rect 17635 26432 17647 26435
rect 17770 26432 17776 26444
rect 17635 26404 17776 26432
rect 17635 26401 17647 26404
rect 17589 26395 17647 26401
rect 17770 26392 17776 26404
rect 17828 26392 17834 26444
rect 18138 26392 18144 26444
rect 18196 26392 18202 26444
rect 17126 26364 17132 26376
rect 16264 26336 16574 26364
rect 17087 26336 17132 26364
rect 16264 26324 16270 26336
rect 17126 26324 17132 26336
rect 17184 26324 17190 26376
rect 17862 26324 17868 26376
rect 17920 26364 17926 26376
rect 18049 26367 18107 26373
rect 18049 26364 18061 26367
rect 17920 26336 18061 26364
rect 17920 26324 17926 26336
rect 18049 26333 18061 26336
rect 18095 26333 18107 26367
rect 18156 26364 18184 26392
rect 18233 26367 18291 26373
rect 18233 26364 18245 26367
rect 18156 26336 18245 26364
rect 18049 26327 18107 26333
rect 18233 26333 18245 26336
rect 18279 26333 18291 26367
rect 18233 26327 18291 26333
rect 19797 26367 19855 26373
rect 19797 26333 19809 26367
rect 19843 26364 19855 26367
rect 20456 26364 20484 26463
rect 21358 26460 21364 26512
rect 21416 26500 21422 26512
rect 22066 26500 22094 26540
rect 23566 26528 23572 26540
rect 23624 26528 23630 26580
rect 23750 26568 23756 26580
rect 23663 26540 23756 26568
rect 23750 26528 23756 26540
rect 23808 26568 23814 26580
rect 26234 26568 26240 26580
rect 23808 26540 26240 26568
rect 23808 26528 23814 26540
rect 26234 26528 26240 26540
rect 26292 26568 26298 26580
rect 26970 26568 26976 26580
rect 26292 26540 26976 26568
rect 26292 26528 26298 26540
rect 26970 26528 26976 26540
rect 27028 26528 27034 26580
rect 33410 26568 33416 26580
rect 33371 26540 33416 26568
rect 33410 26528 33416 26540
rect 33468 26528 33474 26580
rect 36262 26528 36268 26580
rect 36320 26568 36326 26580
rect 36725 26571 36783 26577
rect 36725 26568 36737 26571
rect 36320 26540 36737 26568
rect 36320 26528 36326 26540
rect 36725 26537 36737 26540
rect 36771 26537 36783 26571
rect 38933 26571 38991 26577
rect 38933 26568 38945 26571
rect 36725 26531 36783 26537
rect 37016 26540 38945 26568
rect 24026 26500 24032 26512
rect 21416 26472 22094 26500
rect 22664 26472 24032 26500
rect 21416 26460 21422 26472
rect 21085 26435 21143 26441
rect 21085 26401 21097 26435
rect 21131 26432 21143 26435
rect 22370 26432 22376 26444
rect 21131 26404 22376 26432
rect 21131 26401 21143 26404
rect 21085 26395 21143 26401
rect 22370 26392 22376 26404
rect 22428 26432 22434 26444
rect 22664 26432 22692 26472
rect 24026 26460 24032 26472
rect 24084 26460 24090 26512
rect 31938 26500 31944 26512
rect 25700 26472 31944 26500
rect 24581 26435 24639 26441
rect 24581 26432 24593 26435
rect 22428 26404 22692 26432
rect 23584 26404 24593 26432
rect 22428 26392 22434 26404
rect 20806 26364 20812 26376
rect 19843 26336 20484 26364
rect 20767 26336 20812 26364
rect 19843 26333 19855 26336
rect 19797 26327 19855 26333
rect 20806 26324 20812 26336
rect 20864 26324 20870 26376
rect 23584 26373 23612 26404
rect 24581 26401 24593 26404
rect 24627 26401 24639 26435
rect 25700 26432 25728 26472
rect 31938 26460 31944 26472
rect 31996 26460 32002 26512
rect 32030 26432 32036 26444
rect 24581 26395 24639 26401
rect 24688 26404 25728 26432
rect 31726 26404 32036 26432
rect 23569 26367 23627 26373
rect 23569 26333 23581 26367
rect 23615 26333 23627 26367
rect 23569 26327 23627 26333
rect 23845 26367 23903 26373
rect 23845 26333 23857 26367
rect 23891 26364 23903 26367
rect 23934 26364 23940 26376
rect 23891 26336 23940 26364
rect 23891 26333 23903 26336
rect 23845 26327 23903 26333
rect 23934 26324 23940 26336
rect 23992 26364 23998 26376
rect 24688 26364 24716 26404
rect 23992 26336 24716 26364
rect 24765 26367 24823 26373
rect 23992 26324 23998 26336
rect 24765 26333 24777 26367
rect 24811 26333 24823 26367
rect 24765 26327 24823 26333
rect 25041 26367 25099 26373
rect 25041 26333 25053 26367
rect 25087 26333 25099 26367
rect 25222 26364 25228 26376
rect 25183 26336 25228 26364
rect 25041 26327 25099 26333
rect 24670 26256 24676 26308
rect 24728 26296 24734 26308
rect 24780 26296 24808 26327
rect 24728 26268 24808 26296
rect 25056 26296 25084 26327
rect 25222 26324 25228 26336
rect 25280 26324 25286 26376
rect 25961 26367 26019 26373
rect 25961 26333 25973 26367
rect 26007 26364 26019 26367
rect 26142 26364 26148 26376
rect 26007 26336 26148 26364
rect 26007 26333 26019 26336
rect 25961 26327 26019 26333
rect 26142 26324 26148 26336
rect 26200 26324 26206 26376
rect 26878 26296 26884 26308
rect 25056 26268 26884 26296
rect 24728 26256 24734 26268
rect 26878 26256 26884 26268
rect 26936 26256 26942 26308
rect 12066 26228 12072 26240
rect 12027 26200 12072 26228
rect 12066 26188 12072 26200
rect 12124 26188 12130 26240
rect 16945 26231 17003 26237
rect 16945 26197 16957 26231
rect 16991 26228 17003 26231
rect 17034 26228 17040 26240
rect 16991 26200 17040 26228
rect 16991 26197 17003 26200
rect 16945 26191 17003 26197
rect 17034 26188 17040 26200
rect 17092 26188 17098 26240
rect 19978 26228 19984 26240
rect 19939 26200 19984 26228
rect 19978 26188 19984 26200
rect 20036 26188 20042 26240
rect 20901 26231 20959 26237
rect 20901 26197 20913 26231
rect 20947 26228 20959 26231
rect 21450 26228 21456 26240
rect 20947 26200 21456 26228
rect 20947 26197 20959 26200
rect 20901 26191 20959 26197
rect 21450 26188 21456 26200
rect 21508 26188 21514 26240
rect 23382 26228 23388 26240
rect 23343 26200 23388 26228
rect 23382 26188 23388 26200
rect 23440 26188 23446 26240
rect 31110 26188 31116 26240
rect 31168 26228 31174 26240
rect 31726 26228 31754 26404
rect 32030 26392 32036 26404
rect 32088 26392 32094 26444
rect 37016 26441 37044 26540
rect 38933 26537 38945 26540
rect 38979 26537 38991 26571
rect 44174 26568 44180 26580
rect 44135 26540 44180 26568
rect 38933 26531 38991 26537
rect 44174 26528 44180 26540
rect 44232 26528 44238 26580
rect 37921 26503 37979 26509
rect 37921 26469 37933 26503
rect 37967 26500 37979 26503
rect 38378 26500 38384 26512
rect 37967 26472 38384 26500
rect 37967 26469 37979 26472
rect 37921 26463 37979 26469
rect 38378 26460 38384 26472
rect 38436 26460 38442 26512
rect 40037 26503 40095 26509
rect 40037 26500 40049 26503
rect 39132 26472 40049 26500
rect 37001 26435 37059 26441
rect 37001 26401 37013 26435
rect 37047 26401 37059 26435
rect 37737 26435 37795 26441
rect 37737 26432 37749 26435
rect 37001 26395 37059 26401
rect 37108 26404 37749 26432
rect 34238 26324 34244 26376
rect 34296 26364 34302 26376
rect 37108 26373 37136 26404
rect 37737 26401 37749 26404
rect 37783 26401 37795 26435
rect 37737 26395 37795 26401
rect 38010 26392 38016 26444
rect 38068 26432 38074 26444
rect 38197 26435 38255 26441
rect 38197 26432 38209 26435
rect 38068 26404 38209 26432
rect 38068 26392 38074 26404
rect 38197 26401 38209 26404
rect 38243 26401 38255 26435
rect 38197 26395 38255 26401
rect 34885 26367 34943 26373
rect 34885 26364 34897 26367
rect 34296 26336 34897 26364
rect 34296 26324 34302 26336
rect 34885 26333 34897 26336
rect 34931 26333 34943 26367
rect 34885 26327 34943 26333
rect 37093 26367 37151 26373
rect 37093 26333 37105 26367
rect 37139 26333 37151 26367
rect 37093 26327 37151 26333
rect 38838 26324 38844 26376
rect 38896 26364 38902 26376
rect 39132 26373 39160 26472
rect 40037 26469 40049 26472
rect 40083 26469 40095 26503
rect 40037 26463 40095 26469
rect 39666 26432 39672 26444
rect 39316 26404 39672 26432
rect 39316 26373 39344 26404
rect 39666 26392 39672 26404
rect 39724 26392 39730 26444
rect 40218 26392 40224 26444
rect 40276 26392 40282 26444
rect 46474 26432 46480 26444
rect 46435 26404 46480 26432
rect 46474 26392 46480 26404
rect 46532 26392 46538 26444
rect 46658 26432 46664 26444
rect 46619 26404 46664 26432
rect 46658 26392 46664 26404
rect 46716 26392 46722 26444
rect 47946 26432 47952 26444
rect 47907 26404 47952 26432
rect 47946 26392 47952 26404
rect 48004 26392 48010 26444
rect 39117 26367 39175 26373
rect 39117 26364 39129 26367
rect 38896 26336 39129 26364
rect 38896 26324 38902 26336
rect 39117 26333 39129 26336
rect 39163 26333 39175 26367
rect 39117 26327 39175 26333
rect 39301 26367 39359 26373
rect 39301 26333 39313 26367
rect 39347 26333 39359 26367
rect 39301 26327 39359 26333
rect 39485 26367 39543 26373
rect 39485 26333 39497 26367
rect 39531 26364 39543 26367
rect 40236 26364 40264 26392
rect 39531 26336 40264 26364
rect 39531 26333 39543 26336
rect 39485 26327 39543 26333
rect 40862 26324 40868 26376
rect 40920 26364 40926 26376
rect 41417 26367 41475 26373
rect 41417 26364 41429 26367
rect 40920 26336 41429 26364
rect 40920 26324 40926 26336
rect 41417 26333 41429 26336
rect 41463 26333 41475 26367
rect 43990 26364 43996 26376
rect 43951 26336 43996 26364
rect 41417 26327 41475 26333
rect 43990 26324 43996 26336
rect 44048 26324 44054 26376
rect 32306 26305 32312 26308
rect 32300 26259 32312 26305
rect 32364 26296 32370 26308
rect 35152 26299 35210 26305
rect 32364 26268 32400 26296
rect 32306 26256 32312 26259
rect 32364 26256 32370 26268
rect 35152 26265 35164 26299
rect 35198 26296 35210 26299
rect 35342 26296 35348 26308
rect 35198 26268 35348 26296
rect 35198 26265 35210 26268
rect 35152 26259 35210 26265
rect 35342 26256 35348 26268
rect 35400 26256 35406 26308
rect 38562 26256 38568 26308
rect 38620 26296 38626 26308
rect 39209 26299 39267 26305
rect 39209 26296 39221 26299
rect 38620 26268 39221 26296
rect 38620 26256 38626 26268
rect 39209 26265 39221 26268
rect 39255 26265 39267 26299
rect 39209 26259 39267 26265
rect 40218 26256 40224 26308
rect 40276 26296 40282 26308
rect 41150 26299 41208 26305
rect 41150 26296 41162 26299
rect 40276 26268 41162 26296
rect 40276 26256 40282 26268
rect 41150 26265 41162 26268
rect 41196 26265 41208 26299
rect 41150 26259 41208 26265
rect 31168 26200 31754 26228
rect 36265 26231 36323 26237
rect 31168 26188 31174 26200
rect 36265 26197 36277 26231
rect 36311 26228 36323 26231
rect 36354 26228 36360 26240
rect 36311 26200 36360 26228
rect 36311 26197 36323 26200
rect 36265 26191 36323 26197
rect 36354 26188 36360 26200
rect 36412 26188 36418 26240
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 7926 26024 7932 26036
rect 7887 25996 7932 26024
rect 7926 25984 7932 25996
rect 7984 25984 7990 26036
rect 21450 26024 21456 26036
rect 21411 25996 21456 26024
rect 21450 25984 21456 25996
rect 21508 25984 21514 26036
rect 22002 25984 22008 26036
rect 22060 26024 22066 26036
rect 24305 26027 24363 26033
rect 22060 25996 22968 26024
rect 22060 25984 22066 25996
rect 11968 25959 12026 25965
rect 11968 25925 11980 25959
rect 12014 25956 12026 25959
rect 12066 25956 12072 25968
rect 12014 25928 12072 25956
rect 12014 25925 12026 25928
rect 11968 25919 12026 25925
rect 12066 25916 12072 25928
rect 12124 25916 12130 25968
rect 18417 25959 18475 25965
rect 18417 25925 18429 25959
rect 18463 25956 18475 25959
rect 18506 25956 18512 25968
rect 18463 25928 18512 25956
rect 18463 25925 18475 25928
rect 18417 25919 18475 25925
rect 18506 25916 18512 25928
rect 18564 25956 18570 25968
rect 18564 25928 19196 25956
rect 18564 25916 18570 25928
rect 6816 25891 6874 25897
rect 6816 25857 6828 25891
rect 6862 25888 6874 25891
rect 7098 25888 7104 25900
rect 6862 25860 7104 25888
rect 6862 25857 6874 25860
rect 6816 25851 6874 25857
rect 7098 25848 7104 25860
rect 7156 25848 7162 25900
rect 17773 25891 17831 25897
rect 17773 25857 17785 25891
rect 17819 25888 17831 25891
rect 17862 25888 17868 25900
rect 17819 25860 17868 25888
rect 17819 25857 17831 25860
rect 17773 25851 17831 25857
rect 17862 25848 17868 25860
rect 17920 25848 17926 25900
rect 18601 25891 18659 25897
rect 18601 25857 18613 25891
rect 18647 25857 18659 25891
rect 18601 25851 18659 25857
rect 18693 25891 18751 25897
rect 18693 25857 18705 25891
rect 18739 25888 18751 25891
rect 18874 25888 18880 25900
rect 18739 25860 18880 25888
rect 18739 25857 18751 25860
rect 18693 25851 18751 25857
rect 6454 25780 6460 25832
rect 6512 25820 6518 25832
rect 6549 25823 6607 25829
rect 6549 25820 6561 25823
rect 6512 25792 6561 25820
rect 6512 25780 6518 25792
rect 6549 25789 6561 25792
rect 6595 25789 6607 25823
rect 6549 25783 6607 25789
rect 11701 25823 11759 25829
rect 11701 25789 11713 25823
rect 11747 25789 11759 25823
rect 11701 25783 11759 25789
rect 2317 25687 2375 25693
rect 2317 25653 2329 25687
rect 2363 25684 2375 25687
rect 3418 25684 3424 25696
rect 2363 25656 3424 25684
rect 2363 25653 2375 25656
rect 2317 25647 2375 25653
rect 3418 25644 3424 25656
rect 3476 25644 3482 25696
rect 11716 25684 11744 25783
rect 18138 25712 18144 25764
rect 18196 25752 18202 25764
rect 18417 25755 18475 25761
rect 18417 25752 18429 25755
rect 18196 25724 18429 25752
rect 18196 25712 18202 25724
rect 18417 25721 18429 25724
rect 18463 25721 18475 25755
rect 18616 25752 18644 25851
rect 18874 25848 18880 25860
rect 18932 25848 18938 25900
rect 19168 25897 19196 25928
rect 19978 25916 19984 25968
rect 20036 25956 20042 25968
rect 20318 25959 20376 25965
rect 20318 25956 20330 25959
rect 20036 25928 20330 25956
rect 20036 25916 20042 25928
rect 20318 25925 20330 25928
rect 20364 25925 20376 25959
rect 20318 25919 20376 25925
rect 19153 25891 19211 25897
rect 19153 25857 19165 25891
rect 19199 25888 19211 25891
rect 21468 25888 21496 25984
rect 22940 25897 22968 25996
rect 24305 25993 24317 26027
rect 24351 26024 24363 26027
rect 25222 26024 25228 26036
rect 24351 25996 25228 26024
rect 24351 25993 24363 25996
rect 24305 25987 24363 25993
rect 23192 25959 23250 25965
rect 23192 25925 23204 25959
rect 23238 25956 23250 25959
rect 23382 25956 23388 25968
rect 23238 25928 23388 25956
rect 23238 25925 23250 25928
rect 23192 25919 23250 25925
rect 23382 25916 23388 25928
rect 23440 25916 23446 25968
rect 22005 25891 22063 25897
rect 22005 25888 22017 25891
rect 19199 25860 21128 25888
rect 21468 25860 22017 25888
rect 19199 25857 19211 25860
rect 19153 25851 19211 25857
rect 20073 25823 20131 25829
rect 20073 25789 20085 25823
rect 20119 25789 20131 25823
rect 20073 25783 20131 25789
rect 19518 25752 19524 25764
rect 18616 25724 19524 25752
rect 18417 25715 18475 25721
rect 19518 25712 19524 25724
rect 19576 25712 19582 25764
rect 12434 25684 12440 25696
rect 11716 25656 12440 25684
rect 12434 25644 12440 25656
rect 12492 25644 12498 25696
rect 13078 25684 13084 25696
rect 13039 25656 13084 25684
rect 13078 25644 13084 25656
rect 13136 25644 13142 25696
rect 17865 25687 17923 25693
rect 17865 25653 17877 25687
rect 17911 25684 17923 25687
rect 18598 25684 18604 25696
rect 17911 25656 18604 25684
rect 17911 25653 17923 25656
rect 17865 25647 17923 25653
rect 18598 25644 18604 25656
rect 18656 25644 18662 25696
rect 19610 25684 19616 25696
rect 19571 25656 19616 25684
rect 19610 25644 19616 25656
rect 19668 25644 19674 25696
rect 20088 25684 20116 25783
rect 21100 25752 21128 25860
rect 22005 25857 22017 25860
rect 22051 25857 22063 25891
rect 22005 25851 22063 25857
rect 22189 25891 22247 25897
rect 22189 25857 22201 25891
rect 22235 25857 22247 25891
rect 22189 25851 22247 25857
rect 22925 25891 22983 25897
rect 22925 25857 22937 25891
rect 22971 25857 22983 25891
rect 24320 25888 24348 25987
rect 25222 25984 25228 25996
rect 25280 25984 25286 26036
rect 31662 26024 31668 26036
rect 31588 25996 31668 26024
rect 26510 25956 26516 25968
rect 26252 25928 26516 25956
rect 22925 25851 22983 25857
rect 23032 25860 24348 25888
rect 21634 25780 21640 25832
rect 21692 25820 21698 25832
rect 22204 25820 22232 25851
rect 23032 25820 23060 25860
rect 24946 25848 24952 25900
rect 25004 25888 25010 25900
rect 25317 25891 25375 25897
rect 25317 25888 25329 25891
rect 25004 25860 25329 25888
rect 25004 25848 25010 25860
rect 25317 25857 25329 25860
rect 25363 25888 25375 25891
rect 25682 25888 25688 25900
rect 25363 25860 25688 25888
rect 25363 25857 25375 25860
rect 25317 25851 25375 25857
rect 25682 25848 25688 25860
rect 25740 25848 25746 25900
rect 26252 25897 26280 25928
rect 26510 25916 26516 25928
rect 26568 25916 26574 25968
rect 26237 25891 26295 25897
rect 26237 25857 26249 25891
rect 26283 25857 26295 25891
rect 26237 25851 26295 25857
rect 26421 25891 26479 25897
rect 26421 25857 26433 25891
rect 26467 25888 26479 25891
rect 27154 25888 27160 25900
rect 26467 25860 27160 25888
rect 26467 25857 26479 25860
rect 26421 25851 26479 25857
rect 27154 25848 27160 25860
rect 27212 25848 27218 25900
rect 30673 25891 30731 25897
rect 30673 25857 30685 25891
rect 30719 25888 30731 25891
rect 31202 25888 31208 25900
rect 30719 25860 31208 25888
rect 30719 25857 30731 25860
rect 30673 25851 30731 25857
rect 31202 25848 31208 25860
rect 31260 25848 31266 25900
rect 31588 25832 31616 25996
rect 31662 25984 31668 25996
rect 31720 25984 31726 26036
rect 32858 25984 32864 26036
rect 32916 26024 32922 26036
rect 33045 26027 33103 26033
rect 33045 26024 33057 26027
rect 32916 25996 33057 26024
rect 32916 25984 32922 25996
rect 33045 25993 33057 25996
rect 33091 25993 33103 26027
rect 35434 26024 35440 26036
rect 35395 25996 35440 26024
rect 33045 25987 33103 25993
rect 35434 25984 35440 25996
rect 35492 25984 35498 26036
rect 35802 25984 35808 26036
rect 35860 26024 35866 26036
rect 35897 26027 35955 26033
rect 35897 26024 35909 26027
rect 35860 25996 35909 26024
rect 35860 25984 35866 25996
rect 35897 25993 35909 25996
rect 35943 25993 35955 26027
rect 35897 25987 35955 25993
rect 40221 26027 40279 26033
rect 40221 25993 40233 26027
rect 40267 26024 40279 26027
rect 40494 26024 40500 26036
rect 40267 25996 40500 26024
rect 40267 25993 40279 25996
rect 40221 25987 40279 25993
rect 40494 25984 40500 25996
rect 40552 25984 40558 26036
rect 43809 26027 43867 26033
rect 43809 25993 43821 26027
rect 43855 26024 43867 26027
rect 43990 26024 43996 26036
rect 43855 25996 43996 26024
rect 43855 25993 43867 25996
rect 43809 25987 43867 25993
rect 43990 25984 43996 25996
rect 44048 25984 44054 26036
rect 31754 25916 31760 25968
rect 31812 25956 31818 25968
rect 40126 25956 40132 25968
rect 31812 25928 32904 25956
rect 31812 25916 31818 25928
rect 32876 25900 32904 25928
rect 34808 25928 40132 25956
rect 34808 25900 34836 25928
rect 40126 25916 40132 25928
rect 40184 25916 40190 25968
rect 32401 25891 32459 25897
rect 32401 25857 32413 25891
rect 32447 25857 32459 25891
rect 32582 25888 32588 25900
rect 32543 25860 32588 25888
rect 32401 25851 32459 25857
rect 25590 25820 25596 25832
rect 21692 25792 23060 25820
rect 25551 25792 25596 25820
rect 21692 25780 21698 25792
rect 25590 25780 25596 25792
rect 25648 25780 25654 25832
rect 30929 25823 30987 25829
rect 30929 25789 30941 25823
rect 30975 25820 30987 25823
rect 31110 25820 31116 25832
rect 30975 25792 31116 25820
rect 30975 25789 30987 25792
rect 30929 25783 30987 25789
rect 31110 25780 31116 25792
rect 31168 25780 31174 25832
rect 31570 25780 31576 25832
rect 31628 25780 31634 25832
rect 32416 25820 32444 25851
rect 32582 25848 32588 25860
rect 32640 25848 32646 25900
rect 32858 25888 32864 25900
rect 32819 25860 32864 25888
rect 32858 25848 32864 25860
rect 32916 25848 32922 25900
rect 33134 25848 33140 25900
rect 33192 25888 33198 25900
rect 33873 25891 33931 25897
rect 33873 25888 33885 25891
rect 33192 25860 33885 25888
rect 33192 25848 33198 25860
rect 33873 25857 33885 25860
rect 33919 25888 33931 25891
rect 34790 25888 34796 25900
rect 33919 25860 34796 25888
rect 33919 25857 33931 25860
rect 33873 25851 33931 25857
rect 34790 25848 34796 25860
rect 34848 25848 34854 25900
rect 35805 25891 35863 25897
rect 35805 25857 35817 25891
rect 35851 25888 35863 25891
rect 36354 25888 36360 25900
rect 35851 25860 36360 25888
rect 35851 25857 35863 25860
rect 35805 25851 35863 25857
rect 36354 25848 36360 25860
rect 36412 25848 36418 25900
rect 38010 25888 38016 25900
rect 37971 25860 38016 25888
rect 38010 25848 38016 25860
rect 38068 25848 38074 25900
rect 38105 25891 38163 25897
rect 38105 25857 38117 25891
rect 38151 25857 38163 25891
rect 38105 25851 38163 25857
rect 38197 25891 38255 25897
rect 38197 25857 38209 25891
rect 38243 25888 38255 25891
rect 38838 25888 38844 25900
rect 38243 25860 38844 25888
rect 38243 25857 38255 25860
rect 38197 25851 38255 25857
rect 32674 25820 32680 25832
rect 32416 25792 32680 25820
rect 32674 25780 32680 25792
rect 32732 25780 32738 25832
rect 34238 25780 34244 25832
rect 34296 25820 34302 25832
rect 34609 25823 34667 25829
rect 34609 25820 34621 25823
rect 34296 25792 34621 25820
rect 34296 25780 34302 25792
rect 34609 25789 34621 25792
rect 34655 25789 34667 25823
rect 34609 25783 34667 25789
rect 36081 25823 36139 25829
rect 36081 25789 36093 25823
rect 36127 25820 36139 25823
rect 36630 25820 36636 25832
rect 36127 25792 36636 25820
rect 36127 25789 36139 25792
rect 36081 25783 36139 25789
rect 36630 25780 36636 25792
rect 36688 25820 36694 25832
rect 37182 25820 37188 25832
rect 36688 25792 37188 25820
rect 36688 25780 36694 25792
rect 37182 25780 37188 25792
rect 37240 25780 37246 25832
rect 22005 25755 22063 25761
rect 22005 25752 22017 25755
rect 21100 25724 22017 25752
rect 22005 25721 22017 25724
rect 22051 25721 22063 25755
rect 38120 25752 38148 25851
rect 38838 25848 38844 25860
rect 38896 25848 38902 25900
rect 39022 25888 39028 25900
rect 38983 25860 39028 25888
rect 39022 25848 39028 25860
rect 39080 25848 39086 25900
rect 39117 25891 39175 25897
rect 39117 25857 39129 25891
rect 39163 25857 39175 25891
rect 39117 25851 39175 25857
rect 39209 25891 39267 25897
rect 39209 25857 39221 25891
rect 39255 25857 39267 25891
rect 40037 25891 40095 25897
rect 40037 25888 40049 25891
rect 39209 25851 39267 25857
rect 39408 25860 40049 25888
rect 38378 25780 38384 25832
rect 38436 25820 38442 25832
rect 39132 25820 39160 25851
rect 38436 25792 39160 25820
rect 38436 25780 38442 25792
rect 38562 25752 38568 25764
rect 38120 25724 38568 25752
rect 22005 25715 22063 25721
rect 38562 25712 38568 25724
rect 38620 25712 38626 25764
rect 38654 25712 38660 25764
rect 38712 25752 38718 25764
rect 39224 25752 39252 25851
rect 39408 25761 39436 25860
rect 40037 25857 40049 25860
rect 40083 25857 40095 25891
rect 40310 25888 40316 25900
rect 40271 25860 40316 25888
rect 40037 25851 40095 25857
rect 40310 25848 40316 25860
rect 40368 25848 40374 25900
rect 44177 25891 44235 25897
rect 44177 25857 44189 25891
rect 44223 25888 44235 25891
rect 45186 25888 45192 25900
rect 44223 25860 45192 25888
rect 44223 25857 44235 25860
rect 44177 25851 44235 25857
rect 45186 25848 45192 25860
rect 45244 25848 45250 25900
rect 39853 25823 39911 25829
rect 39853 25789 39865 25823
rect 39899 25820 39911 25823
rect 40218 25820 40224 25832
rect 39899 25792 40224 25820
rect 39899 25789 39911 25792
rect 39853 25783 39911 25789
rect 40218 25780 40224 25792
rect 40276 25780 40282 25832
rect 43070 25780 43076 25832
rect 43128 25820 43134 25832
rect 43990 25820 43996 25832
rect 43128 25792 43996 25820
rect 43128 25780 43134 25792
rect 43990 25780 43996 25792
rect 44048 25820 44054 25832
rect 44269 25823 44327 25829
rect 44269 25820 44281 25823
rect 44048 25792 44281 25820
rect 44048 25780 44054 25792
rect 44269 25789 44281 25792
rect 44315 25789 44327 25823
rect 44269 25783 44327 25789
rect 44450 25780 44456 25832
rect 44508 25820 44514 25832
rect 45278 25820 45284 25832
rect 44508 25792 45284 25820
rect 44508 25780 44514 25792
rect 45278 25780 45284 25792
rect 45336 25780 45342 25832
rect 46750 25820 46756 25832
rect 46711 25792 46756 25820
rect 46750 25780 46756 25792
rect 46808 25780 46814 25832
rect 47026 25820 47032 25832
rect 46987 25792 47032 25820
rect 47026 25780 47032 25792
rect 47084 25780 47090 25832
rect 47210 25820 47216 25832
rect 47171 25792 47216 25820
rect 47210 25780 47216 25792
rect 47268 25780 47274 25832
rect 38712 25724 39252 25752
rect 39393 25755 39451 25761
rect 38712 25712 38718 25724
rect 39393 25721 39405 25755
rect 39439 25721 39451 25755
rect 39393 25715 39451 25721
rect 20346 25684 20352 25696
rect 20088 25656 20352 25684
rect 20346 25644 20352 25656
rect 20404 25644 20410 25696
rect 26418 25684 26424 25696
rect 26379 25656 26424 25684
rect 26418 25644 26424 25656
rect 26476 25644 26482 25696
rect 29546 25684 29552 25696
rect 29507 25656 29552 25684
rect 29546 25644 29552 25656
rect 29604 25644 29610 25696
rect 30190 25644 30196 25696
rect 30248 25684 30254 25696
rect 33686 25684 33692 25696
rect 30248 25656 33692 25684
rect 30248 25644 30254 25656
rect 33686 25644 33692 25656
rect 33744 25644 33750 25696
rect 38286 25644 38292 25696
rect 38344 25684 38350 25696
rect 38381 25687 38439 25693
rect 38381 25684 38393 25687
rect 38344 25656 38393 25684
rect 38344 25644 38350 25656
rect 38381 25653 38393 25656
rect 38427 25653 38439 25687
rect 38381 25647 38439 25653
rect 47949 25687 48007 25693
rect 47949 25653 47961 25687
rect 47995 25684 48007 25687
rect 48314 25684 48320 25696
rect 47995 25656 48320 25684
rect 47995 25653 48007 25656
rect 47949 25647 48007 25653
rect 48314 25644 48320 25656
rect 48372 25644 48378 25696
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 6454 25480 6460 25492
rect 6415 25452 6460 25480
rect 6454 25440 6460 25452
rect 6512 25440 6518 25492
rect 7098 25480 7104 25492
rect 7059 25452 7104 25480
rect 7098 25440 7104 25452
rect 7156 25440 7162 25492
rect 11425 25483 11483 25489
rect 11425 25449 11437 25483
rect 11471 25480 11483 25483
rect 12250 25480 12256 25492
rect 11471 25452 12256 25480
rect 11471 25449 11483 25452
rect 11425 25443 11483 25449
rect 12250 25440 12256 25452
rect 12308 25440 12314 25492
rect 18598 25480 18604 25492
rect 18559 25452 18604 25480
rect 18598 25440 18604 25452
rect 18656 25440 18662 25492
rect 19518 25440 19524 25492
rect 19576 25480 19582 25492
rect 21545 25483 21603 25489
rect 21545 25480 21557 25483
rect 19576 25452 21557 25480
rect 19576 25440 19582 25452
rect 21545 25449 21557 25452
rect 21591 25449 21603 25483
rect 24946 25480 24952 25492
rect 24907 25452 24952 25480
rect 21545 25443 21603 25449
rect 24946 25440 24952 25452
rect 25004 25440 25010 25492
rect 28445 25483 28503 25489
rect 28445 25449 28457 25483
rect 28491 25480 28503 25483
rect 29638 25480 29644 25492
rect 28491 25452 29644 25480
rect 28491 25449 28503 25452
rect 28445 25443 28503 25449
rect 29638 25440 29644 25452
rect 29696 25440 29702 25492
rect 31202 25480 31208 25492
rect 31163 25452 31208 25480
rect 31202 25440 31208 25452
rect 31260 25440 31266 25492
rect 32217 25483 32275 25489
rect 32217 25449 32229 25483
rect 32263 25480 32275 25483
rect 32306 25480 32312 25492
rect 32263 25452 32312 25480
rect 32263 25449 32275 25452
rect 32217 25443 32275 25449
rect 32306 25440 32312 25452
rect 32364 25440 32370 25492
rect 32582 25440 32588 25492
rect 32640 25480 32646 25492
rect 33778 25480 33784 25492
rect 32640 25452 33784 25480
rect 32640 25440 32646 25452
rect 33778 25440 33784 25452
rect 33836 25440 33842 25492
rect 43070 25480 43076 25492
rect 43031 25452 43076 25480
rect 43070 25440 43076 25452
rect 43128 25440 43134 25492
rect 43530 25440 43536 25492
rect 43588 25480 43594 25492
rect 43901 25483 43959 25489
rect 43901 25480 43913 25483
rect 43588 25452 43913 25480
rect 43588 25440 43594 25452
rect 43901 25449 43913 25452
rect 43947 25449 43959 25483
rect 43901 25443 43959 25449
rect 44085 25483 44143 25489
rect 44085 25449 44097 25483
rect 44131 25480 44143 25483
rect 44450 25480 44456 25492
rect 44131 25452 44456 25480
rect 44131 25449 44143 25452
rect 44085 25443 44143 25449
rect 44450 25440 44456 25452
rect 44508 25440 44514 25492
rect 45186 25480 45192 25492
rect 45147 25452 45192 25480
rect 45186 25440 45192 25452
rect 45244 25440 45250 25492
rect 45373 25483 45431 25489
rect 45373 25449 45385 25483
rect 45419 25449 45431 25483
rect 45373 25443 45431 25449
rect 9306 25372 9312 25424
rect 9364 25412 9370 25424
rect 18506 25412 18512 25424
rect 9364 25384 9720 25412
rect 18467 25384 18512 25412
rect 9364 25372 9370 25384
rect 3418 25344 3424 25356
rect 3379 25316 3424 25344
rect 3418 25304 3424 25316
rect 3476 25304 3482 25356
rect 8018 25304 8024 25356
rect 8076 25344 8082 25356
rect 9582 25344 9588 25356
rect 8076 25316 8340 25344
rect 9543 25316 9588 25344
rect 8076 25304 8082 25316
rect 1578 25276 1584 25288
rect 1539 25248 1584 25276
rect 1578 25236 1584 25248
rect 1636 25236 1642 25288
rect 8312 25285 8340 25316
rect 9582 25304 9588 25316
rect 9640 25304 9646 25356
rect 9692 25353 9720 25384
rect 18506 25372 18512 25384
rect 18564 25372 18570 25424
rect 9677 25347 9735 25353
rect 9677 25313 9689 25347
rect 9723 25313 9735 25347
rect 9677 25307 9735 25313
rect 12526 25304 12532 25356
rect 12584 25344 12590 25356
rect 12805 25347 12863 25353
rect 12805 25344 12817 25347
rect 12584 25316 12817 25344
rect 12584 25304 12590 25316
rect 12805 25313 12817 25316
rect 12851 25313 12863 25347
rect 17034 25344 17040 25356
rect 16995 25316 17040 25344
rect 12805 25307 12863 25313
rect 17034 25304 17040 25316
rect 17092 25304 17098 25356
rect 19536 25344 19564 25440
rect 20990 25412 20996 25424
rect 20951 25384 20996 25412
rect 20990 25372 20996 25384
rect 21048 25372 21054 25424
rect 38378 25412 38384 25424
rect 30116 25384 38384 25412
rect 18708 25316 19564 25344
rect 6457 25279 6515 25285
rect 6457 25245 6469 25279
rect 6503 25245 6515 25279
rect 6457 25239 6515 25245
rect 7285 25279 7343 25285
rect 7285 25245 7297 25279
rect 7331 25276 7343 25279
rect 8297 25279 8355 25285
rect 7331 25248 8248 25276
rect 7331 25245 7343 25248
rect 7285 25239 7343 25245
rect 3234 25208 3240 25220
rect 3195 25180 3240 25208
rect 3234 25168 3240 25180
rect 3292 25168 3298 25220
rect 6472 25208 6500 25239
rect 8018 25208 8024 25220
rect 6472 25180 8024 25208
rect 8018 25168 8024 25180
rect 8076 25168 8082 25220
rect 8220 25140 8248 25248
rect 8297 25245 8309 25279
rect 8343 25245 8355 25279
rect 8297 25239 8355 25245
rect 9493 25279 9551 25285
rect 9493 25245 9505 25279
rect 9539 25276 9551 25279
rect 12621 25279 12679 25285
rect 12621 25276 12633 25279
rect 9539 25248 12633 25276
rect 9539 25245 9551 25248
rect 9493 25239 9551 25245
rect 12621 25245 12633 25248
rect 12667 25276 12679 25279
rect 13078 25276 13084 25288
rect 12667 25248 13084 25276
rect 12667 25245 12679 25248
rect 12621 25239 12679 25245
rect 13078 25236 13084 25248
rect 13136 25236 13142 25288
rect 15013 25279 15071 25285
rect 15013 25245 15025 25279
rect 15059 25276 15071 25279
rect 15286 25276 15292 25288
rect 15059 25248 15292 25276
rect 15059 25245 15071 25248
rect 15013 25239 15071 25245
rect 15286 25236 15292 25248
rect 15344 25236 15350 25288
rect 15930 25276 15936 25288
rect 15891 25248 15936 25276
rect 15930 25236 15936 25248
rect 15988 25236 15994 25288
rect 16206 25276 16212 25288
rect 16167 25248 16212 25276
rect 16206 25236 16212 25248
rect 16264 25236 16270 25288
rect 16301 25279 16359 25285
rect 16301 25245 16313 25279
rect 16347 25276 16359 25279
rect 16942 25276 16948 25288
rect 16347 25248 16948 25276
rect 16347 25245 16359 25248
rect 16301 25239 16359 25245
rect 16942 25236 16948 25248
rect 17000 25236 17006 25288
rect 17129 25279 17187 25285
rect 17129 25245 17141 25279
rect 17175 25276 17187 25279
rect 17862 25276 17868 25288
rect 17175 25248 17868 25276
rect 17175 25245 17187 25248
rect 17129 25239 17187 25245
rect 17862 25236 17868 25248
rect 17920 25276 17926 25288
rect 18708 25285 18736 25316
rect 19610 25304 19616 25356
rect 19668 25344 19674 25356
rect 20533 25347 20591 25353
rect 20533 25344 20545 25347
rect 19668 25316 20545 25344
rect 19668 25304 19674 25316
rect 20533 25313 20545 25316
rect 20579 25313 20591 25347
rect 20533 25307 20591 25313
rect 23753 25347 23811 25353
rect 23753 25313 23765 25347
rect 23799 25344 23811 25347
rect 23842 25344 23848 25356
rect 23799 25316 23848 25344
rect 23799 25313 23811 25316
rect 23753 25307 23811 25313
rect 23842 25304 23848 25316
rect 23900 25304 23906 25356
rect 25590 25344 25596 25356
rect 24044 25316 25596 25344
rect 18417 25279 18475 25285
rect 18417 25276 18429 25279
rect 17920 25248 18429 25276
rect 17920 25236 17926 25248
rect 18417 25245 18429 25248
rect 18463 25245 18475 25279
rect 18417 25239 18475 25245
rect 18693 25279 18751 25285
rect 18693 25245 18705 25279
rect 18739 25245 18751 25279
rect 18693 25239 18751 25245
rect 18874 25236 18880 25288
rect 18932 25276 18938 25288
rect 20622 25276 20628 25288
rect 18932 25248 20628 25276
rect 18932 25236 18938 25248
rect 20622 25236 20628 25248
rect 20680 25236 20686 25288
rect 21450 25276 21456 25288
rect 21411 25248 21456 25276
rect 21450 25236 21456 25248
rect 21508 25236 21514 25288
rect 21634 25276 21640 25288
rect 21595 25248 21640 25276
rect 21634 25236 21640 25248
rect 21692 25236 21698 25288
rect 23658 25276 23664 25288
rect 23619 25248 23664 25276
rect 23658 25236 23664 25248
rect 23716 25236 23722 25288
rect 8570 25208 8576 25220
rect 8531 25180 8576 25208
rect 8570 25168 8576 25180
rect 8628 25168 8634 25220
rect 11606 25208 11612 25220
rect 11567 25180 11612 25208
rect 11606 25168 11612 25180
rect 11664 25168 11670 25220
rect 11793 25211 11851 25217
rect 11793 25177 11805 25211
rect 11839 25208 11851 25211
rect 16114 25208 16120 25220
rect 11839 25180 12296 25208
rect 16075 25180 16120 25208
rect 11839 25177 11851 25180
rect 11793 25171 11851 25177
rect 12268 25149 12296 25180
rect 16114 25168 16120 25180
rect 16172 25168 16178 25220
rect 18230 25168 18236 25220
rect 18288 25208 18294 25220
rect 24044 25208 24072 25316
rect 25590 25304 25596 25316
rect 25648 25304 25654 25356
rect 24118 25236 24124 25288
rect 24176 25276 24182 25288
rect 25777 25279 25835 25285
rect 25777 25276 25789 25279
rect 24176 25248 25789 25276
rect 24176 25236 24182 25248
rect 25777 25245 25789 25248
rect 25823 25245 25835 25279
rect 25777 25239 25835 25245
rect 26044 25279 26102 25285
rect 26044 25245 26056 25279
rect 26090 25276 26102 25279
rect 26418 25276 26424 25288
rect 26090 25248 26424 25276
rect 26090 25245 26102 25248
rect 26044 25239 26102 25245
rect 26418 25236 26424 25248
rect 26476 25236 26482 25288
rect 28629 25279 28687 25285
rect 28629 25245 28641 25279
rect 28675 25245 28687 25279
rect 28629 25239 28687 25245
rect 18288 25180 24072 25208
rect 25133 25211 25191 25217
rect 18288 25168 18294 25180
rect 25133 25177 25145 25211
rect 25179 25177 25191 25211
rect 25133 25171 25191 25177
rect 25317 25211 25375 25217
rect 25317 25177 25329 25211
rect 25363 25208 25375 25211
rect 25866 25208 25872 25220
rect 25363 25180 25872 25208
rect 25363 25177 25375 25180
rect 25317 25171 25375 25177
rect 9125 25143 9183 25149
rect 9125 25140 9137 25143
rect 8220 25112 9137 25140
rect 9125 25109 9137 25112
rect 9171 25109 9183 25143
rect 9125 25103 9183 25109
rect 12253 25143 12311 25149
rect 12253 25109 12265 25143
rect 12299 25109 12311 25143
rect 12253 25103 12311 25109
rect 12618 25100 12624 25152
rect 12676 25140 12682 25152
rect 12713 25143 12771 25149
rect 12713 25140 12725 25143
rect 12676 25112 12725 25140
rect 12676 25100 12682 25112
rect 12713 25109 12725 25112
rect 12759 25109 12771 25143
rect 14826 25140 14832 25152
rect 14787 25112 14832 25140
rect 12713 25103 12771 25109
rect 14826 25100 14832 25112
rect 14884 25100 14890 25152
rect 16485 25143 16543 25149
rect 16485 25109 16497 25143
rect 16531 25140 16543 25143
rect 17310 25140 17316 25152
rect 16531 25112 17316 25140
rect 16531 25109 16543 25112
rect 16485 25103 16543 25109
rect 17310 25100 17316 25112
rect 17368 25100 17374 25152
rect 17494 25140 17500 25152
rect 17455 25112 17500 25140
rect 17494 25100 17500 25112
rect 17552 25100 17558 25152
rect 18138 25140 18144 25152
rect 18099 25112 18144 25140
rect 18138 25100 18144 25112
rect 18196 25100 18202 25152
rect 23293 25143 23351 25149
rect 23293 25109 23305 25143
rect 23339 25140 23351 25143
rect 23750 25140 23756 25152
rect 23339 25112 23756 25140
rect 23339 25109 23351 25112
rect 23293 25103 23351 25109
rect 23750 25100 23756 25112
rect 23808 25100 23814 25152
rect 25148 25140 25176 25171
rect 25866 25168 25872 25180
rect 25924 25208 25930 25220
rect 28644 25208 28672 25239
rect 29546 25236 29552 25288
rect 29604 25276 29610 25288
rect 30116 25285 30144 25384
rect 38378 25372 38384 25384
rect 38436 25372 38442 25424
rect 41782 25372 41788 25424
rect 41840 25412 41846 25424
rect 42061 25415 42119 25421
rect 42061 25412 42073 25415
rect 41840 25384 42073 25412
rect 41840 25372 41846 25384
rect 42061 25381 42073 25384
rect 42107 25381 42119 25415
rect 42061 25375 42119 25381
rect 43346 25372 43352 25424
rect 43404 25412 43410 25424
rect 45388 25412 45416 25443
rect 43404 25384 45416 25412
rect 43404 25372 43410 25384
rect 31665 25347 31723 25353
rect 31665 25344 31677 25347
rect 31496 25316 31677 25344
rect 30101 25279 30159 25285
rect 30101 25276 30113 25279
rect 29604 25248 30113 25276
rect 29604 25236 29610 25248
rect 30101 25245 30113 25248
rect 30147 25245 30159 25279
rect 30282 25276 30288 25288
rect 30243 25248 30288 25276
rect 30101 25239 30159 25245
rect 30282 25236 30288 25248
rect 30340 25236 30346 25288
rect 30561 25279 30619 25285
rect 30561 25245 30573 25279
rect 30607 25245 30619 25279
rect 30561 25239 30619 25245
rect 30745 25279 30803 25285
rect 30745 25245 30757 25279
rect 30791 25276 30803 25279
rect 31389 25279 31447 25285
rect 31389 25276 31401 25279
rect 30791 25248 31401 25276
rect 30791 25245 30803 25248
rect 30745 25239 30803 25245
rect 31389 25245 31401 25248
rect 31435 25245 31447 25279
rect 31389 25239 31447 25245
rect 25924 25180 28672 25208
rect 25924 25168 25930 25180
rect 26234 25140 26240 25152
rect 25148 25112 26240 25140
rect 26234 25100 26240 25112
rect 26292 25140 26298 25152
rect 27157 25143 27215 25149
rect 27157 25140 27169 25143
rect 26292 25112 27169 25140
rect 26292 25100 26298 25112
rect 27157 25109 27169 25112
rect 27203 25140 27215 25143
rect 27338 25140 27344 25152
rect 27203 25112 27344 25140
rect 27203 25109 27215 25112
rect 27157 25103 27215 25109
rect 27338 25100 27344 25112
rect 27396 25100 27402 25152
rect 28644 25140 28672 25180
rect 30190 25168 30196 25220
rect 30248 25208 30254 25220
rect 30576 25208 30604 25239
rect 30248 25180 30604 25208
rect 30248 25168 30254 25180
rect 30466 25140 30472 25152
rect 28644 25112 30472 25140
rect 30466 25100 30472 25112
rect 30524 25100 30530 25152
rect 30558 25100 30564 25152
rect 30616 25140 30622 25152
rect 31496 25140 31524 25316
rect 31665 25313 31677 25316
rect 31711 25313 31723 25347
rect 33505 25347 33563 25353
rect 33505 25344 33517 25347
rect 31665 25307 31723 25313
rect 32416 25316 33517 25344
rect 31570 25236 31576 25288
rect 31628 25276 31634 25288
rect 32416 25285 32444 25316
rect 33505 25313 33517 25316
rect 33551 25313 33563 25347
rect 43257 25347 43315 25353
rect 43257 25344 43269 25347
rect 33505 25307 33563 25313
rect 42444 25316 43269 25344
rect 32401 25279 32459 25285
rect 31628 25248 31754 25276
rect 31628 25236 31634 25248
rect 31726 25208 31754 25248
rect 32401 25245 32413 25279
rect 32447 25245 32459 25279
rect 32401 25239 32459 25245
rect 32585 25279 32643 25285
rect 32585 25245 32597 25279
rect 32631 25245 32643 25279
rect 32585 25239 32643 25245
rect 32600 25208 32628 25239
rect 32674 25236 32680 25288
rect 32732 25276 32738 25288
rect 33686 25276 33692 25288
rect 32732 25248 32777 25276
rect 33647 25248 33692 25276
rect 32732 25236 32738 25248
rect 33686 25236 33692 25248
rect 33744 25236 33750 25288
rect 33962 25276 33968 25288
rect 33923 25248 33968 25276
rect 33962 25236 33968 25248
rect 34020 25236 34026 25288
rect 34146 25276 34152 25288
rect 34107 25248 34152 25276
rect 34146 25236 34152 25248
rect 34204 25236 34210 25288
rect 40126 25276 40132 25288
rect 40087 25248 40132 25276
rect 40126 25236 40132 25248
rect 40184 25236 40190 25288
rect 42334 25276 42340 25288
rect 42295 25248 42340 25276
rect 42334 25236 42340 25248
rect 42392 25236 42398 25288
rect 40862 25208 40868 25220
rect 31726 25180 32628 25208
rect 40823 25180 40868 25208
rect 40862 25168 40868 25180
rect 40920 25168 40926 25220
rect 42058 25208 42064 25220
rect 42019 25180 42064 25208
rect 42058 25168 42064 25180
rect 42116 25168 42122 25220
rect 42444 25208 42472 25316
rect 43257 25313 43269 25316
rect 43303 25313 43315 25347
rect 46842 25344 46848 25356
rect 46803 25316 46848 25344
rect 43257 25307 43315 25313
rect 46842 25304 46848 25316
rect 46900 25304 46906 25356
rect 48130 25344 48136 25356
rect 48091 25316 48136 25344
rect 48130 25304 48136 25316
rect 48188 25304 48194 25356
rect 48314 25344 48320 25356
rect 48275 25316 48320 25344
rect 48314 25304 48320 25316
rect 48372 25304 48378 25356
rect 42886 25236 42892 25288
rect 42944 25276 42950 25288
rect 43073 25279 43131 25285
rect 43073 25276 43085 25279
rect 42944 25248 43085 25276
rect 42944 25236 42950 25248
rect 43073 25245 43085 25248
rect 43119 25245 43131 25279
rect 43438 25276 43444 25288
rect 43399 25248 43444 25276
rect 43073 25239 43131 25245
rect 43438 25236 43444 25248
rect 43496 25236 43502 25288
rect 43349 25211 43407 25217
rect 43349 25208 43361 25211
rect 42260 25180 42472 25208
rect 43088 25180 43361 25208
rect 39482 25140 39488 25152
rect 30616 25112 39488 25140
rect 30616 25100 30622 25112
rect 39482 25100 39488 25112
rect 39540 25100 39546 25152
rect 41414 25100 41420 25152
rect 41472 25140 41478 25152
rect 41966 25140 41972 25152
rect 41472 25112 41972 25140
rect 41472 25100 41478 25112
rect 41966 25100 41972 25112
rect 42024 25140 42030 25152
rect 42260 25149 42288 25180
rect 43088 25152 43116 25180
rect 43349 25177 43361 25180
rect 43395 25208 43407 25211
rect 44269 25211 44327 25217
rect 44269 25208 44281 25211
rect 43395 25180 44281 25208
rect 43395 25177 43407 25180
rect 43349 25171 43407 25177
rect 44269 25177 44281 25180
rect 44315 25208 44327 25211
rect 45554 25208 45560 25220
rect 44315 25180 45560 25208
rect 44315 25177 44327 25180
rect 44269 25171 44327 25177
rect 45554 25168 45560 25180
rect 45612 25168 45618 25220
rect 42245 25143 42303 25149
rect 42245 25140 42257 25143
rect 42024 25112 42257 25140
rect 42024 25100 42030 25112
rect 42245 25109 42257 25112
rect 42291 25109 42303 25143
rect 42245 25103 42303 25109
rect 43070 25100 43076 25152
rect 43128 25100 43134 25152
rect 43438 25100 43444 25152
rect 43496 25140 43502 25152
rect 44069 25143 44127 25149
rect 44069 25140 44081 25143
rect 43496 25112 44081 25140
rect 43496 25100 43502 25112
rect 44069 25109 44081 25112
rect 44115 25140 44127 25143
rect 45347 25143 45405 25149
rect 45347 25140 45359 25143
rect 44115 25112 45359 25140
rect 44115 25109 44127 25112
rect 44069 25103 44127 25109
rect 45347 25109 45359 25112
rect 45393 25109 45405 25143
rect 45347 25103 45405 25109
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 9493 24939 9551 24945
rect 9493 24905 9505 24939
rect 9539 24936 9551 24939
rect 9582 24936 9588 24948
rect 9539 24908 9588 24936
rect 9539 24905 9551 24908
rect 9493 24899 9551 24905
rect 9582 24896 9588 24908
rect 9640 24896 9646 24948
rect 11606 24896 11612 24948
rect 11664 24936 11670 24948
rect 13538 24936 13544 24948
rect 11664 24908 13544 24936
rect 11664 24896 11670 24908
rect 13538 24896 13544 24908
rect 13596 24936 13602 24948
rect 15749 24939 15807 24945
rect 13596 24908 13768 24936
rect 13596 24896 13602 24908
rect 10321 24871 10379 24877
rect 10321 24837 10333 24871
rect 10367 24868 10379 24871
rect 12434 24868 12440 24880
rect 10367 24840 11652 24868
rect 10367 24837 10379 24840
rect 10321 24831 10379 24837
rect 2590 24800 2596 24812
rect 2551 24772 2596 24800
rect 2590 24760 2596 24772
rect 2648 24800 2654 24812
rect 5258 24800 5264 24812
rect 2648 24772 5264 24800
rect 2648 24760 2654 24772
rect 5258 24760 5264 24772
rect 5316 24760 5322 24812
rect 7561 24803 7619 24809
rect 7561 24769 7573 24803
rect 7607 24800 7619 24803
rect 8018 24800 8024 24812
rect 7607 24772 8024 24800
rect 7607 24769 7619 24772
rect 7561 24763 7619 24769
rect 8018 24760 8024 24772
rect 8076 24760 8082 24812
rect 8380 24803 8438 24809
rect 8380 24769 8392 24803
rect 8426 24800 8438 24803
rect 8846 24800 8852 24812
rect 8426 24772 8852 24800
rect 8426 24769 8438 24772
rect 8380 24763 8438 24769
rect 8846 24760 8852 24772
rect 8904 24760 8910 24812
rect 10226 24800 10232 24812
rect 10187 24772 10232 24800
rect 10226 24760 10232 24772
rect 10284 24760 10290 24812
rect 2501 24735 2559 24741
rect 2501 24701 2513 24735
rect 2547 24732 2559 24735
rect 3234 24732 3240 24744
rect 2547 24704 3240 24732
rect 2547 24701 2559 24704
rect 2501 24695 2559 24701
rect 3234 24692 3240 24704
rect 3292 24692 3298 24744
rect 7653 24735 7711 24741
rect 7653 24701 7665 24735
rect 7699 24732 7711 24735
rect 8113 24735 8171 24741
rect 8113 24732 8125 24735
rect 7699 24704 8125 24732
rect 7699 24701 7711 24704
rect 7653 24695 7711 24701
rect 8113 24701 8125 24704
rect 8159 24701 8171 24735
rect 8113 24695 8171 24701
rect 9306 24692 9312 24744
rect 9364 24732 9370 24744
rect 10045 24735 10103 24741
rect 10045 24732 10057 24735
rect 9364 24704 10057 24732
rect 9364 24692 9370 24704
rect 10045 24701 10057 24704
rect 10091 24701 10103 24735
rect 10045 24695 10103 24701
rect 10689 24599 10747 24605
rect 10689 24565 10701 24599
rect 10735 24596 10747 24599
rect 11146 24596 11152 24608
rect 10735 24568 11152 24596
rect 10735 24565 10747 24568
rect 10689 24559 10747 24565
rect 11146 24556 11152 24568
rect 11204 24556 11210 24608
rect 11624 24596 11652 24840
rect 11716 24840 12440 24868
rect 11716 24809 11744 24840
rect 12434 24828 12440 24840
rect 12492 24868 12498 24880
rect 12492 24840 13676 24868
rect 12492 24828 12498 24840
rect 11701 24803 11759 24809
rect 11701 24769 11713 24803
rect 11747 24769 11759 24803
rect 11701 24763 11759 24769
rect 11790 24760 11796 24812
rect 11848 24800 11854 24812
rect 11957 24803 12015 24809
rect 11957 24800 11969 24803
rect 11848 24772 11969 24800
rect 11848 24760 11854 24772
rect 11957 24769 11969 24772
rect 12003 24769 12015 24803
rect 11957 24763 12015 24769
rect 12986 24760 12992 24812
rect 13044 24800 13050 24812
rect 13541 24803 13599 24809
rect 13541 24800 13553 24803
rect 13044 24772 13553 24800
rect 13044 24760 13050 24772
rect 13541 24769 13553 24772
rect 13587 24769 13599 24803
rect 13541 24763 13599 24769
rect 13648 24744 13676 24840
rect 13740 24809 13768 24908
rect 15749 24905 15761 24939
rect 15795 24936 15807 24939
rect 16114 24936 16120 24948
rect 15795 24908 16120 24936
rect 15795 24905 15807 24908
rect 15749 24899 15807 24905
rect 16114 24896 16120 24908
rect 16172 24936 16178 24948
rect 17862 24936 17868 24948
rect 16172 24908 16574 24936
rect 17823 24908 17868 24936
rect 16172 24896 16178 24908
rect 14636 24871 14694 24877
rect 14636 24837 14648 24871
rect 14682 24868 14694 24871
rect 14826 24868 14832 24880
rect 14682 24840 14832 24868
rect 14682 24837 14694 24840
rect 14636 24831 14694 24837
rect 14826 24828 14832 24840
rect 14884 24828 14890 24880
rect 13725 24803 13783 24809
rect 13725 24769 13737 24803
rect 13771 24769 13783 24803
rect 16546 24800 16574 24908
rect 17862 24896 17868 24908
rect 17920 24896 17926 24948
rect 20622 24896 20628 24948
rect 20680 24936 20686 24948
rect 23385 24939 23443 24945
rect 23385 24936 23397 24939
rect 20680 24908 23397 24936
rect 20680 24896 20686 24908
rect 23385 24905 23397 24908
rect 23431 24905 23443 24939
rect 27338 24936 27344 24948
rect 27299 24908 27344 24936
rect 23385 24899 23443 24905
rect 27338 24896 27344 24908
rect 27396 24896 27402 24948
rect 30282 24896 30288 24948
rect 30340 24936 30346 24948
rect 32585 24939 32643 24945
rect 30340 24908 31754 24936
rect 30340 24896 30346 24908
rect 24854 24828 24860 24880
rect 24912 24868 24918 24880
rect 25225 24871 25283 24877
rect 25225 24868 25237 24871
rect 24912 24840 25237 24868
rect 24912 24828 24918 24840
rect 25225 24837 25237 24840
rect 25271 24837 25283 24871
rect 25225 24831 25283 24837
rect 16853 24803 16911 24809
rect 16853 24800 16865 24803
rect 16546 24772 16865 24800
rect 13725 24763 13783 24769
rect 16853 24769 16865 24772
rect 16899 24769 16911 24803
rect 16853 24763 16911 24769
rect 17037 24803 17095 24809
rect 17037 24769 17049 24803
rect 17083 24769 17095 24803
rect 17678 24800 17684 24812
rect 17639 24772 17684 24800
rect 17037 24763 17095 24769
rect 13630 24692 13636 24744
rect 13688 24732 13694 24744
rect 14369 24735 14427 24741
rect 14369 24732 14381 24735
rect 13688 24704 14381 24732
rect 13688 24692 13694 24704
rect 14369 24701 14381 24704
rect 14415 24701 14427 24735
rect 14369 24695 14427 24701
rect 16482 24692 16488 24744
rect 16540 24732 16546 24744
rect 17052 24732 17080 24763
rect 17678 24760 17684 24772
rect 17736 24760 17742 24812
rect 17865 24803 17923 24809
rect 17865 24769 17877 24803
rect 17911 24800 17923 24803
rect 18325 24803 18383 24809
rect 18325 24800 18337 24803
rect 17911 24772 18337 24800
rect 17911 24769 17923 24772
rect 17865 24763 17923 24769
rect 18325 24769 18337 24772
rect 18371 24769 18383 24803
rect 18325 24763 18383 24769
rect 18509 24803 18567 24809
rect 18509 24769 18521 24803
rect 18555 24769 18567 24803
rect 18509 24763 18567 24769
rect 16540 24704 17080 24732
rect 17221 24735 17279 24741
rect 16540 24692 16546 24704
rect 17221 24701 17233 24735
rect 17267 24732 17279 24735
rect 17880 24732 17908 24763
rect 17267 24704 17908 24732
rect 17267 24701 17279 24704
rect 17221 24695 17279 24701
rect 17310 24624 17316 24676
rect 17368 24664 17374 24676
rect 18524 24664 18552 24763
rect 19610 24760 19616 24812
rect 19668 24800 19674 24812
rect 19705 24803 19763 24809
rect 19705 24800 19717 24803
rect 19668 24772 19717 24800
rect 19668 24760 19674 24772
rect 19705 24769 19717 24772
rect 19751 24769 19763 24803
rect 22189 24803 22247 24809
rect 22189 24800 22201 24803
rect 19705 24763 19763 24769
rect 19904 24772 22201 24800
rect 19058 24692 19064 24744
rect 19116 24732 19122 24744
rect 19904 24732 19932 24772
rect 22189 24769 22201 24772
rect 22235 24800 22247 24803
rect 23474 24800 23480 24812
rect 22235 24772 23480 24800
rect 22235 24769 22247 24772
rect 22189 24763 22247 24769
rect 23474 24760 23480 24772
rect 23532 24760 23538 24812
rect 23566 24760 23572 24812
rect 23624 24800 23630 24812
rect 23661 24803 23719 24809
rect 23661 24800 23673 24803
rect 23624 24772 23673 24800
rect 23624 24760 23630 24772
rect 23661 24769 23673 24772
rect 23707 24769 23719 24803
rect 25866 24800 25872 24812
rect 25827 24772 25872 24800
rect 23661 24763 23719 24769
rect 25866 24760 25872 24772
rect 25924 24760 25930 24812
rect 26234 24800 26240 24812
rect 26195 24772 26240 24800
rect 26234 24760 26240 24772
rect 26292 24760 26298 24812
rect 27157 24803 27215 24809
rect 27157 24800 27169 24803
rect 26344 24772 27169 24800
rect 19116 24704 19932 24732
rect 19116 24692 19122 24704
rect 19978 24692 19984 24744
rect 20036 24732 20042 24744
rect 23106 24732 23112 24744
rect 20036 24704 22968 24732
rect 23067 24704 23112 24732
rect 20036 24692 20042 24704
rect 17368 24636 18552 24664
rect 17368 24624 17374 24636
rect 12342 24596 12348 24608
rect 11624 24568 12348 24596
rect 12342 24556 12348 24568
rect 12400 24596 12406 24608
rect 13081 24599 13139 24605
rect 13081 24596 13093 24599
rect 12400 24568 13093 24596
rect 12400 24556 12406 24568
rect 13081 24565 13093 24568
rect 13127 24565 13139 24599
rect 13906 24596 13912 24608
rect 13867 24568 13912 24596
rect 13081 24559 13139 24565
rect 13906 24556 13912 24568
rect 13964 24556 13970 24608
rect 17862 24556 17868 24608
rect 17920 24596 17926 24608
rect 18417 24599 18475 24605
rect 18417 24596 18429 24599
rect 17920 24568 18429 24596
rect 17920 24556 17926 24568
rect 18417 24565 18429 24568
rect 18463 24565 18475 24599
rect 18417 24559 18475 24565
rect 19334 24556 19340 24608
rect 19392 24596 19398 24608
rect 19521 24599 19579 24605
rect 19521 24596 19533 24599
rect 19392 24568 19533 24596
rect 19392 24556 19398 24568
rect 19521 24565 19533 24568
rect 19567 24565 19579 24599
rect 19521 24559 19579 24565
rect 19889 24599 19947 24605
rect 19889 24565 19901 24599
rect 19935 24596 19947 24599
rect 20438 24596 20444 24608
rect 19935 24568 20444 24596
rect 19935 24565 19947 24568
rect 19889 24559 19947 24565
rect 20438 24556 20444 24568
rect 20496 24556 20502 24608
rect 22002 24556 22008 24608
rect 22060 24596 22066 24608
rect 22097 24599 22155 24605
rect 22097 24596 22109 24599
rect 22060 24568 22109 24596
rect 22060 24556 22066 24568
rect 22097 24565 22109 24568
rect 22143 24565 22155 24599
rect 22940 24596 22968 24704
rect 23106 24692 23112 24704
rect 23164 24692 23170 24744
rect 23753 24735 23811 24741
rect 23753 24701 23765 24735
rect 23799 24732 23811 24735
rect 23842 24732 23848 24744
rect 23799 24704 23848 24732
rect 23799 24701 23811 24704
rect 23753 24695 23811 24701
rect 23842 24692 23848 24704
rect 23900 24692 23906 24744
rect 26142 24624 26148 24676
rect 26200 24664 26206 24676
rect 26344 24664 26372 24772
rect 27157 24769 27169 24772
rect 27203 24769 27215 24803
rect 27157 24763 27215 24769
rect 27430 24760 27436 24812
rect 27488 24800 27494 24812
rect 30285 24803 30343 24809
rect 27488 24772 27533 24800
rect 27488 24760 27494 24772
rect 30285 24769 30297 24803
rect 30331 24769 30343 24803
rect 30742 24800 30748 24812
rect 30703 24772 30748 24800
rect 30285 24763 30343 24769
rect 27154 24664 27160 24676
rect 26200 24636 26372 24664
rect 27115 24636 27160 24664
rect 26200 24624 26206 24636
rect 27154 24624 27160 24636
rect 27212 24624 27218 24676
rect 28994 24664 29000 24676
rect 28955 24636 29000 24664
rect 28994 24624 29000 24636
rect 29052 24624 29058 24676
rect 30300 24664 30328 24763
rect 30742 24760 30748 24772
rect 30800 24760 30806 24812
rect 30929 24803 30987 24809
rect 30929 24769 30941 24803
rect 30975 24800 30987 24803
rect 31018 24800 31024 24812
rect 30975 24772 31024 24800
rect 30975 24769 30987 24772
rect 30929 24763 30987 24769
rect 31018 24760 31024 24772
rect 31076 24760 31082 24812
rect 31202 24800 31208 24812
rect 31163 24772 31208 24800
rect 31202 24760 31208 24772
rect 31260 24760 31266 24812
rect 31404 24809 31432 24908
rect 31726 24868 31754 24908
rect 32585 24905 32597 24939
rect 32631 24936 32643 24939
rect 32766 24936 32772 24948
rect 32631 24908 32772 24936
rect 32631 24905 32643 24908
rect 32585 24899 32643 24905
rect 32766 24896 32772 24908
rect 32824 24936 32830 24948
rect 36446 24936 36452 24948
rect 32824 24908 36452 24936
rect 32824 24896 32830 24908
rect 36446 24896 36452 24908
rect 36504 24896 36510 24948
rect 41966 24936 41972 24948
rect 41927 24908 41972 24936
rect 41966 24896 41972 24908
rect 42024 24896 42030 24948
rect 45554 24896 45560 24948
rect 45612 24936 45618 24948
rect 45649 24939 45707 24945
rect 45649 24936 45661 24939
rect 45612 24908 45661 24936
rect 45612 24896 45618 24908
rect 45649 24905 45661 24908
rect 45695 24905 45707 24939
rect 45649 24899 45707 24905
rect 33502 24868 33508 24880
rect 31726 24840 33508 24868
rect 33502 24828 33508 24840
rect 33560 24868 33566 24880
rect 33962 24868 33968 24880
rect 33560 24840 33968 24868
rect 33560 24828 33566 24840
rect 33962 24828 33968 24840
rect 34020 24828 34026 24880
rect 43530 24868 43536 24880
rect 38672 24840 41414 24868
rect 38672 24812 38700 24840
rect 31389 24803 31447 24809
rect 31389 24769 31401 24803
rect 31435 24769 31447 24803
rect 31389 24763 31447 24769
rect 31478 24760 31484 24812
rect 31536 24800 31542 24812
rect 32309 24803 32367 24809
rect 32309 24800 32321 24803
rect 31536 24772 32321 24800
rect 31536 24760 31542 24772
rect 32309 24769 32321 24772
rect 32355 24769 32367 24803
rect 32309 24763 32367 24769
rect 32769 24803 32827 24809
rect 32769 24769 32781 24803
rect 32815 24769 32827 24803
rect 32769 24763 32827 24769
rect 30466 24692 30472 24744
rect 30524 24732 30530 24744
rect 32784 24732 32812 24763
rect 32858 24760 32864 24812
rect 32916 24800 32922 24812
rect 33594 24800 33600 24812
rect 32916 24772 33180 24800
rect 33555 24772 33600 24800
rect 32916 24760 32922 24772
rect 30524 24704 32812 24732
rect 33152 24732 33180 24772
rect 33594 24760 33600 24772
rect 33652 24760 33658 24812
rect 33778 24800 33784 24812
rect 33739 24772 33784 24800
rect 33778 24760 33784 24772
rect 33836 24760 33842 24812
rect 34057 24803 34115 24809
rect 34057 24769 34069 24803
rect 34103 24800 34115 24803
rect 37734 24800 37740 24812
rect 34103 24772 37740 24800
rect 34103 24769 34115 24772
rect 34057 24763 34115 24769
rect 34072 24732 34100 24763
rect 37734 24760 37740 24772
rect 37792 24760 37798 24812
rect 38654 24800 38660 24812
rect 38028 24772 38660 24800
rect 33152 24704 34100 24732
rect 30524 24692 30530 24704
rect 34146 24692 34152 24744
rect 34204 24732 34210 24744
rect 38028 24732 38056 24772
rect 38654 24760 38660 24772
rect 38712 24760 38718 24812
rect 38838 24760 38844 24812
rect 38896 24800 38902 24812
rect 39025 24803 39083 24809
rect 39025 24800 39037 24803
rect 38896 24772 39037 24800
rect 38896 24760 38902 24772
rect 39025 24769 39037 24772
rect 39071 24769 39083 24803
rect 39025 24763 39083 24769
rect 34204 24704 38056 24732
rect 34204 24692 34210 24704
rect 38102 24692 38108 24744
rect 38160 24732 38166 24744
rect 38562 24732 38568 24744
rect 38160 24704 38568 24732
rect 38160 24692 38166 24704
rect 38562 24692 38568 24704
rect 38620 24732 38626 24744
rect 38749 24735 38807 24741
rect 38749 24732 38761 24735
rect 38620 24704 38761 24732
rect 38620 24692 38626 24704
rect 38749 24701 38761 24704
rect 38795 24701 38807 24735
rect 41386 24732 41414 24840
rect 43088 24840 43536 24868
rect 41782 24800 41788 24812
rect 41743 24772 41788 24800
rect 41782 24760 41788 24772
rect 41840 24760 41846 24812
rect 42061 24803 42119 24809
rect 42061 24769 42073 24803
rect 42107 24800 42119 24803
rect 43088 24800 43116 24840
rect 43530 24828 43536 24840
rect 43588 24828 43594 24880
rect 42107 24772 43116 24800
rect 42107 24769 42119 24772
rect 42061 24763 42119 24769
rect 43162 24760 43168 24812
rect 43220 24800 43226 24812
rect 43220 24772 43264 24800
rect 43220 24760 43226 24772
rect 43438 24760 43444 24812
rect 43496 24800 43502 24812
rect 44542 24809 44548 24812
rect 44269 24803 44327 24809
rect 44269 24800 44281 24803
rect 43496 24772 44281 24800
rect 43496 24760 43502 24772
rect 44269 24769 44281 24772
rect 44315 24769 44327 24803
rect 44269 24763 44327 24769
rect 44536 24763 44548 24809
rect 44600 24800 44606 24812
rect 46385 24803 46443 24809
rect 44600 24772 44636 24800
rect 44542 24760 44548 24763
rect 44600 24760 44606 24772
rect 46385 24769 46397 24803
rect 46431 24769 46443 24803
rect 46385 24763 46443 24769
rect 46477 24803 46535 24809
rect 46477 24769 46489 24803
rect 46523 24800 46535 24803
rect 47026 24800 47032 24812
rect 46523 24772 47032 24800
rect 46523 24769 46535 24772
rect 46477 24763 46535 24769
rect 41693 24735 41751 24741
rect 41693 24732 41705 24735
rect 41386 24704 41705 24732
rect 38749 24695 38807 24701
rect 41693 24701 41705 24704
rect 41739 24732 41751 24735
rect 42886 24732 42892 24744
rect 41739 24704 42892 24732
rect 41739 24701 41751 24704
rect 41693 24695 41751 24701
rect 42886 24692 42892 24704
rect 42944 24692 42950 24744
rect 43070 24732 43076 24744
rect 43031 24704 43076 24732
rect 43070 24692 43076 24704
rect 43128 24692 43134 24744
rect 43254 24732 43260 24744
rect 43215 24704 43260 24732
rect 43254 24692 43260 24704
rect 43312 24692 43318 24744
rect 43346 24692 43352 24744
rect 43404 24732 43410 24744
rect 46400 24732 46428 24763
rect 47026 24760 47032 24772
rect 47084 24760 47090 24812
rect 47210 24800 47216 24812
rect 47171 24772 47216 24800
rect 47210 24760 47216 24772
rect 47268 24760 47274 24812
rect 48222 24800 48228 24812
rect 48183 24772 48228 24800
rect 48222 24760 48228 24772
rect 48280 24760 48286 24812
rect 47486 24732 47492 24744
rect 43404 24704 43449 24732
rect 46400 24704 47492 24732
rect 43404 24692 43410 24704
rect 47228 24676 47256 24704
rect 47486 24692 47492 24704
rect 47544 24692 47550 24744
rect 30300 24636 44312 24664
rect 31754 24596 31760 24608
rect 22940 24568 31760 24596
rect 22097 24559 22155 24565
rect 31754 24556 31760 24568
rect 31812 24556 31818 24608
rect 31846 24556 31852 24608
rect 31904 24596 31910 24608
rect 33226 24596 33232 24608
rect 31904 24568 33232 24596
rect 31904 24556 31910 24568
rect 33226 24556 33232 24568
rect 33284 24596 33290 24608
rect 34146 24596 34152 24608
rect 33284 24568 34152 24596
rect 33284 24556 33290 24568
rect 34146 24556 34152 24568
rect 34204 24556 34210 24608
rect 34241 24599 34299 24605
rect 34241 24565 34253 24599
rect 34287 24596 34299 24599
rect 34698 24596 34704 24608
rect 34287 24568 34704 24596
rect 34287 24565 34299 24568
rect 34241 24559 34299 24565
rect 34698 24556 34704 24568
rect 34756 24556 34762 24608
rect 36446 24556 36452 24608
rect 36504 24596 36510 24608
rect 37826 24596 37832 24608
rect 36504 24568 37832 24596
rect 36504 24556 36510 24568
rect 37826 24556 37832 24568
rect 37884 24556 37890 24608
rect 38654 24556 38660 24608
rect 38712 24596 38718 24608
rect 38841 24599 38899 24605
rect 38841 24596 38853 24599
rect 38712 24568 38853 24596
rect 38712 24556 38718 24568
rect 38841 24565 38853 24568
rect 38887 24565 38899 24599
rect 39206 24596 39212 24608
rect 39167 24568 39212 24596
rect 38841 24559 38899 24565
rect 39206 24556 39212 24568
rect 39264 24556 39270 24608
rect 41598 24596 41604 24608
rect 41559 24568 41604 24596
rect 41598 24556 41604 24568
rect 41656 24556 41662 24608
rect 42702 24556 42708 24608
rect 42760 24596 42766 24608
rect 43438 24596 43444 24608
rect 42760 24568 43444 24596
rect 42760 24556 42766 24568
rect 43438 24556 43444 24568
rect 43496 24556 43502 24608
rect 43533 24599 43591 24605
rect 43533 24565 43545 24599
rect 43579 24596 43591 24599
rect 44174 24596 44180 24608
rect 43579 24568 44180 24596
rect 43579 24565 43591 24568
rect 43533 24559 43591 24565
rect 44174 24556 44180 24568
rect 44232 24556 44238 24608
rect 44284 24596 44312 24636
rect 47210 24624 47216 24676
rect 47268 24624 47274 24676
rect 48038 24664 48044 24676
rect 47999 24636 48044 24664
rect 48038 24624 48044 24636
rect 48096 24624 48102 24676
rect 45554 24596 45560 24608
rect 44284 24568 45560 24596
rect 45554 24556 45560 24568
rect 45612 24556 45618 24608
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 11790 24392 11796 24404
rect 11751 24364 11796 24392
rect 11790 24352 11796 24364
rect 11848 24352 11854 24404
rect 12986 24392 12992 24404
rect 12947 24364 12992 24392
rect 12986 24352 12992 24364
rect 13044 24352 13050 24404
rect 16666 24392 16672 24404
rect 13096 24364 16672 24392
rect 13096 24324 13124 24364
rect 16666 24352 16672 24364
rect 16724 24352 16730 24404
rect 16761 24395 16819 24401
rect 16761 24361 16773 24395
rect 16807 24392 16819 24395
rect 17678 24392 17684 24404
rect 16807 24364 17684 24392
rect 16807 24361 16819 24364
rect 16761 24355 16819 24361
rect 17678 24352 17684 24364
rect 17736 24352 17742 24404
rect 19610 24392 19616 24404
rect 19571 24364 19616 24392
rect 19610 24352 19616 24364
rect 19668 24352 19674 24404
rect 20070 24352 20076 24404
rect 20128 24392 20134 24404
rect 23014 24392 23020 24404
rect 20128 24364 23020 24392
rect 20128 24352 20134 24364
rect 23014 24352 23020 24364
rect 23072 24392 23078 24404
rect 26142 24392 26148 24404
rect 23072 24364 26148 24392
rect 23072 24352 23078 24364
rect 26142 24352 26148 24364
rect 26200 24352 26206 24404
rect 27157 24395 27215 24401
rect 27157 24361 27169 24395
rect 27203 24392 27215 24395
rect 27430 24392 27436 24404
rect 27203 24364 27436 24392
rect 27203 24361 27215 24364
rect 27157 24355 27215 24361
rect 27430 24352 27436 24364
rect 27488 24352 27494 24404
rect 27816 24364 28764 24392
rect 10980 24296 13124 24324
rect 8570 24216 8576 24268
rect 8628 24256 8634 24268
rect 9125 24259 9183 24265
rect 9125 24256 9137 24259
rect 8628 24228 9137 24256
rect 8628 24216 8634 24228
rect 9125 24225 9137 24228
rect 9171 24225 9183 24259
rect 9125 24219 9183 24225
rect 8202 24148 8208 24200
rect 8260 24188 8266 24200
rect 10980 24188 11008 24296
rect 14550 24284 14556 24336
rect 14608 24324 14614 24336
rect 14608 24296 15332 24324
rect 14608 24284 14614 24296
rect 12434 24256 12440 24268
rect 12395 24228 12440 24256
rect 12434 24216 12440 24228
rect 12492 24216 12498 24268
rect 12529 24259 12587 24265
rect 12529 24225 12541 24259
rect 12575 24256 12587 24259
rect 14734 24256 14740 24268
rect 12575 24228 14740 24256
rect 12575 24225 12587 24228
rect 12529 24219 12587 24225
rect 14734 24216 14740 24228
rect 14792 24216 14798 24268
rect 15304 24256 15332 24296
rect 15378 24284 15384 24336
rect 15436 24324 15442 24336
rect 15930 24324 15936 24336
rect 15436 24296 15936 24324
rect 15436 24284 15442 24296
rect 15930 24284 15936 24296
rect 15988 24324 15994 24336
rect 16482 24324 16488 24336
rect 15988 24296 16488 24324
rect 15988 24284 15994 24296
rect 16482 24284 16488 24296
rect 16540 24324 16546 24336
rect 16540 24296 16896 24324
rect 16540 24284 16546 24296
rect 16025 24259 16083 24265
rect 15304 24228 15608 24256
rect 11146 24188 11152 24200
rect 8260 24160 11008 24188
rect 11107 24160 11152 24188
rect 8260 24148 8266 24160
rect 11146 24148 11152 24160
rect 11204 24148 11210 24200
rect 11609 24191 11667 24197
rect 11609 24157 11621 24191
rect 11655 24188 11667 24191
rect 13906 24188 13912 24200
rect 11655 24160 13912 24188
rect 11655 24157 11667 24160
rect 11609 24151 11667 24157
rect 13906 24148 13912 24160
rect 13964 24148 13970 24200
rect 14550 24188 14556 24200
rect 14511 24160 14556 24188
rect 14550 24148 14556 24160
rect 14608 24148 14614 24200
rect 14829 24191 14887 24197
rect 14829 24157 14841 24191
rect 14875 24188 14887 24191
rect 14918 24188 14924 24200
rect 14875 24160 14924 24188
rect 14875 24157 14887 24160
rect 14829 24151 14887 24157
rect 14918 24148 14924 24160
rect 14976 24148 14982 24200
rect 15013 24191 15071 24197
rect 15013 24157 15025 24191
rect 15059 24188 15071 24191
rect 15378 24188 15384 24200
rect 15059 24160 15384 24188
rect 15059 24157 15071 24160
rect 15013 24151 15071 24157
rect 15378 24148 15384 24160
rect 15436 24148 15442 24200
rect 3326 24080 3332 24132
rect 3384 24120 3390 24132
rect 6365 24123 6423 24129
rect 6365 24120 6377 24123
rect 3384 24092 6377 24120
rect 3384 24080 3390 24092
rect 6365 24089 6377 24092
rect 6411 24089 6423 24123
rect 6365 24083 6423 24089
rect 6638 24080 6644 24132
rect 6696 24120 6702 24132
rect 8021 24123 8079 24129
rect 8021 24120 8033 24123
rect 6696 24092 8033 24120
rect 6696 24080 6702 24092
rect 8021 24089 8033 24092
rect 8067 24089 8079 24123
rect 8021 24083 8079 24089
rect 9392 24123 9450 24129
rect 9392 24089 9404 24123
rect 9438 24120 9450 24123
rect 9438 24092 11008 24120
rect 9438 24089 9450 24092
rect 9392 24083 9450 24089
rect 10134 24012 10140 24064
rect 10192 24052 10198 24064
rect 10980 24061 11008 24092
rect 12342 24080 12348 24132
rect 12400 24120 12406 24132
rect 12621 24123 12679 24129
rect 12621 24120 12633 24123
rect 12400 24092 12633 24120
rect 12400 24080 12406 24092
rect 12621 24089 12633 24092
rect 12667 24089 12679 24123
rect 12621 24083 12679 24089
rect 15286 24080 15292 24132
rect 15344 24120 15350 24132
rect 15344 24092 15516 24120
rect 15344 24080 15350 24092
rect 10505 24055 10563 24061
rect 10505 24052 10517 24055
rect 10192 24024 10517 24052
rect 10192 24012 10198 24024
rect 10505 24021 10517 24024
rect 10551 24021 10563 24055
rect 10505 24015 10563 24021
rect 10965 24055 11023 24061
rect 10965 24021 10977 24055
rect 11011 24021 11023 24055
rect 10965 24015 11023 24021
rect 14369 24055 14427 24061
rect 14369 24021 14381 24055
rect 14415 24052 14427 24055
rect 14458 24052 14464 24064
rect 14415 24024 14464 24052
rect 14415 24021 14427 24024
rect 14369 24015 14427 24021
rect 14458 24012 14464 24024
rect 14516 24012 14522 24064
rect 15488 24061 15516 24092
rect 15473 24055 15531 24061
rect 15473 24021 15485 24055
rect 15519 24021 15531 24055
rect 15580 24052 15608 24228
rect 16025 24225 16037 24259
rect 16071 24256 16083 24259
rect 16390 24256 16396 24268
rect 16071 24228 16396 24256
rect 16071 24225 16083 24228
rect 16025 24219 16083 24225
rect 16390 24216 16396 24228
rect 16448 24216 16454 24268
rect 15933 24191 15991 24197
rect 15933 24157 15945 24191
rect 15979 24188 15991 24191
rect 16114 24188 16120 24200
rect 15979 24160 16120 24188
rect 15979 24157 15991 24160
rect 15933 24151 15991 24157
rect 16114 24148 16120 24160
rect 16172 24188 16178 24200
rect 16868 24197 16896 24296
rect 16942 24284 16948 24336
rect 17000 24324 17006 24336
rect 17000 24296 26464 24324
rect 17000 24284 17006 24296
rect 17494 24216 17500 24268
rect 17552 24256 17558 24268
rect 17773 24259 17831 24265
rect 17773 24256 17785 24259
rect 17552 24228 17785 24256
rect 17552 24216 17558 24228
rect 17773 24225 17785 24228
rect 17819 24225 17831 24259
rect 17773 24219 17831 24225
rect 17865 24259 17923 24265
rect 17865 24225 17877 24259
rect 17911 24256 17923 24259
rect 21358 24256 21364 24268
rect 17911 24228 21364 24256
rect 17911 24225 17923 24228
rect 17865 24219 17923 24225
rect 16669 24191 16727 24197
rect 16669 24188 16681 24191
rect 16172 24160 16681 24188
rect 16172 24148 16178 24160
rect 16669 24157 16681 24160
rect 16715 24157 16727 24191
rect 16669 24151 16727 24157
rect 16853 24191 16911 24197
rect 16853 24157 16865 24191
rect 16899 24157 16911 24191
rect 16853 24151 16911 24157
rect 17586 24148 17592 24200
rect 17644 24188 17650 24200
rect 17880 24188 17908 24219
rect 21358 24216 21364 24228
rect 21416 24216 21422 24268
rect 21836 24265 21864 24296
rect 21821 24259 21879 24265
rect 21821 24225 21833 24259
rect 21867 24225 21879 24259
rect 22002 24256 22008 24268
rect 21963 24228 22008 24256
rect 21821 24219 21879 24225
rect 22002 24216 22008 24228
rect 22060 24216 22066 24268
rect 22830 24256 22836 24268
rect 22791 24228 22836 24256
rect 22830 24216 22836 24228
rect 22888 24216 22894 24268
rect 19794 24188 19800 24200
rect 17644 24160 17908 24188
rect 19755 24160 19800 24188
rect 17644 24148 17650 24160
rect 19794 24148 19800 24160
rect 19852 24148 19858 24200
rect 20070 24188 20076 24200
rect 20031 24160 20076 24188
rect 20070 24148 20076 24160
rect 20128 24148 20134 24200
rect 20257 24191 20315 24197
rect 20257 24157 20269 24191
rect 20303 24157 20315 24191
rect 20257 24151 20315 24157
rect 25685 24191 25743 24197
rect 25685 24157 25697 24191
rect 25731 24188 25743 24191
rect 25866 24188 25872 24200
rect 25731 24160 25872 24188
rect 25731 24157 25743 24160
rect 25685 24151 25743 24157
rect 15841 24123 15899 24129
rect 15841 24089 15853 24123
rect 15887 24120 15899 24123
rect 17681 24123 17739 24129
rect 15887 24092 17356 24120
rect 15887 24089 15899 24092
rect 15841 24083 15899 24089
rect 17126 24052 17132 24064
rect 15580 24024 17132 24052
rect 15473 24015 15531 24021
rect 17126 24012 17132 24024
rect 17184 24012 17190 24064
rect 17328 24061 17356 24092
rect 17681 24089 17693 24123
rect 17727 24120 17739 24123
rect 20272 24120 20300 24151
rect 25866 24148 25872 24160
rect 25924 24148 25930 24200
rect 20622 24120 20628 24132
rect 17727 24092 20628 24120
rect 17727 24089 17739 24092
rect 17681 24083 17739 24089
rect 20622 24080 20628 24092
rect 20680 24080 20686 24132
rect 26436 24120 26464 24296
rect 26605 24259 26663 24265
rect 26605 24225 26617 24259
rect 26651 24256 26663 24259
rect 27614 24256 27620 24268
rect 26651 24228 27620 24256
rect 26651 24225 26663 24228
rect 26605 24219 26663 24225
rect 27614 24216 27620 24228
rect 27672 24216 27678 24268
rect 26786 24188 26792 24200
rect 26699 24160 26792 24188
rect 26786 24148 26792 24160
rect 26844 24188 26850 24200
rect 27816 24188 27844 24364
rect 26844 24160 27844 24188
rect 27908 24228 28672 24256
rect 26844 24148 26850 24160
rect 26436 24092 26832 24120
rect 17313 24055 17371 24061
rect 17313 24021 17325 24055
rect 17359 24021 17371 24055
rect 17313 24015 17371 24021
rect 19794 24012 19800 24064
rect 19852 24052 19858 24064
rect 20162 24052 20168 24064
rect 19852 24024 20168 24052
rect 19852 24012 19858 24024
rect 20162 24012 20168 24024
rect 20220 24012 20226 24064
rect 20254 24012 20260 24064
rect 20312 24052 20318 24064
rect 25869 24055 25927 24061
rect 25869 24052 25881 24055
rect 20312 24024 25881 24052
rect 20312 24012 20318 24024
rect 25869 24021 25881 24024
rect 25915 24052 25927 24055
rect 26050 24052 26056 24064
rect 25915 24024 26056 24052
rect 25915 24021 25927 24024
rect 25869 24015 25927 24021
rect 26050 24012 26056 24024
rect 26108 24012 26114 24064
rect 26694 24052 26700 24064
rect 26655 24024 26700 24052
rect 26694 24012 26700 24024
rect 26752 24012 26758 24064
rect 26804 24052 26832 24092
rect 27614 24080 27620 24132
rect 27672 24120 27678 24132
rect 27908 24120 27936 24228
rect 28353 24191 28411 24197
rect 28353 24157 28365 24191
rect 28399 24157 28411 24191
rect 28534 24188 28540 24200
rect 28495 24160 28540 24188
rect 28353 24151 28411 24157
rect 28368 24120 28396 24151
rect 28534 24148 28540 24160
rect 28592 24148 28598 24200
rect 28644 24197 28672 24228
rect 28736 24197 28764 24364
rect 28994 24352 29000 24404
rect 29052 24392 29058 24404
rect 32490 24392 32496 24404
rect 29052 24364 32496 24392
rect 29052 24352 29058 24364
rect 32490 24352 32496 24364
rect 32548 24352 32554 24404
rect 34514 24392 34520 24404
rect 32876 24364 34520 24392
rect 31202 24324 31208 24336
rect 29012 24296 31208 24324
rect 29012 24265 29040 24296
rect 31202 24284 31208 24296
rect 31260 24284 31266 24336
rect 31754 24284 31760 24336
rect 31812 24324 31818 24336
rect 32876 24324 32904 24364
rect 34514 24352 34520 24364
rect 34572 24352 34578 24404
rect 38102 24392 38108 24404
rect 38063 24364 38108 24392
rect 38102 24352 38108 24364
rect 38160 24352 38166 24404
rect 42058 24352 42064 24404
rect 42116 24392 42122 24404
rect 42705 24395 42763 24401
rect 42705 24392 42717 24395
rect 42116 24364 42717 24392
rect 42116 24352 42122 24364
rect 42705 24361 42717 24364
rect 42751 24361 42763 24395
rect 43530 24392 43536 24404
rect 43491 24364 43536 24392
rect 42705 24355 42763 24361
rect 31812 24296 32904 24324
rect 31812 24284 31818 24296
rect 28997 24259 29055 24265
rect 28997 24225 29009 24259
rect 29043 24225 29055 24259
rect 28997 24219 29055 24225
rect 31110 24216 31116 24268
rect 31168 24256 31174 24268
rect 32861 24259 32919 24265
rect 32861 24256 32873 24259
rect 31168 24228 32873 24256
rect 31168 24216 31174 24228
rect 32861 24225 32873 24228
rect 32907 24225 32919 24259
rect 32861 24219 32919 24225
rect 28629 24191 28687 24197
rect 28629 24157 28641 24191
rect 28675 24157 28687 24191
rect 28629 24151 28687 24157
rect 28721 24191 28779 24197
rect 28721 24157 28733 24191
rect 28767 24157 28779 24191
rect 30929 24191 30987 24197
rect 30929 24188 30941 24191
rect 28721 24151 28779 24157
rect 28828 24160 30941 24188
rect 28442 24120 28448 24132
rect 27672 24092 27936 24120
rect 28355 24092 28448 24120
rect 27672 24080 27678 24092
rect 28442 24080 28448 24092
rect 28500 24120 28506 24132
rect 28828 24120 28856 24160
rect 30929 24157 30941 24160
rect 30975 24188 30987 24191
rect 31478 24188 31484 24200
rect 30975 24160 31484 24188
rect 30975 24157 30987 24160
rect 30929 24151 30987 24157
rect 31478 24148 31484 24160
rect 31536 24148 31542 24200
rect 31573 24191 31631 24197
rect 31573 24157 31585 24191
rect 31619 24157 31631 24191
rect 32876 24188 32904 24219
rect 33962 24216 33968 24268
rect 34020 24256 34026 24268
rect 42720 24256 42748 24355
rect 43530 24352 43536 24364
rect 43588 24352 43594 24404
rect 43162 24256 43168 24268
rect 34020 24228 36216 24256
rect 42720 24228 43168 24256
rect 34020 24216 34026 24228
rect 34238 24188 34244 24200
rect 32876 24160 34244 24188
rect 31573 24151 31631 24157
rect 28500 24092 28856 24120
rect 28500 24080 28506 24092
rect 30466 24080 30472 24132
rect 30524 24120 30530 24132
rect 30745 24123 30803 24129
rect 30745 24120 30757 24123
rect 30524 24092 30757 24120
rect 30524 24080 30530 24092
rect 30745 24089 30757 24092
rect 30791 24089 30803 24123
rect 30745 24083 30803 24089
rect 31113 24123 31171 24129
rect 31113 24089 31125 24123
rect 31159 24120 31171 24123
rect 31588 24120 31616 24151
rect 34238 24148 34244 24160
rect 34296 24188 34302 24200
rect 36081 24191 36139 24197
rect 36081 24188 36093 24191
rect 34296 24160 36093 24188
rect 34296 24148 34302 24160
rect 36081 24157 36093 24160
rect 36127 24157 36139 24191
rect 36188 24188 36216 24228
rect 43162 24216 43168 24228
rect 43220 24216 43226 24268
rect 43990 24256 43996 24268
rect 43951 24228 43996 24256
rect 43990 24216 43996 24228
rect 44048 24216 44054 24268
rect 48130 24256 48136 24268
rect 48091 24228 48136 24256
rect 48130 24216 48136 24228
rect 48188 24216 48194 24268
rect 36188 24160 38884 24188
rect 36081 24151 36139 24157
rect 31846 24120 31852 24132
rect 31159 24092 31616 24120
rect 31807 24092 31852 24120
rect 31159 24089 31171 24092
rect 31113 24083 31171 24089
rect 31846 24080 31852 24092
rect 31904 24080 31910 24132
rect 33134 24129 33140 24132
rect 33128 24083 33140 24129
rect 33192 24120 33198 24132
rect 33192 24092 33228 24120
rect 33704 24092 35020 24120
rect 33134 24080 33140 24083
rect 33192 24080 33198 24092
rect 33704 24052 33732 24092
rect 26804 24024 33732 24052
rect 33778 24012 33784 24064
rect 33836 24052 33842 24064
rect 34241 24055 34299 24061
rect 34241 24052 34253 24055
rect 33836 24024 34253 24052
rect 33836 24012 33842 24024
rect 34241 24021 34253 24024
rect 34287 24052 34299 24055
rect 34882 24052 34888 24064
rect 34287 24024 34888 24052
rect 34287 24021 34299 24024
rect 34241 24015 34299 24021
rect 34882 24012 34888 24024
rect 34940 24012 34946 24064
rect 34992 24052 35020 24092
rect 36170 24080 36176 24132
rect 36228 24120 36234 24132
rect 36326 24123 36384 24129
rect 36326 24120 36338 24123
rect 36228 24092 36338 24120
rect 36228 24080 36234 24092
rect 36326 24089 36338 24092
rect 36372 24089 36384 24123
rect 38856 24120 38884 24160
rect 38930 24148 38936 24200
rect 38988 24188 38994 24200
rect 39485 24191 39543 24197
rect 39485 24188 39497 24191
rect 38988 24160 39497 24188
rect 38988 24148 38994 24160
rect 39485 24157 39497 24160
rect 39531 24188 39543 24191
rect 40862 24188 40868 24200
rect 39531 24160 40868 24188
rect 39531 24157 39543 24160
rect 39485 24151 39543 24157
rect 40862 24148 40868 24160
rect 40920 24188 40926 24200
rect 41325 24191 41383 24197
rect 41325 24188 41337 24191
rect 40920 24160 41337 24188
rect 40920 24148 40926 24160
rect 41325 24157 41337 24160
rect 41371 24188 41383 24191
rect 42702 24188 42708 24200
rect 41371 24160 42708 24188
rect 41371 24157 41383 24160
rect 41325 24151 41383 24157
rect 42702 24148 42708 24160
rect 42760 24148 42766 24200
rect 43346 24188 43352 24200
rect 43259 24160 43352 24188
rect 43346 24148 43352 24160
rect 43404 24148 43410 24200
rect 44174 24188 44180 24200
rect 44135 24160 44180 24188
rect 44174 24148 44180 24160
rect 44232 24148 44238 24200
rect 46474 24188 46480 24200
rect 46435 24160 46480 24188
rect 46474 24148 46480 24160
rect 46532 24148 46538 24200
rect 39114 24120 39120 24132
rect 36326 24083 36384 24089
rect 36556 24092 38240 24120
rect 38856 24092 39120 24120
rect 36556 24052 36584 24092
rect 34992 24024 36584 24052
rect 36722 24012 36728 24064
rect 36780 24052 36786 24064
rect 37461 24055 37519 24061
rect 37461 24052 37473 24055
rect 36780 24024 37473 24052
rect 36780 24012 36786 24024
rect 37461 24021 37473 24024
rect 37507 24021 37519 24055
rect 38212 24052 38240 24092
rect 39114 24080 39120 24092
rect 39172 24080 39178 24132
rect 39206 24080 39212 24132
rect 39264 24129 39270 24132
rect 41598 24129 41604 24132
rect 39264 24120 39276 24129
rect 41592 24120 41604 24129
rect 39264 24092 39309 24120
rect 41559 24092 41604 24120
rect 39264 24083 39276 24092
rect 41592 24083 41604 24092
rect 39264 24080 39270 24083
rect 41598 24080 41604 24083
rect 41656 24080 41662 24132
rect 42334 24080 42340 24132
rect 42392 24120 42398 24132
rect 43364 24120 43392 24148
rect 42392 24092 43392 24120
rect 46661 24123 46719 24129
rect 42392 24080 42398 24092
rect 46661 24089 46673 24123
rect 46707 24120 46719 24123
rect 47854 24120 47860 24132
rect 46707 24092 47860 24120
rect 46707 24089 46719 24092
rect 46661 24083 46719 24089
rect 47854 24080 47860 24092
rect 47912 24080 47918 24132
rect 42794 24052 42800 24064
rect 38212 24024 42800 24052
rect 37461 24015 37519 24021
rect 42794 24012 42800 24024
rect 42852 24012 42858 24064
rect 44266 24012 44272 24064
rect 44324 24052 44330 24064
rect 44361 24055 44419 24061
rect 44361 24052 44373 24055
rect 44324 24024 44373 24052
rect 44324 24012 44330 24024
rect 44361 24021 44373 24024
rect 44407 24021 44419 24055
rect 44361 24015 44419 24021
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 6638 23848 6644 23860
rect 6599 23820 6644 23848
rect 6638 23808 6644 23820
rect 6696 23808 6702 23860
rect 8846 23848 8852 23860
rect 8807 23820 8852 23848
rect 8846 23808 8852 23820
rect 8904 23808 8910 23860
rect 9677 23851 9735 23857
rect 9677 23817 9689 23851
rect 9723 23817 9735 23851
rect 10134 23848 10140 23860
rect 10095 23820 10140 23848
rect 9677 23811 9735 23817
rect 6546 23712 6552 23724
rect 6507 23684 6552 23712
rect 6546 23672 6552 23684
rect 6604 23672 6610 23724
rect 9033 23715 9091 23721
rect 9033 23681 9045 23715
rect 9079 23712 9091 23715
rect 9692 23712 9720 23811
rect 10134 23808 10140 23820
rect 10192 23808 10198 23860
rect 15378 23848 15384 23860
rect 15339 23820 15384 23848
rect 15378 23808 15384 23820
rect 15436 23808 15442 23860
rect 17126 23808 17132 23860
rect 17184 23848 17190 23860
rect 20254 23848 20260 23860
rect 17184 23820 20260 23848
rect 17184 23808 17190 23820
rect 20254 23808 20260 23820
rect 20312 23808 20318 23860
rect 20622 23848 20628 23860
rect 20583 23820 20628 23848
rect 20622 23808 20628 23820
rect 20680 23808 20686 23860
rect 22741 23851 22799 23857
rect 22741 23817 22753 23851
rect 22787 23848 22799 23851
rect 23106 23848 23112 23860
rect 22787 23820 23112 23848
rect 22787 23817 22799 23820
rect 22741 23811 22799 23817
rect 23106 23808 23112 23820
rect 23164 23808 23170 23860
rect 23566 23848 23572 23860
rect 23527 23820 23572 23848
rect 23566 23808 23572 23820
rect 23624 23808 23630 23860
rect 23658 23808 23664 23860
rect 23716 23848 23722 23860
rect 24029 23851 24087 23857
rect 24029 23848 24041 23851
rect 23716 23820 24041 23848
rect 23716 23808 23722 23820
rect 24029 23817 24041 23820
rect 24075 23817 24087 23851
rect 24029 23811 24087 23817
rect 26326 23808 26332 23860
rect 26384 23848 26390 23860
rect 26421 23851 26479 23857
rect 26421 23848 26433 23851
rect 26384 23820 26433 23848
rect 26384 23808 26390 23820
rect 26421 23817 26433 23820
rect 26467 23817 26479 23851
rect 27157 23851 27215 23857
rect 27157 23848 27169 23851
rect 26421 23811 26479 23817
rect 26528 23820 27169 23848
rect 20346 23780 20352 23792
rect 19260 23752 20352 23780
rect 9079 23684 9720 23712
rect 10045 23715 10103 23721
rect 9079 23681 9091 23684
rect 9033 23675 9091 23681
rect 10045 23681 10057 23715
rect 10091 23712 10103 23715
rect 11698 23712 11704 23724
rect 10091 23684 11704 23712
rect 10091 23681 10103 23684
rect 10045 23675 10103 23681
rect 11698 23672 11704 23684
rect 11756 23672 11762 23724
rect 14274 23721 14280 23724
rect 14268 23675 14280 23721
rect 14332 23712 14338 23724
rect 19260 23721 19288 23752
rect 20346 23740 20352 23752
rect 20404 23740 20410 23792
rect 23124 23780 23152 23808
rect 23584 23780 23612 23808
rect 22572 23752 22876 23780
rect 23124 23752 23520 23780
rect 23584 23752 24256 23780
rect 19245 23715 19303 23721
rect 14332 23684 14368 23712
rect 14274 23672 14280 23675
rect 14332 23672 14338 23684
rect 19245 23681 19257 23715
rect 19291 23681 19303 23715
rect 19245 23675 19303 23681
rect 19334 23672 19340 23724
rect 19392 23712 19398 23724
rect 22572 23721 22600 23752
rect 19501 23715 19559 23721
rect 19501 23712 19513 23715
rect 19392 23684 19513 23712
rect 19392 23672 19398 23684
rect 19501 23681 19513 23684
rect 19547 23681 19559 23715
rect 19501 23675 19559 23681
rect 22557 23715 22615 23721
rect 22557 23681 22569 23715
rect 22603 23681 22615 23715
rect 22557 23675 22615 23681
rect 22741 23715 22799 23721
rect 22741 23681 22753 23715
rect 22787 23681 22799 23715
rect 22848 23712 22876 23752
rect 23198 23712 23204 23724
rect 22848 23684 23204 23712
rect 22741 23675 22799 23681
rect 9306 23604 9312 23656
rect 9364 23644 9370 23656
rect 10229 23647 10287 23653
rect 10229 23644 10241 23647
rect 9364 23616 10241 23644
rect 9364 23604 9370 23616
rect 10229 23613 10241 23616
rect 10275 23613 10287 23647
rect 10229 23607 10287 23613
rect 13078 23604 13084 23656
rect 13136 23644 13142 23656
rect 13630 23644 13636 23656
rect 13136 23616 13636 23644
rect 13136 23604 13142 23616
rect 13630 23604 13636 23616
rect 13688 23644 13694 23656
rect 14001 23647 14059 23653
rect 14001 23644 14013 23647
rect 13688 23616 14013 23644
rect 13688 23604 13694 23616
rect 14001 23613 14013 23616
rect 14047 23613 14059 23647
rect 14001 23607 14059 23613
rect 22756 23576 22784 23675
rect 23198 23672 23204 23684
rect 23256 23672 23262 23724
rect 23385 23715 23443 23721
rect 23385 23681 23397 23715
rect 23431 23681 23443 23715
rect 23492 23712 23520 23752
rect 24228 23721 24256 23752
rect 24029 23715 24087 23721
rect 24029 23712 24041 23715
rect 23492 23684 24041 23712
rect 23385 23675 23443 23681
rect 24029 23681 24041 23684
rect 24075 23681 24087 23715
rect 24029 23675 24087 23681
rect 24213 23715 24271 23721
rect 24213 23681 24225 23715
rect 24259 23681 24271 23715
rect 24213 23675 24271 23681
rect 23400 23644 23428 23675
rect 25498 23644 25504 23656
rect 23400 23616 25504 23644
rect 23400 23576 23428 23616
rect 25498 23604 25504 23616
rect 25556 23604 25562 23656
rect 26436 23644 26464 23811
rect 26528 23789 26556 23820
rect 27157 23817 27169 23820
rect 27203 23817 27215 23851
rect 27157 23811 27215 23817
rect 28442 23808 28448 23860
rect 28500 23848 28506 23860
rect 28537 23851 28595 23857
rect 28537 23848 28549 23851
rect 28500 23820 28549 23848
rect 28500 23808 28506 23820
rect 28537 23817 28549 23820
rect 28583 23817 28595 23851
rect 28537 23811 28595 23817
rect 28644 23820 31754 23848
rect 26513 23783 26571 23789
rect 26513 23749 26525 23783
rect 26559 23749 26571 23783
rect 26513 23743 26571 23749
rect 27706 23712 27712 23724
rect 27667 23684 27712 23712
rect 27706 23672 27712 23684
rect 27764 23672 27770 23724
rect 27154 23644 27160 23656
rect 26436 23616 27160 23644
rect 27154 23604 27160 23616
rect 27212 23604 27218 23656
rect 27433 23647 27491 23653
rect 27433 23613 27445 23647
rect 27479 23644 27491 23647
rect 27614 23644 27620 23656
rect 27479 23616 27620 23644
rect 27479 23613 27491 23616
rect 27433 23607 27491 23613
rect 27614 23604 27620 23616
rect 27672 23604 27678 23656
rect 22756 23548 23428 23576
rect 23474 23536 23480 23588
rect 23532 23576 23538 23588
rect 28644 23576 28672 23820
rect 29672 23783 29730 23789
rect 29672 23749 29684 23783
rect 29718 23780 29730 23783
rect 30742 23780 30748 23792
rect 29718 23752 30748 23780
rect 29718 23749 29730 23752
rect 29672 23743 29730 23749
rect 30742 23740 30748 23752
rect 30800 23740 30806 23792
rect 31726 23780 31754 23820
rect 32490 23808 32496 23860
rect 32548 23848 32554 23860
rect 33042 23848 33048 23860
rect 32548 23820 33048 23848
rect 32548 23808 32554 23820
rect 33042 23808 33048 23820
rect 33100 23808 33106 23860
rect 36081 23851 36139 23857
rect 36081 23817 36093 23851
rect 36127 23848 36139 23851
rect 36170 23848 36176 23860
rect 36127 23820 36176 23848
rect 36127 23817 36139 23820
rect 36081 23811 36139 23817
rect 36170 23808 36176 23820
rect 36228 23808 36234 23860
rect 38838 23848 38844 23860
rect 38799 23820 38844 23848
rect 38838 23808 38844 23820
rect 38896 23808 38902 23860
rect 39022 23808 39028 23860
rect 39080 23848 39086 23860
rect 43622 23848 43628 23860
rect 39080 23820 43628 23848
rect 39080 23808 39086 23820
rect 43622 23808 43628 23820
rect 43680 23808 43686 23860
rect 44453 23851 44511 23857
rect 44453 23817 44465 23851
rect 44499 23848 44511 23851
rect 44542 23848 44548 23860
rect 44499 23820 44548 23848
rect 44499 23817 44511 23820
rect 44453 23811 44511 23817
rect 44542 23808 44548 23820
rect 44600 23808 44606 23860
rect 47854 23848 47860 23860
rect 47815 23820 47860 23848
rect 47854 23808 47860 23820
rect 47912 23808 47918 23860
rect 47118 23780 47124 23792
rect 31726 23752 47124 23780
rect 47118 23740 47124 23752
rect 47176 23780 47182 23792
rect 47176 23752 47808 23780
rect 47176 23740 47182 23752
rect 30374 23712 30380 23724
rect 30335 23684 30380 23712
rect 30374 23672 30380 23684
rect 30432 23672 30438 23724
rect 30466 23672 30472 23724
rect 30524 23712 30530 23724
rect 31481 23715 31539 23721
rect 31481 23712 31493 23715
rect 30524 23684 31493 23712
rect 30524 23672 30530 23684
rect 31481 23681 31493 23684
rect 31527 23681 31539 23715
rect 31481 23675 31539 23681
rect 33321 23715 33379 23721
rect 33321 23681 33333 23715
rect 33367 23681 33379 23715
rect 33321 23675 33379 23681
rect 29917 23647 29975 23653
rect 29917 23613 29929 23647
rect 29963 23644 29975 23647
rect 31110 23644 31116 23656
rect 29963 23616 31116 23644
rect 29963 23613 29975 23616
rect 29917 23607 29975 23613
rect 31110 23604 31116 23616
rect 31168 23604 31174 23656
rect 33336 23644 33364 23675
rect 33502 23672 33508 23724
rect 33560 23712 33566 23724
rect 33597 23715 33655 23721
rect 33597 23712 33609 23715
rect 33560 23684 33609 23712
rect 33560 23672 33566 23684
rect 33597 23681 33609 23684
rect 33643 23681 33655 23715
rect 33778 23712 33784 23724
rect 33739 23684 33784 23712
rect 33597 23675 33655 23681
rect 33778 23672 33784 23684
rect 33836 23672 33842 23724
rect 34238 23712 34244 23724
rect 34199 23684 34244 23712
rect 34238 23672 34244 23684
rect 34296 23672 34302 23724
rect 34508 23715 34566 23721
rect 34508 23681 34520 23715
rect 34554 23712 34566 23715
rect 34790 23712 34796 23724
rect 34554 23684 34796 23712
rect 34554 23681 34566 23684
rect 34508 23675 34566 23681
rect 34790 23672 34796 23684
rect 34848 23672 34854 23724
rect 34882 23672 34888 23724
rect 34940 23712 34946 23724
rect 36265 23715 36323 23721
rect 36265 23712 36277 23715
rect 34940 23684 36277 23712
rect 34940 23672 34946 23684
rect 36265 23681 36277 23684
rect 36311 23681 36323 23715
rect 36630 23712 36636 23724
rect 36591 23684 36636 23712
rect 36265 23675 36323 23681
rect 36630 23672 36636 23684
rect 36688 23672 36694 23724
rect 36817 23715 36875 23721
rect 36817 23681 36829 23715
rect 36863 23712 36875 23715
rect 37642 23712 37648 23724
rect 36863 23684 37648 23712
rect 36863 23681 36875 23684
rect 36817 23675 36875 23681
rect 37642 23672 37648 23684
rect 37700 23672 37706 23724
rect 37734 23672 37740 23724
rect 37792 23712 37798 23724
rect 39025 23715 39083 23721
rect 39025 23712 39037 23715
rect 37792 23684 39037 23712
rect 37792 23672 37798 23684
rect 39025 23681 39037 23684
rect 39071 23681 39083 23715
rect 39025 23675 39083 23681
rect 39114 23672 39120 23724
rect 39172 23712 39178 23724
rect 39301 23715 39359 23721
rect 39301 23712 39313 23715
rect 39172 23684 39313 23712
rect 39172 23672 39178 23684
rect 39301 23681 39313 23684
rect 39347 23681 39359 23715
rect 39482 23712 39488 23724
rect 39443 23684 39488 23712
rect 39301 23675 39359 23681
rect 33686 23644 33692 23656
rect 33336 23616 33692 23644
rect 33686 23604 33692 23616
rect 33744 23604 33750 23656
rect 36446 23644 36452 23656
rect 36407 23616 36452 23644
rect 36446 23604 36452 23616
rect 36504 23604 36510 23656
rect 36541 23647 36599 23653
rect 36541 23613 36553 23647
rect 36587 23644 36599 23647
rect 36722 23644 36728 23656
rect 36587 23616 36728 23644
rect 36587 23613 36599 23616
rect 36541 23607 36599 23613
rect 36722 23604 36728 23616
rect 36780 23604 36786 23656
rect 39316 23644 39344 23675
rect 39482 23672 39488 23684
rect 39540 23672 39546 23724
rect 40681 23715 40739 23721
rect 40681 23681 40693 23715
rect 40727 23712 40739 23715
rect 43254 23712 43260 23724
rect 40727 23684 43260 23712
rect 40727 23681 40739 23684
rect 40681 23675 40739 23681
rect 43254 23672 43260 23684
rect 43312 23672 43318 23724
rect 44266 23712 44272 23724
rect 44227 23684 44272 23712
rect 44266 23672 44272 23684
rect 44324 23672 44330 23724
rect 46474 23672 46480 23724
rect 46532 23712 46538 23724
rect 47780 23721 47808 23752
rect 47029 23715 47087 23721
rect 47029 23712 47041 23715
rect 46532 23684 47041 23712
rect 46532 23672 46538 23684
rect 47029 23681 47041 23684
rect 47075 23681 47087 23715
rect 47029 23675 47087 23681
rect 47765 23715 47823 23721
rect 47765 23681 47777 23715
rect 47811 23681 47823 23715
rect 47765 23675 47823 23681
rect 39390 23644 39396 23656
rect 39316 23616 39396 23644
rect 39390 23604 39396 23616
rect 39448 23604 39454 23656
rect 23532 23548 28672 23576
rect 23532 23536 23538 23548
rect 30282 23536 30288 23588
rect 30340 23576 30346 23588
rect 30561 23579 30619 23585
rect 30561 23576 30573 23579
rect 30340 23548 30573 23576
rect 30340 23536 30346 23548
rect 30561 23545 30573 23548
rect 30607 23545 30619 23579
rect 39022 23576 39028 23588
rect 30561 23539 30619 23545
rect 30668 23548 34284 23576
rect 20530 23468 20536 23520
rect 20588 23508 20594 23520
rect 26602 23508 26608 23520
rect 20588 23480 26608 23508
rect 20588 23468 20594 23480
rect 26602 23468 26608 23480
rect 26660 23508 26666 23520
rect 27341 23511 27399 23517
rect 27341 23508 27353 23511
rect 26660 23480 27353 23508
rect 26660 23468 26666 23480
rect 27341 23477 27353 23480
rect 27387 23508 27399 23511
rect 27798 23508 27804 23520
rect 27387 23480 27804 23508
rect 27387 23477 27399 23480
rect 27341 23471 27399 23477
rect 27798 23468 27804 23480
rect 27856 23468 27862 23520
rect 29270 23468 29276 23520
rect 29328 23508 29334 23520
rect 30668 23508 30696 23548
rect 31662 23508 31668 23520
rect 29328 23480 30696 23508
rect 31623 23480 31668 23508
rect 29328 23468 29334 23480
rect 31662 23468 31668 23480
rect 31720 23468 31726 23520
rect 33137 23511 33195 23517
rect 33137 23477 33149 23511
rect 33183 23508 33195 23511
rect 33226 23508 33232 23520
rect 33183 23480 33232 23508
rect 33183 23477 33195 23480
rect 33137 23471 33195 23477
rect 33226 23468 33232 23480
rect 33284 23468 33290 23520
rect 34256 23508 34284 23548
rect 35176 23548 39028 23576
rect 35176 23508 35204 23548
rect 39022 23536 39028 23548
rect 39080 23536 39086 23588
rect 35618 23508 35624 23520
rect 34256 23480 35204 23508
rect 35579 23480 35624 23508
rect 35618 23468 35624 23480
rect 35676 23468 35682 23520
rect 36078 23468 36084 23520
rect 36136 23508 36142 23520
rect 36630 23508 36636 23520
rect 36136 23480 36636 23508
rect 36136 23468 36142 23480
rect 36630 23468 36636 23480
rect 36688 23468 36694 23520
rect 40402 23508 40408 23520
rect 40363 23480 40408 23508
rect 40402 23468 40408 23480
rect 40460 23508 40466 23520
rect 42794 23508 42800 23520
rect 40460 23480 42800 23508
rect 40460 23468 40466 23480
rect 42794 23468 42800 23480
rect 42852 23508 42858 23520
rect 42978 23508 42984 23520
rect 42852 23480 42984 23508
rect 42852 23468 42858 23480
rect 42978 23468 42984 23480
rect 43036 23468 43042 23520
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 14274 23304 14280 23316
rect 14235 23276 14280 23304
rect 14274 23264 14280 23276
rect 14332 23264 14338 23316
rect 21266 23264 21272 23316
rect 21324 23304 21330 23316
rect 26329 23307 26387 23313
rect 21324 23276 22094 23304
rect 21324 23264 21330 23276
rect 14642 23196 14648 23248
rect 14700 23196 14706 23248
rect 22066 23236 22094 23276
rect 26329 23273 26341 23307
rect 26375 23304 26387 23307
rect 26694 23304 26700 23316
rect 26375 23276 26700 23304
rect 26375 23273 26387 23276
rect 26329 23267 26387 23273
rect 26694 23264 26700 23276
rect 26752 23304 26758 23316
rect 31757 23307 31815 23313
rect 26752 23276 27752 23304
rect 26752 23264 26758 23276
rect 27724 23248 27752 23276
rect 31757 23273 31769 23307
rect 31803 23304 31815 23307
rect 32582 23304 32588 23316
rect 31803 23276 32588 23304
rect 31803 23273 31815 23276
rect 31757 23267 31815 23273
rect 32582 23264 32588 23276
rect 32640 23264 32646 23316
rect 33045 23307 33103 23313
rect 33045 23273 33057 23307
rect 33091 23304 33103 23307
rect 33134 23304 33140 23316
rect 33091 23276 33140 23304
rect 33091 23273 33103 23276
rect 33045 23267 33103 23273
rect 33134 23264 33140 23276
rect 33192 23264 33198 23316
rect 34790 23264 34796 23316
rect 34848 23304 34854 23316
rect 34885 23307 34943 23313
rect 34885 23304 34897 23307
rect 34848 23276 34897 23304
rect 34848 23264 34854 23276
rect 34885 23273 34897 23276
rect 34931 23273 34943 23307
rect 37642 23304 37648 23316
rect 37603 23276 37648 23304
rect 34885 23267 34943 23273
rect 37642 23264 37648 23276
rect 37700 23264 37706 23316
rect 42334 23304 42340 23316
rect 42295 23276 42340 23304
rect 42334 23264 42340 23276
rect 42392 23264 42398 23316
rect 48038 23304 48044 23316
rect 42536 23276 48044 23304
rect 27706 23236 27712 23248
rect 22066 23208 27476 23236
rect 27619 23208 27712 23236
rect 12345 23171 12403 23177
rect 12345 23137 12357 23171
rect 12391 23168 12403 23171
rect 12434 23168 12440 23180
rect 12391 23140 12440 23168
rect 12391 23137 12403 23140
rect 12345 23131 12403 23137
rect 11698 23060 11704 23112
rect 11756 23100 11762 23112
rect 12069 23103 12127 23109
rect 12069 23100 12081 23103
rect 11756 23072 12081 23100
rect 11756 23060 11762 23072
rect 12069 23069 12081 23072
rect 12115 23069 12127 23103
rect 12069 23063 12127 23069
rect 12360 23032 12388 23131
rect 12434 23128 12440 23140
rect 12492 23128 12498 23180
rect 14660 23168 14688 23196
rect 14737 23171 14795 23177
rect 14737 23168 14749 23171
rect 14660 23140 14749 23168
rect 14737 23137 14749 23140
rect 14783 23168 14795 23171
rect 19978 23168 19984 23180
rect 14783 23140 19984 23168
rect 14783 23137 14795 23140
rect 14737 23131 14795 23137
rect 19978 23128 19984 23140
rect 20036 23128 20042 23180
rect 22370 23168 22376 23180
rect 22331 23140 22376 23168
rect 22370 23128 22376 23140
rect 22428 23128 22434 23180
rect 22465 23171 22523 23177
rect 22465 23137 22477 23171
rect 22511 23168 22523 23171
rect 23198 23168 23204 23180
rect 22511 23140 23204 23168
rect 22511 23137 22523 23140
rect 22465 23131 22523 23137
rect 23198 23128 23204 23140
rect 23256 23128 23262 23180
rect 24949 23171 25007 23177
rect 24949 23137 24961 23171
rect 24995 23168 25007 23171
rect 26970 23168 26976 23180
rect 24995 23140 26976 23168
rect 24995 23137 25007 23140
rect 24949 23131 25007 23137
rect 26970 23128 26976 23140
rect 27028 23128 27034 23180
rect 14458 23100 14464 23112
rect 14419 23072 14464 23100
rect 14458 23060 14464 23072
rect 14516 23060 14522 23112
rect 14642 23060 14648 23112
rect 14700 23100 14706 23112
rect 15010 23100 15016 23112
rect 14700 23072 15016 23100
rect 14700 23060 14706 23072
rect 15010 23060 15016 23072
rect 15068 23060 15074 23112
rect 19889 23103 19947 23109
rect 19889 23069 19901 23103
rect 19935 23069 19947 23103
rect 24762 23100 24768 23112
rect 24723 23072 24768 23100
rect 19889 23063 19947 23069
rect 19613 23035 19671 23041
rect 19613 23032 19625 23035
rect 12360 23004 19625 23032
rect 19613 23001 19625 23004
rect 19659 23001 19671 23035
rect 19904 23032 19932 23063
rect 24762 23060 24768 23072
rect 24820 23060 24826 23112
rect 25038 23060 25044 23112
rect 25096 23100 25102 23112
rect 27338 23100 27344 23112
rect 25096 23072 25141 23100
rect 26436 23072 27344 23100
rect 25096 23060 25102 23072
rect 26313 23035 26371 23041
rect 19904 23004 26188 23032
rect 19613 22995 19671 23001
rect 11606 22924 11612 22976
rect 11664 22964 11670 22976
rect 11701 22967 11759 22973
rect 11701 22964 11713 22967
rect 11664 22936 11713 22964
rect 11664 22924 11670 22936
rect 11701 22933 11713 22936
rect 11747 22933 11759 22967
rect 11701 22927 11759 22933
rect 12161 22967 12219 22973
rect 12161 22933 12173 22967
rect 12207 22964 12219 22967
rect 12802 22964 12808 22976
rect 12207 22936 12808 22964
rect 12207 22933 12219 22936
rect 12161 22927 12219 22933
rect 12802 22924 12808 22936
rect 12860 22924 12866 22976
rect 16206 22924 16212 22976
rect 16264 22964 16270 22976
rect 17586 22964 17592 22976
rect 16264 22936 17592 22964
rect 16264 22924 16270 22936
rect 17586 22924 17592 22936
rect 17644 22924 17650 22976
rect 22557 22967 22615 22973
rect 22557 22933 22569 22967
rect 22603 22964 22615 22967
rect 22646 22964 22652 22976
rect 22603 22936 22652 22964
rect 22603 22933 22615 22936
rect 22557 22927 22615 22933
rect 22646 22924 22652 22936
rect 22704 22924 22710 22976
rect 22738 22924 22744 22976
rect 22796 22964 22802 22976
rect 22925 22967 22983 22973
rect 22925 22964 22937 22967
rect 22796 22936 22937 22964
rect 22796 22924 22802 22936
rect 22925 22933 22937 22936
rect 22971 22933 22983 22967
rect 24578 22964 24584 22976
rect 24539 22936 24584 22964
rect 22925 22927 22983 22933
rect 24578 22924 24584 22936
rect 24636 22924 24642 22976
rect 26160 22973 26188 23004
rect 26313 23001 26325 23035
rect 26359 23032 26371 23035
rect 26436 23032 26464 23072
rect 27338 23060 27344 23072
rect 27396 23060 27402 23112
rect 26359 23004 26464 23032
rect 26513 23035 26571 23041
rect 26359 23001 26371 23004
rect 26313 22995 26371 23001
rect 26513 23001 26525 23035
rect 26559 23032 26571 23035
rect 26602 23032 26608 23044
rect 26559 23004 26608 23032
rect 26559 23001 26571 23004
rect 26513 22995 26571 23001
rect 26602 22992 26608 23004
rect 26660 22992 26666 23044
rect 27448 23032 27476 23208
rect 27706 23196 27712 23208
rect 27764 23236 27770 23248
rect 29270 23236 29276 23248
rect 27764 23208 29276 23236
rect 27764 23196 27770 23208
rect 29270 23196 29276 23208
rect 29328 23196 29334 23248
rect 32214 23196 32220 23248
rect 32272 23236 32278 23248
rect 42536 23236 42564 23276
rect 48038 23264 48044 23276
rect 48096 23264 48102 23316
rect 32272 23208 42564 23236
rect 42613 23239 42671 23245
rect 32272 23196 32278 23208
rect 42613 23205 42625 23239
rect 42659 23236 42671 23239
rect 43254 23236 43260 23248
rect 42659 23208 43260 23236
rect 42659 23205 42671 23208
rect 42613 23199 42671 23205
rect 43254 23196 43260 23208
rect 43312 23196 43318 23248
rect 27724 23168 27752 23196
rect 27632 23140 27752 23168
rect 27985 23171 28043 23177
rect 27632 23112 27660 23140
rect 27985 23137 27997 23171
rect 28031 23168 28043 23171
rect 28031 23140 28580 23168
rect 28031 23137 28043 23140
rect 27985 23131 28043 23137
rect 28552 23112 28580 23140
rect 30098 23128 30104 23180
rect 30156 23168 30162 23180
rect 31570 23168 31576 23180
rect 30156 23140 31576 23168
rect 30156 23128 30162 23140
rect 31570 23128 31576 23140
rect 31628 23168 31634 23180
rect 33413 23171 33471 23177
rect 33413 23168 33425 23171
rect 31628 23140 33425 23168
rect 31628 23128 31634 23140
rect 33413 23137 33425 23140
rect 33459 23137 33471 23171
rect 33413 23131 33471 23137
rect 33505 23171 33563 23177
rect 33505 23137 33517 23171
rect 33551 23168 33563 23171
rect 33594 23168 33600 23180
rect 33551 23140 33600 23168
rect 33551 23137 33563 23140
rect 33505 23131 33563 23137
rect 33594 23128 33600 23140
rect 33652 23128 33658 23180
rect 35345 23171 35403 23177
rect 35345 23137 35357 23171
rect 35391 23168 35403 23171
rect 35618 23168 35624 23180
rect 35391 23140 35624 23168
rect 35391 23137 35403 23140
rect 35345 23131 35403 23137
rect 35618 23128 35624 23140
rect 35676 23168 35682 23180
rect 39850 23168 39856 23180
rect 35676 23140 36584 23168
rect 35676 23128 35682 23140
rect 27614 23100 27620 23112
rect 27527 23072 27620 23100
rect 27614 23060 27620 23072
rect 27672 23060 27678 23112
rect 28442 23100 28448 23112
rect 27724 23072 28304 23100
rect 28403 23072 28448 23100
rect 27724 23032 27752 23072
rect 27448 23004 27752 23032
rect 27798 22992 27804 23044
rect 27856 23032 27862 23044
rect 27856 23004 27901 23032
rect 27856 22992 27862 23004
rect 26145 22967 26203 22973
rect 26145 22933 26157 22967
rect 26191 22933 26203 22967
rect 28276 22964 28304 23072
rect 28442 23060 28448 23072
rect 28500 23060 28506 23112
rect 28534 23060 28540 23112
rect 28592 23100 28598 23112
rect 28629 23103 28687 23109
rect 28629 23100 28641 23103
rect 28592 23072 28641 23100
rect 28592 23060 28598 23072
rect 28629 23069 28641 23072
rect 28675 23069 28687 23103
rect 30282 23100 30288 23112
rect 30243 23072 30288 23100
rect 28629 23063 28687 23069
rect 30282 23060 30288 23072
rect 30340 23060 30346 23112
rect 30466 23100 30472 23112
rect 30427 23072 30472 23100
rect 30466 23060 30472 23072
rect 30524 23060 30530 23112
rect 30745 23103 30803 23109
rect 30745 23069 30757 23103
rect 30791 23100 30803 23103
rect 31662 23100 31668 23112
rect 30791 23072 31668 23100
rect 30791 23069 30803 23072
rect 30745 23063 30803 23069
rect 31662 23060 31668 23072
rect 31720 23060 31726 23112
rect 33226 23100 33232 23112
rect 33187 23072 33232 23100
rect 33226 23060 33232 23072
rect 33284 23060 33290 23112
rect 34698 23060 34704 23112
rect 34756 23100 34762 23112
rect 36556 23109 36584 23140
rect 37568 23140 39856 23168
rect 35069 23103 35127 23109
rect 35069 23100 35081 23103
rect 34756 23072 35081 23100
rect 34756 23060 34762 23072
rect 35069 23069 35081 23072
rect 35115 23069 35127 23103
rect 35069 23063 35127 23069
rect 35253 23103 35311 23109
rect 35253 23069 35265 23103
rect 35299 23069 35311 23103
rect 35253 23063 35311 23069
rect 36541 23103 36599 23109
rect 36541 23069 36553 23103
rect 36587 23069 36599 23103
rect 36722 23100 36728 23112
rect 36683 23072 36728 23100
rect 36541 23063 36599 23069
rect 28813 23035 28871 23041
rect 28813 23001 28825 23035
rect 28859 23032 28871 23035
rect 30374 23032 30380 23044
rect 28859 23004 30380 23032
rect 28859 23001 28871 23004
rect 28813 22995 28871 23001
rect 30374 22992 30380 23004
rect 30432 22992 30438 23044
rect 30484 23032 30512 23060
rect 31481 23035 31539 23041
rect 31481 23032 31493 23035
rect 30484 23004 31493 23032
rect 31481 23001 31493 23004
rect 31527 23001 31539 23035
rect 31481 22995 31539 23001
rect 32950 22992 32956 23044
rect 33008 23032 33014 23044
rect 35268 23032 35296 23063
rect 36722 23060 36728 23072
rect 36780 23060 36786 23112
rect 37568 23109 37596 23140
rect 39850 23128 39856 23140
rect 39908 23168 39914 23180
rect 40402 23168 40408 23180
rect 39908 23140 40408 23168
rect 39908 23128 39914 23140
rect 40402 23128 40408 23140
rect 40460 23128 40466 23180
rect 42705 23171 42763 23177
rect 42705 23137 42717 23171
rect 42751 23168 42763 23171
rect 43162 23168 43168 23180
rect 42751 23140 43168 23168
rect 42751 23137 42763 23140
rect 42705 23131 42763 23137
rect 43162 23128 43168 23140
rect 43220 23128 43226 23180
rect 37553 23103 37611 23109
rect 37553 23069 37565 23103
rect 37599 23069 37611 23103
rect 37734 23100 37740 23112
rect 37695 23072 37740 23100
rect 37553 23063 37611 23069
rect 37734 23060 37740 23072
rect 37792 23060 37798 23112
rect 42521 23103 42579 23109
rect 42521 23069 42533 23103
rect 42567 23069 42579 23103
rect 42521 23063 42579 23069
rect 42797 23103 42855 23109
rect 42797 23069 42809 23103
rect 42843 23100 42855 23103
rect 43438 23100 43444 23112
rect 42843 23072 43444 23100
rect 42843 23069 42855 23072
rect 42797 23063 42855 23069
rect 38654 23032 38660 23044
rect 33008 23004 38660 23032
rect 33008 22992 33014 23004
rect 38654 22992 38660 23004
rect 38712 22992 38718 23044
rect 42536 23032 42564 23063
rect 43438 23060 43444 23072
rect 43496 23060 43502 23112
rect 43070 23032 43076 23044
rect 42536 23004 43076 23032
rect 43070 22992 43076 23004
rect 43128 22992 43134 23044
rect 30558 22964 30564 22976
rect 28276 22936 30564 22964
rect 26145 22927 26203 22933
rect 30558 22924 30564 22936
rect 30616 22924 30622 22976
rect 30929 22967 30987 22973
rect 30929 22933 30941 22967
rect 30975 22964 30987 22967
rect 31294 22964 31300 22976
rect 30975 22936 31300 22964
rect 30975 22933 30987 22936
rect 30929 22927 30987 22933
rect 31294 22924 31300 22936
rect 31352 22924 31358 22976
rect 36354 22964 36360 22976
rect 36315 22936 36360 22964
rect 36354 22924 36360 22936
rect 36412 22924 36418 22976
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 11149 22763 11207 22769
rect 11149 22729 11161 22763
rect 11195 22729 11207 22763
rect 11698 22760 11704 22772
rect 11659 22732 11704 22760
rect 11149 22723 11207 22729
rect 11164 22692 11192 22723
rect 11698 22720 11704 22732
rect 11756 22720 11762 22772
rect 23198 22720 23204 22772
rect 23256 22760 23262 22772
rect 23385 22763 23443 22769
rect 23385 22760 23397 22763
rect 23256 22732 23397 22760
rect 23256 22720 23262 22732
rect 23385 22729 23397 22732
rect 23431 22729 23443 22763
rect 23385 22723 23443 22729
rect 27433 22763 27491 22769
rect 27433 22729 27445 22763
rect 27479 22760 27491 22763
rect 27522 22760 27528 22772
rect 27479 22732 27528 22760
rect 27479 22729 27491 22732
rect 27433 22723 27491 22729
rect 27522 22720 27528 22732
rect 27580 22760 27586 22772
rect 27706 22760 27712 22772
rect 27580 22732 27712 22760
rect 27580 22720 27586 22732
rect 27706 22720 27712 22732
rect 27764 22720 27770 22772
rect 42794 22720 42800 22772
rect 42852 22720 42858 22772
rect 42886 22720 42892 22772
rect 42944 22760 42950 22772
rect 42944 22732 43116 22760
rect 42944 22720 42950 22732
rect 12814 22695 12872 22701
rect 12814 22692 12826 22695
rect 11164 22664 12826 22692
rect 12814 22661 12826 22664
rect 12860 22661 12872 22695
rect 12814 22655 12872 22661
rect 20104 22695 20162 22701
rect 20104 22661 20116 22695
rect 20150 22692 20162 22695
rect 20809 22695 20867 22701
rect 20809 22692 20821 22695
rect 20150 22664 20821 22692
rect 20150 22661 20162 22664
rect 20104 22655 20162 22661
rect 20809 22661 20821 22664
rect 20855 22661 20867 22695
rect 20809 22655 20867 22661
rect 24388 22695 24446 22701
rect 24388 22661 24400 22695
rect 24434 22692 24446 22695
rect 24578 22692 24584 22704
rect 24434 22664 24584 22692
rect 24434 22661 24446 22664
rect 24388 22655 24446 22661
rect 24578 22652 24584 22664
rect 24636 22652 24642 22704
rect 26513 22695 26571 22701
rect 26513 22661 26525 22695
rect 26559 22692 26571 22695
rect 26786 22692 26792 22704
rect 26559 22664 26792 22692
rect 26559 22661 26571 22664
rect 26513 22655 26571 22661
rect 26786 22652 26792 22664
rect 26844 22692 26850 22704
rect 27338 22692 27344 22704
rect 26844 22664 27344 22692
rect 26844 22652 26850 22664
rect 27338 22652 27344 22664
rect 27396 22652 27402 22704
rect 28261 22695 28319 22701
rect 28261 22661 28273 22695
rect 28307 22692 28319 22695
rect 28534 22692 28540 22704
rect 28307 22664 28540 22692
rect 28307 22661 28319 22664
rect 28261 22655 28319 22661
rect 28534 22652 28540 22664
rect 28592 22652 28598 22704
rect 29241 22695 29299 22701
rect 29241 22692 29253 22695
rect 29104 22664 29253 22692
rect 2590 22624 2596 22636
rect 2503 22596 2596 22624
rect 2590 22584 2596 22596
rect 2648 22624 2654 22636
rect 7558 22624 7564 22636
rect 2648 22596 7564 22624
rect 2648 22584 2654 22596
rect 7558 22584 7564 22596
rect 7616 22584 7622 22636
rect 10965 22627 11023 22633
rect 10965 22593 10977 22627
rect 11011 22624 11023 22627
rect 11422 22624 11428 22636
rect 11011 22596 11428 22624
rect 11011 22593 11023 22596
rect 10965 22587 11023 22593
rect 11422 22584 11428 22596
rect 11480 22584 11486 22636
rect 16298 22624 16304 22636
rect 16259 22596 16304 22624
rect 16298 22584 16304 22596
rect 16356 22584 16362 22636
rect 16390 22584 16396 22636
rect 16448 22624 16454 22636
rect 16853 22627 16911 22633
rect 16853 22624 16865 22627
rect 16448 22596 16865 22624
rect 16448 22584 16454 22596
rect 16853 22593 16865 22596
rect 16899 22593 16911 22627
rect 17034 22624 17040 22636
rect 16995 22596 17040 22624
rect 16853 22587 16911 22593
rect 17034 22584 17040 22596
rect 17092 22584 17098 22636
rect 20990 22624 20996 22636
rect 20951 22596 20996 22624
rect 20990 22584 20996 22596
rect 21048 22584 21054 22636
rect 21266 22624 21272 22636
rect 21227 22596 21272 22624
rect 21266 22584 21272 22596
rect 21324 22584 21330 22636
rect 22272 22627 22330 22633
rect 22272 22593 22284 22627
rect 22318 22624 22330 22627
rect 22554 22624 22560 22636
rect 22318 22596 22560 22624
rect 22318 22593 22330 22596
rect 22272 22587 22330 22593
rect 22554 22584 22560 22596
rect 22612 22584 22618 22636
rect 24118 22624 24124 22636
rect 24079 22596 24124 22624
rect 24118 22584 24124 22596
rect 24176 22584 24182 22636
rect 26421 22627 26479 22633
rect 26421 22593 26433 22627
rect 26467 22624 26479 22627
rect 26602 22624 26608 22636
rect 26467 22596 26608 22624
rect 26467 22593 26479 22596
rect 26421 22587 26479 22593
rect 26602 22584 26608 22596
rect 26660 22584 26666 22636
rect 27430 22624 27436 22636
rect 27391 22596 27436 22624
rect 27430 22584 27436 22596
rect 27488 22584 27494 22636
rect 27706 22584 27712 22636
rect 27764 22624 27770 22636
rect 28442 22624 28448 22636
rect 27764 22596 28448 22624
rect 27764 22584 27770 22596
rect 28442 22584 28448 22596
rect 28500 22624 28506 22636
rect 29104 22624 29132 22664
rect 29241 22661 29253 22664
rect 29287 22661 29299 22695
rect 29241 22655 29299 22661
rect 29457 22695 29515 22701
rect 29457 22661 29469 22695
rect 29503 22661 29515 22695
rect 29457 22655 29515 22661
rect 28500 22596 29132 22624
rect 28500 22584 28506 22596
rect 13078 22556 13084 22568
rect 13039 22528 13084 22556
rect 13078 22516 13084 22528
rect 13136 22516 13142 22568
rect 15562 22556 15568 22568
rect 15523 22528 15568 22556
rect 15562 22516 15568 22528
rect 15620 22516 15626 22568
rect 20346 22516 20352 22568
rect 20404 22556 20410 22568
rect 22002 22556 22008 22568
rect 20404 22528 20497 22556
rect 21963 22528 22008 22556
rect 20404 22516 20410 22528
rect 22002 22516 22008 22528
rect 22060 22516 22066 22568
rect 27338 22516 27344 22568
rect 27396 22556 27402 22568
rect 29472 22556 29500 22655
rect 30006 22652 30012 22704
rect 30064 22692 30070 22704
rect 30193 22695 30251 22701
rect 30193 22692 30205 22695
rect 30064 22664 30205 22692
rect 30064 22652 30070 22664
rect 30193 22661 30205 22664
rect 30239 22692 30251 22695
rect 32950 22692 32956 22704
rect 30239 22664 32956 22692
rect 30239 22661 30251 22664
rect 30193 22655 30251 22661
rect 30561 22627 30619 22633
rect 30561 22593 30573 22627
rect 30607 22624 30619 22627
rect 30834 22624 30840 22636
rect 30607 22596 30840 22624
rect 30607 22593 30619 22596
rect 30561 22587 30619 22593
rect 30834 22584 30840 22596
rect 30892 22584 30898 22636
rect 31294 22624 31300 22636
rect 31255 22596 31300 22624
rect 31294 22584 31300 22596
rect 31352 22584 31358 22636
rect 31496 22633 31524 22664
rect 32950 22652 32956 22664
rect 33008 22652 33014 22704
rect 33597 22695 33655 22701
rect 33597 22661 33609 22695
rect 33643 22692 33655 22695
rect 34146 22692 34152 22704
rect 33643 22664 34152 22692
rect 33643 22661 33655 22664
rect 33597 22655 33655 22661
rect 34146 22652 34152 22664
rect 34204 22652 34210 22704
rect 36354 22652 36360 22704
rect 36412 22692 36418 22704
rect 42812 22692 42840 22720
rect 43088 22701 43116 22732
rect 42982 22695 43040 22701
rect 42982 22692 42994 22695
rect 36412 22664 37688 22692
rect 42812 22664 42994 22692
rect 36412 22652 36418 22664
rect 31481 22627 31539 22633
rect 31481 22593 31493 22627
rect 31527 22593 31539 22627
rect 31481 22587 31539 22593
rect 31573 22627 31631 22633
rect 31573 22593 31585 22627
rect 31619 22624 31631 22627
rect 33778 22624 33784 22636
rect 31619 22596 33784 22624
rect 31619 22593 31631 22596
rect 31573 22587 31631 22593
rect 33778 22584 33784 22596
rect 33836 22584 33842 22636
rect 35618 22584 35624 22636
rect 35676 22624 35682 22636
rect 36265 22627 36323 22633
rect 36265 22624 36277 22627
rect 35676 22596 36277 22624
rect 35676 22584 35682 22596
rect 36265 22593 36277 22596
rect 36311 22593 36323 22627
rect 36265 22587 36323 22593
rect 36449 22627 36507 22633
rect 36449 22593 36461 22627
rect 36495 22624 36507 22627
rect 36722 22624 36728 22636
rect 36495 22596 36728 22624
rect 36495 22593 36507 22596
rect 36449 22587 36507 22593
rect 36722 22584 36728 22596
rect 36780 22584 36786 22636
rect 37660 22633 37688 22664
rect 42982 22661 42994 22664
rect 43028 22661 43040 22695
rect 43088 22695 43157 22701
rect 43088 22664 43111 22695
rect 42982 22655 43040 22661
rect 43099 22661 43111 22664
rect 43145 22661 43157 22695
rect 44174 22692 44180 22704
rect 43099 22655 43157 22661
rect 43272 22664 44180 22692
rect 37461 22627 37519 22633
rect 37461 22593 37473 22627
rect 37507 22593 37519 22627
rect 37461 22587 37519 22593
rect 37645 22627 37703 22633
rect 37645 22593 37657 22627
rect 37691 22593 37703 22627
rect 38930 22624 38936 22636
rect 38891 22596 38936 22624
rect 37645 22587 37703 22593
rect 27396 22528 29500 22556
rect 36357 22559 36415 22565
rect 27396 22516 27402 22528
rect 36357 22525 36369 22559
rect 36403 22556 36415 22559
rect 36814 22556 36820 22568
rect 36403 22528 36820 22556
rect 36403 22525 36415 22528
rect 36357 22519 36415 22525
rect 36814 22516 36820 22528
rect 36872 22556 36878 22568
rect 37476 22556 37504 22587
rect 38930 22584 38936 22596
rect 38988 22584 38994 22636
rect 39022 22584 39028 22636
rect 39080 22624 39086 22636
rect 39189 22627 39247 22633
rect 39189 22624 39201 22627
rect 39080 22596 39201 22624
rect 39080 22584 39086 22596
rect 39189 22593 39201 22596
rect 39235 22593 39247 22627
rect 39189 22587 39247 22593
rect 41782 22584 41788 22636
rect 41840 22624 41846 22636
rect 41877 22627 41935 22633
rect 41877 22624 41889 22627
rect 41840 22596 41889 22624
rect 41840 22584 41846 22596
rect 41877 22593 41889 22596
rect 41923 22593 41935 22627
rect 42794 22624 42800 22636
rect 42755 22596 42800 22624
rect 41877 22587 41935 22593
rect 41690 22556 41696 22568
rect 36872 22528 37504 22556
rect 41651 22528 41696 22556
rect 36872 22516 36878 22528
rect 41690 22516 41696 22528
rect 41748 22516 41754 22568
rect 41892 22556 41920 22587
rect 42794 22584 42800 22596
rect 42852 22584 42858 22636
rect 42889 22627 42947 22633
rect 42889 22593 42901 22627
rect 42935 22624 42947 22627
rect 43272 22624 43300 22664
rect 44174 22652 44180 22664
rect 44232 22652 44238 22704
rect 42935 22596 43300 22624
rect 43717 22627 43775 22633
rect 42935 22593 42947 22596
rect 42889 22587 42947 22593
rect 43717 22593 43729 22627
rect 43763 22593 43775 22627
rect 43898 22624 43904 22636
rect 43859 22596 43904 22624
rect 43717 22587 43775 22593
rect 43257 22559 43315 22565
rect 43257 22556 43269 22559
rect 41892 22528 43269 22556
rect 43257 22525 43269 22528
rect 43303 22556 43315 22559
rect 43732 22556 43760 22587
rect 43898 22584 43904 22596
rect 43956 22584 43962 22636
rect 43303 22528 43760 22556
rect 43303 22525 43315 22528
rect 43257 22519 43315 22525
rect 20364 22488 20392 22516
rect 20714 22488 20720 22500
rect 20364 22460 20720 22488
rect 20714 22448 20720 22460
rect 20772 22488 20778 22500
rect 22020 22488 22048 22516
rect 33410 22488 33416 22500
rect 20772 22460 22048 22488
rect 25056 22460 33416 22488
rect 20772 22448 20778 22460
rect 25056 22432 25084 22460
rect 33410 22448 33416 22460
rect 33468 22488 33474 22500
rect 34054 22488 34060 22500
rect 33468 22460 34060 22488
rect 33468 22448 33474 22460
rect 34054 22448 34060 22460
rect 34112 22448 34118 22500
rect 42061 22491 42119 22497
rect 42061 22457 42073 22491
rect 42107 22488 42119 22491
rect 42886 22488 42892 22500
rect 42107 22460 42892 22488
rect 42107 22457 42119 22460
rect 42061 22451 42119 22457
rect 42886 22448 42892 22460
rect 42944 22448 42950 22500
rect 43438 22448 43444 22500
rect 43496 22488 43502 22500
rect 44085 22491 44143 22497
rect 44085 22488 44097 22491
rect 43496 22460 44097 22488
rect 43496 22448 43502 22460
rect 44085 22457 44097 22460
rect 44131 22457 44143 22491
rect 44085 22451 44143 22457
rect 2501 22423 2559 22429
rect 2501 22389 2513 22423
rect 2547 22420 2559 22423
rect 3234 22420 3240 22432
rect 2547 22392 3240 22420
rect 2547 22389 2559 22392
rect 2501 22383 2559 22389
rect 3234 22380 3240 22392
rect 3292 22380 3298 22432
rect 16758 22380 16764 22432
rect 16816 22420 16822 22432
rect 17037 22423 17095 22429
rect 17037 22420 17049 22423
rect 16816 22392 17049 22420
rect 16816 22380 16822 22392
rect 17037 22389 17049 22392
rect 17083 22389 17095 22423
rect 18966 22420 18972 22432
rect 18927 22392 18972 22420
rect 17037 22383 17095 22389
rect 18966 22380 18972 22392
rect 19024 22380 19030 22432
rect 20438 22380 20444 22432
rect 20496 22420 20502 22432
rect 21177 22423 21235 22429
rect 21177 22420 21189 22423
rect 20496 22392 21189 22420
rect 20496 22380 20502 22392
rect 21177 22389 21189 22392
rect 21223 22389 21235 22423
rect 21177 22383 21235 22389
rect 25038 22380 25044 22432
rect 25096 22380 25102 22432
rect 25498 22420 25504 22432
rect 25459 22392 25504 22420
rect 25498 22380 25504 22392
rect 25556 22380 25562 22432
rect 28626 22420 28632 22432
rect 28587 22392 28632 22420
rect 28626 22380 28632 22392
rect 28684 22380 28690 22432
rect 29086 22420 29092 22432
rect 29047 22392 29092 22420
rect 29086 22380 29092 22392
rect 29144 22380 29150 22432
rect 29270 22420 29276 22432
rect 29231 22392 29276 22420
rect 29270 22380 29276 22392
rect 29328 22380 29334 22432
rect 31113 22423 31171 22429
rect 31113 22389 31125 22423
rect 31159 22420 31171 22423
rect 31202 22420 31208 22432
rect 31159 22392 31208 22420
rect 31159 22389 31171 22392
rect 31113 22383 31171 22389
rect 31202 22380 31208 22392
rect 31260 22380 31266 22432
rect 33965 22423 34023 22429
rect 33965 22389 33977 22423
rect 34011 22420 34023 22423
rect 34790 22420 34796 22432
rect 34011 22392 34796 22420
rect 34011 22389 34023 22392
rect 33965 22383 34023 22389
rect 34790 22380 34796 22392
rect 34848 22420 34854 22432
rect 35434 22420 35440 22432
rect 34848 22392 35440 22420
rect 34848 22380 34854 22392
rect 35434 22380 35440 22392
rect 35492 22380 35498 22432
rect 37366 22380 37372 22432
rect 37424 22420 37430 22432
rect 37553 22423 37611 22429
rect 37553 22420 37565 22423
rect 37424 22392 37565 22420
rect 37424 22380 37430 22392
rect 37553 22389 37565 22392
rect 37599 22389 37611 22423
rect 40310 22420 40316 22432
rect 40271 22392 40316 22420
rect 37553 22383 37611 22389
rect 40310 22380 40316 22392
rect 40368 22380 40374 22432
rect 42426 22380 42432 22432
rect 42484 22420 42490 22432
rect 42613 22423 42671 22429
rect 42613 22420 42625 22423
rect 42484 22392 42625 22420
rect 42484 22380 42490 22392
rect 42613 22389 42625 22392
rect 42659 22389 42671 22423
rect 42613 22383 42671 22389
rect 43254 22380 43260 22432
rect 43312 22420 43318 22432
rect 44266 22420 44272 22432
rect 43312 22392 44272 22420
rect 43312 22380 43318 22392
rect 44266 22380 44272 22392
rect 44324 22380 44330 22432
rect 47949 22423 48007 22429
rect 47949 22389 47961 22423
rect 47995 22420 48007 22423
rect 48314 22420 48320 22432
rect 47995 22392 48320 22420
rect 47995 22389 48007 22392
rect 47949 22383 48007 22389
rect 48314 22380 48320 22392
rect 48372 22380 48378 22432
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 14642 22216 14648 22228
rect 14603 22188 14648 22216
rect 14642 22176 14648 22188
rect 14700 22176 14706 22228
rect 16482 22176 16488 22228
rect 16540 22216 16546 22228
rect 18230 22216 18236 22228
rect 16540 22188 18236 22216
rect 16540 22176 16546 22188
rect 18230 22176 18236 22188
rect 18288 22176 18294 22228
rect 22554 22216 22560 22228
rect 22515 22188 22560 22216
rect 22554 22176 22560 22188
rect 22612 22176 22618 22228
rect 22646 22176 22652 22228
rect 22704 22216 22710 22228
rect 23201 22219 23259 22225
rect 23201 22216 23213 22219
rect 22704 22188 23213 22216
rect 22704 22176 22710 22188
rect 23201 22185 23213 22188
rect 23247 22185 23259 22219
rect 23201 22179 23259 22185
rect 24581 22219 24639 22225
rect 24581 22185 24593 22219
rect 24627 22216 24639 22219
rect 24762 22216 24768 22228
rect 24627 22188 24768 22216
rect 24627 22185 24639 22188
rect 24581 22179 24639 22185
rect 24762 22176 24768 22188
rect 24820 22176 24826 22228
rect 24854 22176 24860 22228
rect 24912 22176 24918 22228
rect 26605 22219 26663 22225
rect 26605 22185 26617 22219
rect 26651 22185 26663 22219
rect 26605 22179 26663 22185
rect 11606 22148 11612 22160
rect 11567 22120 11612 22148
rect 11606 22108 11612 22120
rect 11664 22108 11670 22160
rect 18322 22148 18328 22160
rect 18156 22120 18328 22148
rect 3234 22080 3240 22092
rect 3195 22052 3240 22080
rect 3234 22040 3240 22052
rect 3292 22040 3298 22092
rect 11422 22080 11428 22092
rect 11383 22052 11428 22080
rect 11422 22040 11428 22052
rect 11480 22040 11486 22092
rect 11882 22080 11888 22092
rect 11843 22052 11888 22080
rect 11882 22040 11888 22052
rect 11940 22040 11946 22092
rect 13078 22040 13084 22092
rect 13136 22080 13142 22092
rect 15562 22080 15568 22092
rect 13136 22052 15568 22080
rect 13136 22040 13142 22052
rect 15562 22040 15568 22052
rect 15620 22080 15626 22092
rect 16117 22083 16175 22089
rect 16117 22080 16129 22083
rect 15620 22052 16129 22080
rect 15620 22040 15626 22052
rect 16117 22049 16129 22052
rect 16163 22049 16175 22083
rect 16117 22043 16175 22049
rect 3418 21972 3424 22024
rect 3476 22012 3482 22024
rect 14458 22012 14464 22024
rect 3476 21984 3521 22012
rect 14419 21984 14464 22012
rect 3476 21972 3482 21984
rect 14458 21972 14464 21984
rect 14516 21972 14522 22024
rect 14734 22012 14740 22024
rect 14647 21984 14740 22012
rect 14734 21972 14740 21984
rect 14792 22012 14798 22024
rect 17862 22012 17868 22024
rect 14792 21984 17868 22012
rect 14792 21972 14798 21984
rect 17862 21972 17868 21984
rect 17920 21972 17926 22024
rect 18156 22021 18184 22120
rect 18322 22108 18328 22120
rect 18380 22108 18386 22160
rect 23842 22148 23848 22160
rect 23755 22120 23848 22148
rect 18966 22080 18972 22092
rect 18248 22052 18972 22080
rect 18248 22021 18276 22052
rect 18966 22040 18972 22052
rect 19024 22080 19030 22092
rect 20073 22083 20131 22089
rect 19024 22052 19472 22080
rect 19024 22040 19030 22052
rect 18141 22015 18199 22021
rect 18141 21981 18153 22015
rect 18187 21981 18199 22015
rect 18141 21975 18199 21981
rect 18233 22015 18291 22021
rect 18233 21981 18245 22015
rect 18279 21981 18291 22015
rect 18233 21975 18291 21981
rect 18322 21972 18328 22024
rect 18380 22012 18386 22024
rect 19444 22021 19472 22052
rect 20073 22049 20085 22083
rect 20119 22080 20131 22083
rect 20990 22080 20996 22092
rect 20119 22052 20996 22080
rect 20119 22049 20131 22052
rect 20073 22043 20131 22049
rect 20990 22040 20996 22052
rect 21048 22040 21054 22092
rect 22002 22080 22008 22092
rect 21915 22052 22008 22080
rect 22002 22040 22008 22052
rect 22060 22080 22066 22092
rect 23566 22080 23572 22092
rect 22060 22052 23572 22080
rect 22060 22040 22066 22052
rect 23566 22040 23572 22052
rect 23624 22040 23630 22092
rect 23768 22089 23796 22120
rect 23842 22108 23848 22120
rect 23900 22148 23906 22160
rect 24872 22148 24900 22176
rect 23900 22120 24900 22148
rect 26620 22148 26648 22179
rect 27246 22176 27252 22228
rect 27304 22216 27310 22228
rect 27430 22216 27436 22228
rect 27304 22188 27436 22216
rect 27304 22176 27310 22188
rect 27430 22176 27436 22188
rect 27488 22216 27494 22228
rect 27893 22219 27951 22225
rect 27893 22216 27905 22219
rect 27488 22188 27905 22216
rect 27488 22176 27494 22188
rect 27893 22185 27905 22188
rect 27939 22216 27951 22219
rect 32214 22216 32220 22228
rect 27939 22188 32220 22216
rect 27939 22185 27951 22188
rect 27893 22179 27951 22185
rect 32214 22176 32220 22188
rect 32272 22176 32278 22228
rect 32309 22219 32367 22225
rect 32309 22185 32321 22219
rect 32355 22216 32367 22219
rect 33778 22216 33784 22228
rect 32355 22188 33784 22216
rect 32355 22185 32367 22188
rect 32309 22179 32367 22185
rect 33778 22176 33784 22188
rect 33836 22176 33842 22228
rect 37734 22176 37740 22228
rect 37792 22216 37798 22228
rect 37829 22219 37887 22225
rect 37829 22216 37841 22219
rect 37792 22188 37841 22216
rect 37792 22176 37798 22188
rect 37829 22185 37841 22188
rect 37875 22185 37887 22219
rect 39022 22216 39028 22228
rect 38983 22188 39028 22216
rect 37829 22179 37887 22185
rect 39022 22176 39028 22188
rect 39080 22176 39086 22228
rect 41325 22219 41383 22225
rect 41325 22185 41337 22219
rect 41371 22216 41383 22219
rect 41782 22216 41788 22228
rect 41371 22188 41788 22216
rect 41371 22185 41383 22188
rect 41325 22179 41383 22185
rect 41782 22176 41788 22188
rect 41840 22176 41846 22228
rect 42886 22176 42892 22228
rect 42944 22216 42950 22228
rect 43162 22216 43168 22228
rect 42944 22188 43168 22216
rect 42944 22176 42950 22188
rect 43162 22176 43168 22188
rect 43220 22176 43226 22228
rect 43346 22176 43352 22228
rect 43404 22216 43410 22228
rect 43898 22216 43904 22228
rect 43404 22188 43904 22216
rect 43404 22176 43410 22188
rect 43898 22176 43904 22188
rect 43956 22176 43962 22228
rect 44174 22216 44180 22228
rect 44135 22188 44180 22216
rect 44174 22176 44180 22188
rect 44232 22176 44238 22228
rect 44266 22176 44272 22228
rect 44324 22216 44330 22228
rect 44324 22188 44369 22216
rect 44324 22176 44330 22188
rect 27706 22148 27712 22160
rect 26620 22120 27712 22148
rect 23900 22108 23906 22120
rect 27706 22108 27712 22120
rect 27764 22108 27770 22160
rect 43438 22148 43444 22160
rect 43399 22120 43444 22148
rect 43438 22108 43444 22120
rect 43496 22108 43502 22160
rect 43548 22120 44220 22148
rect 23753 22083 23811 22089
rect 23753 22049 23765 22083
rect 23799 22080 23811 22083
rect 23799 22052 23833 22080
rect 23799 22049 23811 22052
rect 23753 22043 23811 22049
rect 26510 22040 26516 22092
rect 26568 22080 26574 22092
rect 26568 22052 31064 22080
rect 26568 22040 26574 22052
rect 18509 22015 18567 22021
rect 18380 21984 18425 22012
rect 18380 21972 18386 21984
rect 18509 21981 18521 22015
rect 18555 21981 18567 22015
rect 18509 21975 18567 21981
rect 19429 22015 19487 22021
rect 19429 21981 19441 22015
rect 19475 21981 19487 22015
rect 19429 21975 19487 21981
rect 19613 22015 19671 22021
rect 19613 21981 19625 22015
rect 19659 21981 19671 22015
rect 19613 21975 19671 21981
rect 19889 22015 19947 22021
rect 19889 21981 19901 22015
rect 19935 22012 19947 22015
rect 22738 22012 22744 22024
rect 19935 21984 20116 22012
rect 22699 21984 22744 22012
rect 19935 21981 19947 21984
rect 19889 21975 19947 21981
rect 1578 21944 1584 21956
rect 1539 21916 1584 21944
rect 1578 21904 1584 21916
rect 1636 21904 1642 21956
rect 16384 21947 16442 21953
rect 16384 21913 16396 21947
rect 16430 21944 16442 21947
rect 16850 21944 16856 21956
rect 16430 21916 16856 21944
rect 16430 21913 16442 21916
rect 16384 21907 16442 21913
rect 16850 21904 16856 21916
rect 16908 21904 16914 21956
rect 17034 21904 17040 21956
rect 17092 21944 17098 21956
rect 18524 21944 18552 21975
rect 17092 21916 18552 21944
rect 19628 21944 19656 21975
rect 20088 21956 20116 21984
rect 22738 21972 22744 21984
rect 22796 21972 22802 22024
rect 23584 22012 23612 22040
rect 31036 22024 31064 22052
rect 33870 22040 33876 22092
rect 33928 22080 33934 22092
rect 36078 22080 36084 22092
rect 33928 22052 36084 22080
rect 33928 22040 33934 22052
rect 36078 22040 36084 22052
rect 36136 22040 36142 22092
rect 36354 22080 36360 22092
rect 36315 22052 36360 22080
rect 36354 22040 36360 22052
rect 36412 22040 36418 22092
rect 36814 22080 36820 22092
rect 36775 22052 36820 22080
rect 36814 22040 36820 22052
rect 36872 22040 36878 22092
rect 37366 22080 37372 22092
rect 37327 22052 37372 22080
rect 37366 22040 37372 22052
rect 37424 22040 37430 22092
rect 37918 22040 37924 22092
rect 37976 22080 37982 22092
rect 43162 22080 43168 22092
rect 37976 22052 38516 22080
rect 43123 22052 43168 22080
rect 37976 22040 37982 22052
rect 24118 22012 24124 22024
rect 23584 21984 24124 22012
rect 24118 21972 24124 21984
rect 24176 21972 24182 22024
rect 24670 21972 24676 22024
rect 24728 22012 24734 22024
rect 24765 22015 24823 22021
rect 24765 22012 24777 22015
rect 24728 21984 24777 22012
rect 24728 21972 24734 21984
rect 24765 21981 24777 21984
rect 24811 21981 24823 22015
rect 24765 21975 24823 21981
rect 24946 21972 24952 22024
rect 25004 22012 25010 22024
rect 25041 22015 25099 22021
rect 25041 22012 25053 22015
rect 25004 21984 25053 22012
rect 25004 21972 25010 21984
rect 25041 21981 25053 21984
rect 25087 21981 25099 22015
rect 25041 21975 25099 21981
rect 25225 22015 25283 22021
rect 25225 21981 25237 22015
rect 25271 22012 25283 22015
rect 25498 22012 25504 22024
rect 25271 21984 25504 22012
rect 25271 21981 25283 21984
rect 25225 21975 25283 21981
rect 25498 21972 25504 21984
rect 25556 21972 25562 22024
rect 26234 21972 26240 22024
rect 26292 22012 26298 22024
rect 26786 22012 26792 22024
rect 26292 21984 26792 22012
rect 26292 21972 26298 21984
rect 26786 21972 26792 21984
rect 26844 21972 26850 22024
rect 26973 22015 27031 22021
rect 26973 21981 26985 22015
rect 27019 22012 27031 22015
rect 27522 22012 27528 22024
rect 27019 21984 27528 22012
rect 27019 21981 27031 21984
rect 26973 21975 27031 21981
rect 27522 21972 27528 21984
rect 27580 21972 27586 22024
rect 27798 22012 27804 22024
rect 27759 21984 27804 22012
rect 27798 21972 27804 21984
rect 27856 21972 27862 22024
rect 28997 22015 29055 22021
rect 28997 21981 29009 22015
rect 29043 22012 29055 22015
rect 29086 22012 29092 22024
rect 29043 21984 29092 22012
rect 29043 21981 29055 21984
rect 28997 21975 29055 21981
rect 29086 21972 29092 21984
rect 29144 21972 29150 22024
rect 29914 22012 29920 22024
rect 29875 21984 29920 22012
rect 29914 21972 29920 21984
rect 29972 21972 29978 22024
rect 30098 22012 30104 22024
rect 30059 21984 30104 22012
rect 30098 21972 30104 21984
rect 30156 21972 30162 22024
rect 30193 22015 30251 22021
rect 30193 21981 30205 22015
rect 30239 22012 30251 22015
rect 30282 22012 30288 22024
rect 30239 21984 30288 22012
rect 30239 21981 30251 21984
rect 30193 21975 30251 21981
rect 30282 21972 30288 21984
rect 30340 21972 30346 22024
rect 30929 22015 30987 22021
rect 30929 21981 30941 22015
rect 30975 21981 30987 22015
rect 30929 21975 30987 21981
rect 19978 21944 19984 21956
rect 19628 21916 19984 21944
rect 17092 21904 17098 21916
rect 14274 21876 14280 21888
rect 14235 21848 14280 21876
rect 14274 21836 14280 21848
rect 14332 21836 14338 21888
rect 16574 21836 16580 21888
rect 16632 21876 16638 21888
rect 17052 21876 17080 21904
rect 17512 21885 17540 21916
rect 19978 21904 19984 21916
rect 20036 21904 20042 21956
rect 20070 21904 20076 21956
rect 20128 21904 20134 21956
rect 21174 21944 21180 21956
rect 21135 21916 21180 21944
rect 21174 21904 21180 21916
rect 21232 21944 21238 21956
rect 28902 21944 28908 21956
rect 21232 21916 28908 21944
rect 21232 21904 21238 21916
rect 28902 21904 28908 21916
rect 28960 21904 28966 21956
rect 29181 21947 29239 21953
rect 29181 21913 29193 21947
rect 29227 21944 29239 21947
rect 30834 21944 30840 21956
rect 29227 21916 30840 21944
rect 29227 21913 29239 21916
rect 29181 21907 29239 21913
rect 30834 21904 30840 21916
rect 30892 21904 30898 21956
rect 30944 21888 30972 21975
rect 31018 21972 31024 22024
rect 31076 21972 31082 22024
rect 31202 22021 31208 22024
rect 31196 21975 31208 22021
rect 31260 22012 31266 22024
rect 32769 22015 32827 22021
rect 31260 21984 31296 22012
rect 31202 21972 31208 21975
rect 31260 21972 31266 21984
rect 32769 21981 32781 22015
rect 32815 21981 32827 22015
rect 35250 22012 35256 22024
rect 35211 21984 35256 22012
rect 32769 21975 32827 21981
rect 16632 21848 17080 21876
rect 17497 21879 17555 21885
rect 16632 21836 16638 21848
rect 17497 21845 17509 21879
rect 17543 21845 17555 21879
rect 17497 21839 17555 21845
rect 17770 21836 17776 21888
rect 17828 21876 17834 21888
rect 17957 21879 18015 21885
rect 17957 21876 17969 21879
rect 17828 21848 17969 21876
rect 17828 21836 17834 21848
rect 17957 21845 17969 21848
rect 18003 21845 18015 21879
rect 17957 21839 18015 21845
rect 18230 21836 18236 21888
rect 18288 21876 18294 21888
rect 22278 21876 22284 21888
rect 18288 21848 22284 21876
rect 18288 21836 18294 21848
rect 22278 21836 22284 21848
rect 22336 21836 22342 21888
rect 22370 21836 22376 21888
rect 22428 21876 22434 21888
rect 23569 21879 23627 21885
rect 23569 21876 23581 21879
rect 22428 21848 23581 21876
rect 22428 21836 22434 21848
rect 23569 21845 23581 21848
rect 23615 21845 23627 21879
rect 23569 21839 23627 21845
rect 23658 21836 23664 21888
rect 23716 21876 23722 21888
rect 26418 21876 26424 21888
rect 23716 21848 23761 21876
rect 26379 21848 26424 21876
rect 23716 21836 23722 21848
rect 26418 21836 26424 21848
rect 26476 21836 26482 21888
rect 26602 21876 26608 21888
rect 26563 21848 26608 21876
rect 26602 21836 26608 21848
rect 26660 21836 26666 21888
rect 28074 21876 28080 21888
rect 28035 21848 28080 21876
rect 28074 21836 28080 21848
rect 28132 21836 28138 21888
rect 29733 21879 29791 21885
rect 29733 21845 29745 21879
rect 29779 21876 29791 21879
rect 29822 21876 29828 21888
rect 29779 21848 29828 21876
rect 29779 21845 29791 21848
rect 29733 21839 29791 21845
rect 29822 21836 29828 21848
rect 29880 21836 29886 21888
rect 30926 21876 30932 21888
rect 30839 21848 30932 21876
rect 30926 21836 30932 21848
rect 30984 21876 30990 21888
rect 31662 21876 31668 21888
rect 30984 21848 31668 21876
rect 30984 21836 30990 21848
rect 31662 21836 31668 21848
rect 31720 21876 31726 21888
rect 32784 21876 32812 21975
rect 35250 21972 35256 21984
rect 35308 21972 35314 22024
rect 35434 22012 35440 22024
rect 35395 21984 35440 22012
rect 35434 21972 35440 21984
rect 35492 21972 35498 22024
rect 36449 22015 36507 22021
rect 36449 21981 36461 22015
rect 36495 22012 36507 22015
rect 37461 22015 37519 22021
rect 37461 22012 37473 22015
rect 36495 21984 37473 22012
rect 36495 21981 36507 21984
rect 36449 21975 36507 21981
rect 37461 21981 37473 21984
rect 37507 21981 37519 22015
rect 38286 22012 38292 22024
rect 38247 21984 38292 22012
rect 37461 21975 37519 21981
rect 33036 21947 33094 21953
rect 33036 21913 33048 21947
rect 33082 21944 33094 21947
rect 33318 21944 33324 21956
rect 33082 21916 33324 21944
rect 33082 21913 33094 21916
rect 33036 21907 33094 21913
rect 33318 21904 33324 21916
rect 33376 21904 33382 21956
rect 35345 21947 35403 21953
rect 35345 21913 35357 21947
rect 35391 21944 35403 21947
rect 35618 21944 35624 21956
rect 35391 21916 35624 21944
rect 35391 21913 35403 21916
rect 35345 21907 35403 21913
rect 35618 21904 35624 21916
rect 35676 21904 35682 21956
rect 37476 21944 37504 21975
rect 38286 21972 38292 21984
rect 38344 21972 38350 22024
rect 38488 22021 38516 22052
rect 43162 22040 43168 22052
rect 43220 22040 43226 22092
rect 38473 22015 38531 22021
rect 38473 21981 38485 22015
rect 38519 21981 38531 22015
rect 39206 22012 39212 22024
rect 39167 21984 39212 22012
rect 38473 21975 38531 21981
rect 39206 21972 39212 21984
rect 39264 21972 39270 22024
rect 39482 22012 39488 22024
rect 39443 21984 39488 22012
rect 39482 21972 39488 21984
rect 39540 21972 39546 22024
rect 40310 21972 40316 22024
rect 40368 22012 40374 22024
rect 40405 22015 40463 22021
rect 40405 22012 40417 22015
rect 40368 21984 40417 22012
rect 40368 21972 40374 21984
rect 40405 21981 40417 21984
rect 40451 21981 40463 22015
rect 41874 22012 41880 22024
rect 40405 21975 40463 21981
rect 41386 21984 41880 22012
rect 38381 21947 38439 21953
rect 38381 21944 38393 21947
rect 37476 21916 38393 21944
rect 38381 21913 38393 21916
rect 38427 21913 38439 21947
rect 38381 21907 38439 21913
rect 40773 21947 40831 21953
rect 40773 21913 40785 21947
rect 40819 21944 40831 21947
rect 41386 21944 41414 21984
rect 41874 21972 41880 21984
rect 41932 21972 41938 22024
rect 42426 22012 42432 22024
rect 42484 22021 42490 22024
rect 42396 21984 42432 22012
rect 42426 21972 42432 21984
rect 42484 21975 42496 22021
rect 42702 22012 42708 22024
rect 42663 21984 42708 22012
rect 42484 21972 42490 21975
rect 42702 21972 42708 21984
rect 42760 21972 42766 22024
rect 43070 21972 43076 22024
rect 43128 22012 43134 22024
rect 43548 22012 43576 22120
rect 44085 22083 44143 22089
rect 44085 22080 44097 22083
rect 43128 21984 43576 22012
rect 43640 22052 44097 22080
rect 43128 21972 43134 21984
rect 40819 21916 41414 21944
rect 40819 21913 40831 21916
rect 40773 21907 40831 21913
rect 41690 21904 41696 21956
rect 41748 21944 41754 21956
rect 43346 21944 43352 21956
rect 41748 21916 43352 21944
rect 41748 21904 41754 21916
rect 43346 21904 43352 21916
rect 43404 21904 43410 21956
rect 34146 21876 34152 21888
rect 31720 21848 32812 21876
rect 34107 21848 34152 21876
rect 31720 21836 31726 21848
rect 34146 21836 34152 21848
rect 34204 21836 34210 21888
rect 35526 21836 35532 21888
rect 35584 21876 35590 21888
rect 36173 21879 36231 21885
rect 36173 21876 36185 21879
rect 35584 21848 36185 21876
rect 35584 21836 35590 21848
rect 36173 21845 36185 21848
rect 36219 21845 36231 21879
rect 36173 21839 36231 21845
rect 39393 21879 39451 21885
rect 39393 21845 39405 21879
rect 39439 21876 39451 21879
rect 40954 21876 40960 21888
rect 39439 21848 40960 21876
rect 39439 21845 39451 21848
rect 39393 21839 39451 21845
rect 40954 21836 40960 21848
rect 41012 21876 41018 21888
rect 41708 21876 41736 21904
rect 43640 21888 43668 22052
rect 44085 22049 44097 22052
rect 44131 22049 44143 22083
rect 44192 22080 44220 22120
rect 46842 22080 46848 22092
rect 44192 22052 44404 22080
rect 46803 22052 46848 22080
rect 44085 22043 44143 22049
rect 44376 22021 44404 22052
rect 46842 22040 46848 22052
rect 46900 22040 46906 22092
rect 48314 22080 48320 22092
rect 48275 22052 48320 22080
rect 48314 22040 48320 22052
rect 48372 22040 48378 22092
rect 44361 22015 44419 22021
rect 44361 21981 44373 22015
rect 44407 21981 44419 22015
rect 44361 21975 44419 21981
rect 47854 21904 47860 21956
rect 47912 21944 47918 21956
rect 48133 21947 48191 21953
rect 48133 21944 48145 21947
rect 47912 21916 48145 21944
rect 47912 21904 47918 21916
rect 48133 21913 48145 21916
rect 48179 21913 48191 21947
rect 48133 21907 48191 21913
rect 43622 21876 43628 21888
rect 41012 21848 41736 21876
rect 43583 21848 43628 21876
rect 41012 21836 41018 21848
rect 43622 21836 43628 21848
rect 43680 21836 43686 21888
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 11882 21632 11888 21684
rect 11940 21672 11946 21684
rect 22281 21675 22339 21681
rect 11940 21644 22094 21672
rect 11940 21632 11946 21644
rect 13532 21607 13590 21613
rect 13532 21573 13544 21607
rect 13578 21604 13590 21607
rect 14274 21604 14280 21616
rect 13578 21576 14280 21604
rect 13578 21573 13590 21576
rect 13532 21567 13590 21573
rect 14274 21564 14280 21576
rect 14332 21564 14338 21616
rect 16301 21607 16359 21613
rect 16301 21573 16313 21607
rect 16347 21604 16359 21607
rect 16942 21604 16948 21616
rect 16347 21576 16948 21604
rect 16347 21573 16359 21576
rect 16301 21567 16359 21573
rect 16942 21564 16948 21576
rect 17000 21604 17006 21616
rect 17000 21576 17908 21604
rect 17000 21564 17006 21576
rect 2317 21539 2375 21545
rect 2317 21505 2329 21539
rect 2363 21536 2375 21539
rect 3418 21536 3424 21548
rect 2363 21508 3424 21536
rect 2363 21505 2375 21508
rect 2317 21499 2375 21505
rect 3418 21496 3424 21508
rect 3476 21496 3482 21548
rect 13078 21496 13084 21548
rect 13136 21536 13142 21548
rect 13265 21539 13323 21545
rect 13265 21536 13277 21539
rect 13136 21508 13277 21536
rect 13136 21496 13142 21508
rect 13265 21505 13277 21508
rect 13311 21505 13323 21539
rect 13265 21499 13323 21505
rect 16117 21539 16175 21545
rect 16117 21505 16129 21539
rect 16163 21536 16175 21539
rect 16574 21536 16580 21548
rect 16163 21508 16580 21536
rect 16163 21505 16175 21508
rect 16117 21499 16175 21505
rect 16574 21496 16580 21508
rect 16632 21496 16638 21548
rect 17218 21536 17224 21548
rect 17179 21508 17224 21536
rect 17218 21496 17224 21508
rect 17276 21496 17282 21548
rect 17313 21539 17371 21545
rect 17313 21505 17325 21539
rect 17359 21536 17371 21539
rect 17770 21536 17776 21548
rect 17359 21508 17776 21536
rect 17359 21505 17371 21508
rect 17313 21499 17371 21505
rect 17770 21496 17776 21508
rect 17828 21496 17834 21548
rect 17880 21545 17908 21576
rect 17954 21564 17960 21616
rect 18012 21604 18018 21616
rect 21266 21604 21272 21616
rect 18012 21576 21272 21604
rect 18012 21564 18018 21576
rect 21266 21564 21272 21576
rect 21324 21564 21330 21616
rect 17865 21539 17923 21545
rect 17865 21505 17877 21539
rect 17911 21505 17923 21539
rect 18233 21539 18291 21545
rect 18233 21536 18245 21539
rect 17865 21499 17923 21505
rect 17972 21508 18245 21536
rect 15933 21471 15991 21477
rect 15933 21468 15945 21471
rect 14660 21440 15945 21468
rect 14660 21409 14688 21440
rect 15933 21437 15945 21440
rect 15979 21468 15991 21471
rect 16390 21468 16396 21480
rect 15979 21440 16396 21468
rect 15979 21437 15991 21440
rect 15933 21431 15991 21437
rect 16390 21428 16396 21440
rect 16448 21428 16454 21480
rect 16850 21468 16856 21480
rect 16811 21440 16856 21468
rect 16850 21428 16856 21440
rect 16908 21428 16914 21480
rect 17034 21468 17040 21480
rect 16995 21440 17040 21468
rect 17034 21428 17040 21440
rect 17092 21428 17098 21480
rect 17129 21471 17187 21477
rect 17129 21437 17141 21471
rect 17175 21437 17187 21471
rect 17236 21468 17264 21496
rect 17494 21468 17500 21480
rect 17236 21440 17500 21468
rect 17129 21431 17187 21437
rect 14645 21403 14703 21409
rect 14645 21369 14657 21403
rect 14691 21369 14703 21403
rect 17144 21400 17172 21431
rect 17494 21428 17500 21440
rect 17552 21428 17558 21480
rect 17586 21428 17592 21480
rect 17644 21468 17650 21480
rect 17972 21468 18000 21508
rect 18233 21505 18245 21508
rect 18279 21505 18291 21539
rect 22066 21536 22094 21644
rect 22281 21641 22293 21675
rect 22327 21672 22339 21675
rect 22370 21672 22376 21684
rect 22327 21644 22376 21672
rect 22327 21641 22339 21644
rect 22281 21635 22339 21641
rect 22370 21632 22376 21644
rect 22428 21632 22434 21684
rect 23106 21632 23112 21684
rect 23164 21672 23170 21684
rect 24946 21672 24952 21684
rect 23164 21644 24952 21672
rect 23164 21632 23170 21644
rect 24946 21632 24952 21644
rect 25004 21672 25010 21684
rect 26234 21672 26240 21684
rect 25004 21644 26240 21672
rect 25004 21632 25010 21644
rect 26234 21632 26240 21644
rect 26292 21632 26298 21684
rect 26513 21675 26571 21681
rect 26513 21641 26525 21675
rect 26559 21672 26571 21675
rect 26559 21644 26740 21672
rect 26559 21641 26571 21644
rect 26513 21635 26571 21641
rect 26712 21616 26740 21644
rect 29730 21632 29736 21684
rect 29788 21672 29794 21684
rect 30282 21672 30288 21684
rect 29788 21644 30288 21672
rect 29788 21632 29794 21644
rect 30282 21632 30288 21644
rect 30340 21632 30346 21684
rect 33134 21672 33140 21684
rect 32876 21644 33140 21672
rect 23416 21607 23474 21613
rect 23416 21573 23428 21607
rect 23462 21604 23474 21607
rect 24121 21607 24179 21613
rect 24121 21604 24133 21607
rect 23462 21576 24133 21604
rect 23462 21573 23474 21576
rect 23416 21567 23474 21573
rect 24121 21573 24133 21576
rect 24167 21573 24179 21607
rect 24121 21567 24179 21573
rect 25501 21607 25559 21613
rect 25501 21573 25513 21607
rect 25547 21604 25559 21607
rect 25547 21576 26648 21604
rect 25547 21573 25559 21576
rect 25501 21567 25559 21573
rect 22066 21508 23612 21536
rect 18233 21499 18291 21505
rect 18138 21468 18144 21480
rect 17644 21440 18000 21468
rect 18099 21440 18144 21468
rect 17644 21428 17650 21440
rect 18138 21428 18144 21440
rect 18196 21428 18202 21480
rect 23584 21468 23612 21508
rect 23658 21496 23664 21548
rect 23716 21536 23722 21548
rect 24302 21536 24308 21548
rect 23716 21508 23761 21536
rect 24263 21508 24308 21536
rect 23716 21496 23722 21508
rect 24302 21496 24308 21508
rect 24360 21496 24366 21548
rect 24581 21539 24639 21545
rect 24581 21505 24593 21539
rect 24627 21536 24639 21539
rect 25038 21536 25044 21548
rect 24627 21508 25044 21536
rect 24627 21505 24639 21508
rect 24581 21499 24639 21505
rect 25038 21496 25044 21508
rect 25096 21496 25102 21548
rect 26329 21539 26387 21545
rect 26329 21505 26341 21539
rect 26375 21536 26387 21539
rect 26418 21536 26424 21548
rect 26375 21508 26424 21536
rect 26375 21505 26387 21508
rect 26329 21499 26387 21505
rect 26418 21496 26424 21508
rect 26476 21496 26482 21548
rect 25225 21471 25283 21477
rect 25225 21468 25237 21471
rect 23584 21440 25237 21468
rect 25225 21437 25237 21440
rect 25271 21468 25283 21471
rect 26510 21468 26516 21480
rect 25271 21440 26516 21468
rect 25271 21437 25283 21440
rect 25225 21431 25283 21437
rect 26510 21428 26516 21440
rect 26568 21428 26574 21480
rect 26620 21468 26648 21576
rect 26694 21564 26700 21616
rect 26752 21564 26758 21616
rect 27062 21564 27068 21616
rect 27120 21604 27126 21616
rect 27246 21604 27252 21616
rect 27120 21576 27252 21604
rect 27120 21564 27126 21576
rect 27246 21564 27252 21576
rect 27304 21604 27310 21616
rect 27433 21607 27491 21613
rect 27433 21604 27445 21607
rect 27304 21576 27445 21604
rect 27304 21564 27310 21576
rect 27433 21573 27445 21576
rect 27479 21573 27491 21607
rect 27433 21567 27491 21573
rect 27617 21607 27675 21613
rect 27617 21573 27629 21607
rect 27663 21573 27675 21607
rect 27617 21567 27675 21573
rect 27338 21496 27344 21548
rect 27396 21536 27402 21548
rect 27632 21536 27660 21567
rect 28626 21564 28632 21616
rect 28684 21604 28690 21616
rect 28721 21607 28779 21613
rect 28721 21604 28733 21607
rect 28684 21576 28733 21604
rect 28684 21564 28690 21576
rect 28721 21573 28733 21576
rect 28767 21573 28779 21607
rect 30926 21604 30932 21616
rect 28721 21567 28779 21573
rect 29564 21576 30932 21604
rect 29564 21545 29592 21576
rect 30926 21564 30932 21576
rect 30984 21564 30990 21616
rect 31389 21607 31447 21613
rect 31389 21573 31401 21607
rect 31435 21604 31447 21607
rect 32490 21604 32496 21616
rect 31435 21576 32496 21604
rect 31435 21573 31447 21576
rect 31389 21567 31447 21573
rect 32490 21564 32496 21576
rect 32548 21564 32554 21616
rect 29822 21545 29828 21548
rect 27396 21508 27660 21536
rect 29549 21539 29607 21545
rect 27396 21496 27402 21508
rect 29549 21505 29561 21539
rect 29595 21505 29607 21539
rect 29816 21536 29828 21545
rect 29783 21508 29828 21536
rect 29549 21499 29607 21505
rect 29816 21499 29828 21508
rect 29822 21496 29828 21499
rect 29880 21496 29886 21548
rect 32876 21545 32904 21644
rect 33134 21632 33140 21644
rect 33192 21632 33198 21684
rect 33318 21672 33324 21684
rect 33279 21644 33324 21672
rect 33318 21632 33324 21644
rect 33376 21632 33382 21684
rect 33873 21675 33931 21681
rect 33873 21641 33885 21675
rect 33919 21672 33931 21675
rect 35250 21672 35256 21684
rect 33919 21644 35256 21672
rect 33919 21641 33931 21644
rect 33873 21635 33931 21641
rect 35250 21632 35256 21644
rect 35308 21632 35314 21684
rect 37829 21675 37887 21681
rect 37829 21641 37841 21675
rect 37875 21672 37887 21675
rect 38286 21672 38292 21684
rect 37875 21644 38292 21672
rect 37875 21641 37887 21644
rect 37829 21635 37887 21641
rect 38286 21632 38292 21644
rect 38344 21632 38350 21684
rect 42613 21675 42671 21681
rect 42613 21641 42625 21675
rect 42659 21672 42671 21675
rect 42794 21672 42800 21684
rect 42659 21644 42800 21672
rect 42659 21641 42671 21644
rect 42613 21635 42671 21641
rect 42794 21632 42800 21644
rect 42852 21632 42858 21684
rect 43346 21632 43352 21684
rect 43404 21672 43410 21684
rect 45281 21675 45339 21681
rect 45281 21672 45293 21675
rect 43404 21644 45293 21672
rect 43404 21632 43410 21644
rect 45281 21641 45293 21644
rect 45327 21641 45339 21675
rect 47854 21672 47860 21684
rect 47815 21644 47860 21672
rect 45281 21635 45339 21641
rect 47854 21632 47860 21644
rect 47912 21632 47918 21684
rect 34146 21604 34152 21616
rect 33152 21576 34152 21604
rect 33152 21545 33180 21576
rect 31573 21539 31631 21545
rect 31573 21505 31585 21539
rect 31619 21505 31631 21539
rect 31573 21499 31631 21505
rect 31757 21539 31815 21545
rect 31757 21505 31769 21539
rect 31803 21536 31815 21539
rect 32585 21539 32643 21545
rect 32585 21536 32597 21539
rect 31803 21508 32597 21536
rect 31803 21505 31815 21508
rect 31757 21499 31815 21505
rect 32585 21505 32597 21508
rect 32631 21505 32643 21539
rect 32585 21499 32643 21505
rect 32769 21539 32827 21545
rect 32769 21505 32781 21539
rect 32815 21505 32827 21539
rect 32769 21499 32827 21505
rect 32861 21539 32919 21545
rect 32861 21505 32873 21539
rect 32907 21505 32919 21539
rect 32861 21499 32919 21505
rect 33137 21539 33195 21545
rect 33137 21505 33149 21539
rect 33183 21505 33195 21539
rect 33778 21536 33784 21548
rect 33739 21508 33784 21536
rect 33137 21499 33195 21505
rect 27706 21468 27712 21480
rect 26620 21440 27712 21468
rect 27706 21428 27712 21440
rect 27764 21428 27770 21480
rect 18049 21403 18107 21409
rect 18049 21400 18061 21403
rect 17144 21372 18061 21400
rect 14645 21363 14703 21369
rect 18049 21369 18061 21372
rect 18095 21369 18107 21403
rect 18049 21363 18107 21369
rect 22066 21372 22416 21400
rect 17862 21292 17868 21344
rect 17920 21332 17926 21344
rect 17957 21335 18015 21341
rect 17957 21332 17969 21335
rect 17920 21304 17969 21332
rect 17920 21292 17926 21304
rect 17957 21301 17969 21304
rect 18003 21301 18015 21335
rect 17957 21295 18015 21301
rect 20438 21292 20444 21344
rect 20496 21332 20502 21344
rect 22066 21332 22094 21372
rect 20496 21304 22094 21332
rect 22388 21332 22416 21372
rect 26326 21360 26332 21412
rect 26384 21400 26390 21412
rect 27249 21403 27307 21409
rect 27249 21400 27261 21403
rect 26384 21372 27261 21400
rect 26384 21360 26390 21372
rect 27249 21369 27261 21372
rect 27295 21369 27307 21403
rect 28902 21400 28908 21412
rect 27249 21363 27307 21369
rect 27356 21372 28764 21400
rect 28863 21372 28908 21400
rect 24489 21335 24547 21341
rect 24489 21332 24501 21335
rect 22388 21304 24501 21332
rect 20496 21292 20502 21304
rect 24489 21301 24501 21304
rect 24535 21301 24547 21335
rect 24489 21295 24547 21301
rect 24670 21292 24676 21344
rect 24728 21332 24734 21344
rect 27356 21332 27384 21372
rect 24728 21304 27384 21332
rect 27433 21335 27491 21341
rect 24728 21292 24734 21304
rect 27433 21301 27445 21335
rect 27479 21332 27491 21335
rect 27522 21332 27528 21344
rect 27479 21304 27528 21332
rect 27479 21301 27491 21304
rect 27433 21295 27491 21301
rect 27522 21292 27528 21304
rect 27580 21292 27586 21344
rect 28736 21332 28764 21372
rect 28902 21360 28908 21372
rect 28960 21360 28966 21412
rect 30650 21360 30656 21412
rect 30708 21400 30714 21412
rect 30929 21403 30987 21409
rect 30929 21400 30941 21403
rect 30708 21372 30941 21400
rect 30708 21360 30714 21372
rect 30929 21369 30941 21372
rect 30975 21400 30987 21403
rect 31588 21400 31616 21499
rect 30975 21372 31616 21400
rect 32784 21400 32812 21499
rect 33778 21496 33784 21508
rect 33836 21496 33842 21548
rect 33980 21545 34008 21576
rect 34146 21564 34152 21576
rect 34204 21564 34210 21616
rect 35268 21604 35296 21632
rect 35268 21576 36400 21604
rect 33965 21539 34023 21545
rect 33965 21505 33977 21539
rect 34011 21505 34023 21539
rect 35526 21536 35532 21548
rect 35487 21508 35532 21536
rect 33965 21499 34023 21505
rect 35526 21496 35532 21508
rect 35584 21496 35590 21548
rect 36372 21545 36400 21576
rect 36357 21539 36415 21545
rect 36357 21505 36369 21539
rect 36403 21505 36415 21539
rect 36357 21499 36415 21505
rect 36541 21539 36599 21545
rect 36541 21505 36553 21539
rect 36587 21536 36599 21539
rect 36814 21536 36820 21548
rect 36587 21508 36820 21536
rect 36587 21505 36599 21508
rect 36541 21499 36599 21505
rect 36814 21496 36820 21508
rect 36872 21496 36878 21548
rect 36906 21496 36912 21548
rect 36964 21536 36970 21548
rect 37645 21539 37703 21545
rect 37645 21536 37657 21539
rect 36964 21508 37657 21536
rect 36964 21496 36970 21508
rect 37645 21505 37657 21508
rect 37691 21505 37703 21539
rect 37918 21536 37924 21548
rect 37879 21508 37924 21536
rect 37645 21499 37703 21505
rect 37918 21496 37924 21508
rect 37976 21496 37982 21548
rect 42981 21539 43039 21545
rect 42981 21505 42993 21539
rect 43027 21536 43039 21539
rect 43622 21536 43628 21548
rect 43027 21508 43628 21536
rect 43027 21505 43039 21508
rect 42981 21499 43039 21505
rect 43622 21496 43628 21508
rect 43680 21496 43686 21548
rect 44453 21539 44511 21545
rect 44453 21505 44465 21539
rect 44499 21536 44511 21539
rect 44634 21536 44640 21548
rect 44499 21508 44640 21536
rect 44499 21505 44511 21508
rect 44453 21499 44511 21505
rect 44634 21496 44640 21508
rect 44692 21536 44698 21548
rect 45097 21539 45155 21545
rect 45097 21536 45109 21539
rect 44692 21508 45109 21536
rect 44692 21496 44698 21508
rect 45097 21505 45109 21508
rect 45143 21505 45155 21539
rect 46382 21536 46388 21548
rect 46343 21508 46388 21536
rect 45097 21499 45155 21505
rect 46382 21496 46388 21508
rect 46440 21536 46446 21548
rect 47578 21536 47584 21548
rect 46440 21508 47584 21536
rect 46440 21496 46446 21508
rect 47578 21496 47584 21508
rect 47636 21496 47642 21548
rect 47762 21536 47768 21548
rect 47723 21508 47768 21536
rect 47762 21496 47768 21508
rect 47820 21496 47826 21548
rect 32953 21471 33011 21477
rect 32953 21437 32965 21471
rect 32999 21468 33011 21471
rect 33870 21468 33876 21480
rect 32999 21440 33876 21468
rect 32999 21437 33011 21440
rect 32953 21431 33011 21437
rect 33870 21428 33876 21440
rect 33928 21428 33934 21480
rect 35618 21468 35624 21480
rect 35579 21440 35624 21468
rect 35618 21428 35624 21440
rect 35676 21428 35682 21480
rect 42886 21468 42892 21480
rect 42847 21440 42892 21468
rect 42886 21428 42892 21440
rect 42944 21468 42950 21480
rect 43070 21468 43076 21480
rect 42944 21440 43076 21468
rect 42944 21428 42950 21440
rect 43070 21428 43076 21440
rect 43128 21428 43134 21480
rect 44361 21471 44419 21477
rect 44361 21437 44373 21471
rect 44407 21468 44419 21471
rect 44407 21440 44496 21468
rect 44407 21437 44419 21440
rect 44361 21431 44419 21437
rect 44468 21412 44496 21440
rect 35161 21403 35219 21409
rect 35161 21400 35173 21403
rect 32784 21372 35173 21400
rect 30975 21369 30987 21372
rect 30929 21363 30987 21369
rect 35161 21369 35173 21372
rect 35207 21369 35219 21403
rect 39206 21400 39212 21412
rect 35161 21363 35219 21369
rect 35452 21372 39212 21400
rect 30742 21332 30748 21344
rect 28736 21304 30748 21332
rect 30742 21292 30748 21304
rect 30800 21292 30806 21344
rect 31018 21292 31024 21344
rect 31076 21332 31082 21344
rect 35452 21332 35480 21372
rect 39206 21360 39212 21372
rect 39264 21360 39270 21412
rect 43990 21360 43996 21412
rect 44048 21400 44054 21412
rect 44085 21403 44143 21409
rect 44085 21400 44097 21403
rect 44048 21372 44097 21400
rect 44048 21360 44054 21372
rect 44085 21369 44097 21372
rect 44131 21369 44143 21403
rect 44085 21363 44143 21369
rect 44450 21360 44456 21412
rect 44508 21360 44514 21412
rect 31076 21304 35480 21332
rect 31076 21292 31082 21304
rect 35986 21292 35992 21344
rect 36044 21332 36050 21344
rect 36173 21335 36231 21341
rect 36173 21332 36185 21335
rect 36044 21304 36185 21332
rect 36044 21292 36050 21304
rect 36173 21301 36185 21304
rect 36219 21301 36231 21335
rect 36173 21295 36231 21301
rect 37461 21335 37519 21341
rect 37461 21301 37473 21335
rect 37507 21332 37519 21335
rect 37550 21332 37556 21344
rect 37507 21304 37556 21332
rect 37507 21301 37519 21304
rect 37461 21295 37519 21301
rect 37550 21292 37556 21304
rect 37608 21292 37614 21344
rect 42794 21332 42800 21344
rect 42755 21304 42800 21332
rect 42794 21292 42800 21304
rect 42852 21332 42858 21344
rect 43254 21332 43260 21344
rect 42852 21304 43260 21332
rect 42852 21292 42858 21304
rect 43254 21292 43260 21304
rect 43312 21292 43318 21344
rect 46477 21335 46535 21341
rect 46477 21301 46489 21335
rect 46523 21332 46535 21335
rect 46658 21332 46664 21344
rect 46523 21304 46664 21332
rect 46523 21301 46535 21304
rect 46477 21295 46535 21301
rect 46658 21292 46664 21304
rect 46716 21292 46722 21344
rect 47026 21332 47032 21344
rect 46987 21304 47032 21332
rect 47026 21292 47032 21304
rect 47084 21292 47090 21344
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 14277 21131 14335 21137
rect 14277 21097 14289 21131
rect 14323 21128 14335 21131
rect 14458 21128 14464 21140
rect 14323 21100 14464 21128
rect 14323 21097 14335 21100
rect 14277 21091 14335 21097
rect 14458 21088 14464 21100
rect 14516 21088 14522 21140
rect 14918 21128 14924 21140
rect 14660 21100 14924 21128
rect 13814 20952 13820 21004
rect 13872 20992 13878 21004
rect 14660 20992 14688 21100
rect 14918 21088 14924 21100
rect 14976 21128 14982 21140
rect 19981 21131 20039 21137
rect 14976 21100 18000 21128
rect 14976 21088 14982 21100
rect 17034 21020 17040 21072
rect 17092 21060 17098 21072
rect 17313 21063 17371 21069
rect 17313 21060 17325 21063
rect 17092 21032 17325 21060
rect 17092 21020 17098 21032
rect 17313 21029 17325 21032
rect 17359 21029 17371 21063
rect 17313 21023 17371 21029
rect 17862 20992 17868 21004
rect 13872 20964 14688 20992
rect 13872 20952 13878 20964
rect 2038 20884 2044 20936
rect 2096 20924 2102 20936
rect 2133 20927 2191 20933
rect 2133 20924 2145 20927
rect 2096 20896 2145 20924
rect 2096 20884 2102 20896
rect 2133 20893 2145 20896
rect 2179 20893 2191 20927
rect 2133 20887 2191 20893
rect 14461 20927 14519 20933
rect 14461 20893 14473 20927
rect 14507 20924 14519 20927
rect 14550 20924 14556 20936
rect 14507 20896 14556 20924
rect 14507 20893 14519 20896
rect 14461 20887 14519 20893
rect 14550 20884 14556 20896
rect 14608 20884 14614 20936
rect 14660 20924 14688 20964
rect 14936 20964 16344 20992
rect 14936 20933 14964 20964
rect 16316 20933 16344 20964
rect 16776 20964 17868 20992
rect 16776 20936 16804 20964
rect 17862 20952 17868 20964
rect 17920 20952 17926 21004
rect 17972 20992 18000 21100
rect 19981 21097 19993 21131
rect 20027 21128 20039 21131
rect 20070 21128 20076 21140
rect 20027 21100 20076 21128
rect 20027 21097 20039 21100
rect 19981 21091 20039 21097
rect 20070 21088 20076 21100
rect 20128 21128 20134 21140
rect 20438 21128 20444 21140
rect 20128 21100 20444 21128
rect 20128 21088 20134 21100
rect 20438 21088 20444 21100
rect 20496 21088 20502 21140
rect 23569 21131 23627 21137
rect 23216 21100 23428 21128
rect 23106 21060 23112 21072
rect 21376 21032 23112 21060
rect 21376 20992 21404 21032
rect 23106 21020 23112 21032
rect 23164 21020 23170 21072
rect 23216 20992 23244 21100
rect 17972 20964 21404 20992
rect 22066 20964 23244 20992
rect 23400 20992 23428 21100
rect 23569 21097 23581 21131
rect 23615 21128 23627 21131
rect 24302 21128 24308 21140
rect 23615 21100 24308 21128
rect 23615 21097 23627 21100
rect 23569 21091 23627 21097
rect 24302 21088 24308 21100
rect 24360 21088 24366 21140
rect 25593 21131 25651 21137
rect 25593 21097 25605 21131
rect 25639 21128 25651 21131
rect 26142 21128 26148 21140
rect 25639 21100 26148 21128
rect 25639 21097 25651 21100
rect 25593 21091 25651 21097
rect 23474 21020 23480 21072
rect 23532 21060 23538 21072
rect 25608 21060 25636 21091
rect 26142 21088 26148 21100
rect 26200 21088 26206 21140
rect 26234 21088 26240 21140
rect 26292 21128 26298 21140
rect 26329 21131 26387 21137
rect 26329 21128 26341 21131
rect 26292 21100 26341 21128
rect 26292 21088 26298 21100
rect 26329 21097 26341 21100
rect 26375 21097 26387 21131
rect 26329 21091 26387 21097
rect 27249 21131 27307 21137
rect 27249 21097 27261 21131
rect 27295 21128 27307 21131
rect 27522 21128 27528 21140
rect 27295 21100 27528 21128
rect 27295 21097 27307 21100
rect 27249 21091 27307 21097
rect 27522 21088 27528 21100
rect 27580 21088 27586 21140
rect 29914 21088 29920 21140
rect 29972 21128 29978 21140
rect 30009 21131 30067 21137
rect 30009 21128 30021 21131
rect 29972 21100 30021 21128
rect 29972 21088 29978 21100
rect 30009 21097 30021 21100
rect 30055 21097 30067 21131
rect 30009 21091 30067 21097
rect 35253 21131 35311 21137
rect 35253 21097 35265 21131
rect 35299 21128 35311 21131
rect 35526 21128 35532 21140
rect 35299 21100 35532 21128
rect 35299 21097 35311 21100
rect 35253 21091 35311 21097
rect 35526 21088 35532 21100
rect 35584 21088 35590 21140
rect 35618 21088 35624 21140
rect 35676 21128 35682 21140
rect 36541 21131 36599 21137
rect 36541 21128 36553 21131
rect 35676 21100 36553 21128
rect 35676 21088 35682 21100
rect 36541 21097 36553 21100
rect 36587 21097 36599 21131
rect 36906 21128 36912 21140
rect 36867 21100 36912 21128
rect 36541 21091 36599 21097
rect 36906 21088 36912 21100
rect 36964 21088 36970 21140
rect 23532 21032 25636 21060
rect 28813 21063 28871 21069
rect 23532 21020 23538 21032
rect 28813 21029 28825 21063
rect 28859 21060 28871 21063
rect 30466 21060 30472 21072
rect 28859 21032 30472 21060
rect 28859 21029 28871 21032
rect 28813 21023 28871 21029
rect 30466 21020 30472 21032
rect 30524 21020 30530 21072
rect 47026 21060 47032 21072
rect 46492 21032 47032 21060
rect 32674 20992 32680 21004
rect 23400 20964 32680 20992
rect 14737 20927 14795 20933
rect 14737 20924 14749 20927
rect 14660 20896 14749 20924
rect 14737 20893 14749 20896
rect 14783 20893 14795 20927
rect 14737 20887 14795 20893
rect 14921 20927 14979 20933
rect 14921 20893 14933 20927
rect 14967 20893 14979 20927
rect 14921 20887 14979 20893
rect 16117 20927 16175 20933
rect 16117 20893 16129 20927
rect 16163 20893 16175 20927
rect 16117 20887 16175 20893
rect 16301 20927 16359 20933
rect 16301 20893 16313 20927
rect 16347 20924 16359 20927
rect 16390 20924 16396 20936
rect 16347 20896 16396 20924
rect 16347 20893 16359 20896
rect 16301 20887 16359 20893
rect 16132 20856 16160 20887
rect 16390 20884 16396 20896
rect 16448 20884 16454 20936
rect 16758 20924 16764 20936
rect 16719 20896 16764 20924
rect 16758 20884 16764 20896
rect 16816 20884 16822 20936
rect 16853 20927 16911 20933
rect 16853 20893 16865 20927
rect 16899 20924 16911 20927
rect 16942 20924 16948 20936
rect 16899 20896 16948 20924
rect 16899 20893 16911 20896
rect 16853 20887 16911 20893
rect 16942 20884 16948 20896
rect 17000 20884 17006 20936
rect 17037 20927 17095 20933
rect 17037 20893 17049 20927
rect 17083 20893 17095 20927
rect 17037 20887 17095 20893
rect 17129 20927 17187 20933
rect 17129 20893 17141 20927
rect 17175 20924 17187 20927
rect 17586 20924 17592 20936
rect 17175 20896 17592 20924
rect 17175 20893 17187 20896
rect 17129 20887 17187 20893
rect 16574 20856 16580 20868
rect 16132 20828 16580 20856
rect 16574 20816 16580 20828
rect 16632 20816 16638 20868
rect 17052 20856 17080 20887
rect 17586 20884 17592 20896
rect 17644 20884 17650 20936
rect 19426 20884 19432 20936
rect 19484 20924 19490 20936
rect 19797 20927 19855 20933
rect 19797 20924 19809 20927
rect 19484 20896 19809 20924
rect 19484 20884 19490 20896
rect 19797 20893 19809 20896
rect 19843 20893 19855 20927
rect 19797 20887 19855 20893
rect 20073 20927 20131 20933
rect 20073 20893 20085 20927
rect 20119 20924 20131 20927
rect 20438 20924 20444 20936
rect 20119 20896 20444 20924
rect 20119 20893 20131 20896
rect 20073 20887 20131 20893
rect 20438 20884 20444 20896
rect 20496 20924 20502 20936
rect 22066 20924 22094 20964
rect 32674 20952 32680 20964
rect 32732 20952 32738 21004
rect 42702 20952 42708 21004
rect 42760 20992 42766 21004
rect 46492 21001 46520 21032
rect 47026 21020 47032 21032
rect 47084 21020 47090 21072
rect 43257 20995 43315 21001
rect 43257 20992 43269 20995
rect 42760 20964 43269 20992
rect 42760 20952 42766 20964
rect 43257 20961 43269 20964
rect 43303 20961 43315 20995
rect 43257 20955 43315 20961
rect 46477 20995 46535 21001
rect 46477 20961 46489 20995
rect 46523 20961 46535 20995
rect 46658 20992 46664 21004
rect 46619 20964 46664 20992
rect 46477 20955 46535 20961
rect 46658 20952 46664 20964
rect 46716 20952 46722 21004
rect 48222 20992 48228 21004
rect 48183 20964 48228 20992
rect 48222 20952 48228 20964
rect 48280 20952 48286 21004
rect 20496 20896 22094 20924
rect 20496 20884 20502 20896
rect 22370 20884 22376 20936
rect 22428 20924 22434 20936
rect 22925 20927 22983 20933
rect 22925 20924 22937 20927
rect 22428 20896 22937 20924
rect 22428 20884 22434 20896
rect 22925 20893 22937 20896
rect 22971 20893 22983 20927
rect 22925 20887 22983 20893
rect 23109 20927 23167 20933
rect 23109 20893 23121 20927
rect 23155 20924 23167 20927
rect 23290 20924 23296 20936
rect 23155 20896 23296 20924
rect 23155 20893 23167 20896
rect 23109 20887 23167 20893
rect 17770 20856 17776 20868
rect 17052 20828 17776 20856
rect 17770 20816 17776 20828
rect 17828 20856 17834 20868
rect 18138 20856 18144 20868
rect 17828 20828 18144 20856
rect 17828 20816 17834 20828
rect 18138 20816 18144 20828
rect 18196 20816 18202 20868
rect 22002 20816 22008 20868
rect 22060 20856 22066 20868
rect 23124 20856 23152 20887
rect 23290 20884 23296 20896
rect 23348 20884 23354 20936
rect 23385 20927 23443 20933
rect 23385 20893 23397 20927
rect 23431 20924 23443 20927
rect 25222 20924 25228 20936
rect 23431 20896 25228 20924
rect 23431 20893 23443 20896
rect 23385 20887 23443 20893
rect 22060 20828 23152 20856
rect 22060 20816 22066 20828
rect 16301 20791 16359 20797
rect 16301 20757 16313 20791
rect 16347 20788 16359 20791
rect 17402 20788 17408 20800
rect 16347 20760 17408 20788
rect 16347 20757 16359 20760
rect 16301 20751 16359 20757
rect 17402 20748 17408 20760
rect 17460 20748 17466 20800
rect 17494 20748 17500 20800
rect 17552 20788 17558 20800
rect 18046 20788 18052 20800
rect 17552 20760 18052 20788
rect 17552 20748 17558 20760
rect 18046 20748 18052 20760
rect 18104 20748 18110 20800
rect 19334 20748 19340 20800
rect 19392 20788 19398 20800
rect 19613 20791 19671 20797
rect 19613 20788 19625 20791
rect 19392 20760 19625 20788
rect 19392 20748 19398 20760
rect 19613 20757 19625 20760
rect 19659 20757 19671 20791
rect 19613 20751 19671 20757
rect 19978 20748 19984 20800
rect 20036 20788 20042 20800
rect 22922 20788 22928 20800
rect 20036 20760 22928 20788
rect 20036 20748 20042 20760
rect 22922 20748 22928 20760
rect 22980 20788 22986 20800
rect 23400 20788 23428 20887
rect 25222 20884 25228 20896
rect 25280 20884 25286 20936
rect 26237 20927 26295 20933
rect 26237 20893 26249 20927
rect 26283 20924 26295 20927
rect 26326 20924 26332 20936
rect 26283 20896 26332 20924
rect 26283 20893 26295 20896
rect 26237 20887 26295 20893
rect 26326 20884 26332 20896
rect 26384 20884 26390 20936
rect 27062 20924 27068 20936
rect 27023 20896 27068 20924
rect 27062 20884 27068 20896
rect 27120 20884 27126 20936
rect 27249 20927 27307 20933
rect 27249 20893 27261 20927
rect 27295 20924 27307 20927
rect 27338 20924 27344 20936
rect 27295 20896 27344 20924
rect 27295 20893 27307 20896
rect 27249 20887 27307 20893
rect 27338 20884 27344 20896
rect 27396 20884 27402 20936
rect 27893 20927 27951 20933
rect 27893 20924 27905 20927
rect 27448 20896 27905 20924
rect 25317 20859 25375 20865
rect 25317 20825 25329 20859
rect 25363 20825 25375 20859
rect 25317 20819 25375 20825
rect 22980 20760 23428 20788
rect 25332 20788 25360 20819
rect 26694 20788 26700 20800
rect 25332 20760 26700 20788
rect 22980 20748 22986 20760
rect 26694 20748 26700 20760
rect 26752 20788 26758 20800
rect 27246 20788 27252 20800
rect 26752 20760 27252 20788
rect 26752 20748 26758 20760
rect 27246 20748 27252 20760
rect 27304 20748 27310 20800
rect 27448 20797 27476 20896
rect 27893 20893 27905 20896
rect 27939 20893 27951 20927
rect 27893 20887 27951 20893
rect 28074 20884 28080 20936
rect 28132 20924 28138 20936
rect 28629 20927 28687 20933
rect 28629 20924 28641 20927
rect 28132 20896 28641 20924
rect 28132 20884 28138 20896
rect 28629 20893 28641 20896
rect 28675 20893 28687 20927
rect 28629 20887 28687 20893
rect 29914 20884 29920 20936
rect 29972 20924 29978 20936
rect 30190 20924 30196 20936
rect 29972 20896 30196 20924
rect 29972 20884 29978 20896
rect 30190 20884 30196 20896
rect 30248 20884 30254 20936
rect 30374 20884 30380 20936
rect 30432 20924 30438 20936
rect 30469 20927 30527 20933
rect 30469 20924 30481 20927
rect 30432 20896 30481 20924
rect 30432 20884 30438 20896
rect 30469 20893 30481 20896
rect 30515 20893 30527 20927
rect 30650 20924 30656 20936
rect 30611 20896 30656 20924
rect 30469 20887 30527 20893
rect 30650 20884 30656 20896
rect 30708 20884 30714 20936
rect 35342 20924 35348 20936
rect 35303 20896 35348 20924
rect 35342 20884 35348 20896
rect 35400 20884 35406 20936
rect 36538 20924 36544 20936
rect 36499 20896 36544 20924
rect 36538 20884 36544 20896
rect 36596 20884 36602 20936
rect 36725 20927 36783 20933
rect 36725 20893 36737 20927
rect 36771 20924 36783 20927
rect 37366 20924 37372 20936
rect 36771 20896 37372 20924
rect 36771 20893 36783 20896
rect 36725 20887 36783 20893
rect 37366 20884 37372 20896
rect 37424 20884 37430 20936
rect 43524 20859 43582 20865
rect 43524 20825 43536 20859
rect 43570 20856 43582 20859
rect 43714 20856 43720 20868
rect 43570 20828 43720 20856
rect 43570 20825 43582 20828
rect 43524 20819 43582 20825
rect 43714 20816 43720 20828
rect 43772 20816 43778 20868
rect 27433 20791 27491 20797
rect 27433 20757 27445 20791
rect 27479 20757 27491 20791
rect 27433 20751 27491 20757
rect 27614 20748 27620 20800
rect 27672 20788 27678 20800
rect 28077 20791 28135 20797
rect 28077 20788 28089 20791
rect 27672 20760 28089 20788
rect 27672 20748 27678 20760
rect 28077 20757 28089 20760
rect 28123 20788 28135 20791
rect 28626 20788 28632 20800
rect 28123 20760 28632 20788
rect 28123 20757 28135 20760
rect 28077 20751 28135 20757
rect 28626 20748 28632 20760
rect 28684 20748 28690 20800
rect 34882 20788 34888 20800
rect 34843 20760 34888 20788
rect 34882 20748 34888 20760
rect 34940 20748 34946 20800
rect 44450 20748 44456 20800
rect 44508 20788 44514 20800
rect 44637 20791 44695 20797
rect 44637 20788 44649 20791
rect 44508 20760 44649 20788
rect 44508 20748 44514 20760
rect 44637 20757 44649 20760
rect 44683 20757 44695 20791
rect 44637 20751 44695 20757
rect 47302 20748 47308 20800
rect 47360 20788 47366 20800
rect 47762 20788 47768 20800
rect 47360 20760 47768 20788
rect 47360 20748 47366 20760
rect 47762 20748 47768 20760
rect 47820 20748 47826 20800
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 14642 20584 14648 20596
rect 12728 20556 14648 20584
rect 12728 20460 12756 20556
rect 14642 20544 14648 20556
rect 14700 20544 14706 20596
rect 16298 20544 16304 20596
rect 16356 20584 16362 20596
rect 21174 20584 21180 20596
rect 16356 20556 21180 20584
rect 16356 20544 16362 20556
rect 21174 20544 21180 20556
rect 21232 20544 21238 20596
rect 29733 20587 29791 20593
rect 29733 20553 29745 20587
rect 29779 20584 29791 20587
rect 30098 20584 30104 20596
rect 29779 20556 30104 20584
rect 29779 20553 29791 20556
rect 29733 20547 29791 20553
rect 30098 20544 30104 20556
rect 30156 20544 30162 20596
rect 33873 20587 33931 20593
rect 33873 20553 33885 20587
rect 33919 20584 33931 20587
rect 33919 20556 34836 20584
rect 33919 20553 33931 20556
rect 33873 20547 33931 20553
rect 34808 20528 34836 20556
rect 40586 20544 40592 20596
rect 40644 20584 40650 20596
rect 43714 20584 43720 20596
rect 40644 20556 43576 20584
rect 43675 20556 43720 20584
rect 40644 20544 40650 20556
rect 15197 20519 15255 20525
rect 15197 20485 15209 20519
rect 15243 20516 15255 20519
rect 16942 20516 16948 20528
rect 15243 20488 16948 20516
rect 15243 20485 15255 20488
rect 15197 20479 15255 20485
rect 16942 20476 16948 20488
rect 17000 20476 17006 20528
rect 17494 20516 17500 20528
rect 17329 20488 17500 20516
rect 2038 20448 2044 20460
rect 1999 20420 2044 20448
rect 2038 20408 2044 20420
rect 2096 20408 2102 20460
rect 12526 20448 12532 20460
rect 12487 20420 12532 20448
rect 12526 20408 12532 20420
rect 12584 20408 12590 20460
rect 12710 20408 12716 20460
rect 12768 20448 12774 20460
rect 14093 20451 14151 20457
rect 12768 20420 12861 20448
rect 12768 20408 12774 20420
rect 14093 20417 14105 20451
rect 14139 20448 14151 20451
rect 14642 20448 14648 20460
rect 14139 20420 14648 20448
rect 14139 20417 14151 20420
rect 14093 20411 14151 20417
rect 14642 20408 14648 20420
rect 14700 20408 14706 20460
rect 15102 20448 15108 20460
rect 15063 20420 15108 20448
rect 15102 20408 15108 20420
rect 15160 20408 15166 20460
rect 15286 20448 15292 20460
rect 15247 20420 15292 20448
rect 15286 20408 15292 20420
rect 15344 20408 15350 20460
rect 15933 20451 15991 20457
rect 15933 20417 15945 20451
rect 15979 20417 15991 20451
rect 15933 20411 15991 20417
rect 16025 20451 16083 20457
rect 16025 20417 16037 20451
rect 16071 20417 16083 20451
rect 16025 20411 16083 20417
rect 16301 20451 16359 20457
rect 16301 20417 16313 20451
rect 16347 20448 16359 20451
rect 16666 20448 16672 20460
rect 16347 20420 16672 20448
rect 16347 20417 16359 20420
rect 16301 20411 16359 20417
rect 2225 20383 2283 20389
rect 2225 20349 2237 20383
rect 2271 20380 2283 20383
rect 2406 20380 2412 20392
rect 2271 20352 2412 20380
rect 2271 20349 2283 20352
rect 2225 20343 2283 20349
rect 2406 20340 2412 20352
rect 2464 20340 2470 20392
rect 2774 20340 2780 20392
rect 2832 20380 2838 20392
rect 12802 20380 12808 20392
rect 2832 20352 2877 20380
rect 12763 20352 12808 20380
rect 2832 20340 2838 20352
rect 12802 20340 12808 20352
rect 12860 20340 12866 20392
rect 15948 20312 15976 20411
rect 16040 20380 16068 20411
rect 16666 20408 16672 20420
rect 16724 20408 16730 20460
rect 17034 20448 17040 20460
rect 16995 20420 17040 20448
rect 17034 20408 17040 20420
rect 17092 20408 17098 20460
rect 17329 20457 17357 20488
rect 17494 20476 17500 20488
rect 17552 20476 17558 20528
rect 17678 20476 17684 20528
rect 17736 20516 17742 20528
rect 17865 20519 17923 20525
rect 17865 20516 17877 20519
rect 17736 20488 17877 20516
rect 17736 20476 17742 20488
rect 17865 20485 17877 20488
rect 17911 20485 17923 20519
rect 20714 20516 20720 20528
rect 17865 20479 17923 20485
rect 19260 20488 20720 20516
rect 17221 20451 17279 20457
rect 17221 20417 17233 20451
rect 17267 20417 17279 20451
rect 17221 20411 17279 20417
rect 17313 20451 17371 20457
rect 17313 20417 17325 20451
rect 17359 20417 17371 20451
rect 17313 20411 17371 20417
rect 16853 20383 16911 20389
rect 16853 20380 16865 20383
rect 16040 20352 16865 20380
rect 16853 20349 16865 20352
rect 16899 20349 16911 20383
rect 17126 20380 17132 20392
rect 17088 20352 17132 20380
rect 16853 20343 16911 20349
rect 17126 20340 17132 20352
rect 17184 20340 17190 20392
rect 17236 20324 17264 20411
rect 17402 20408 17408 20460
rect 17460 20448 17466 20460
rect 18049 20451 18107 20457
rect 18049 20448 18061 20451
rect 17460 20438 17908 20448
rect 17972 20438 18061 20448
rect 17460 20420 18061 20438
rect 17460 20408 17466 20420
rect 17880 20410 18000 20420
rect 18049 20417 18061 20420
rect 18095 20417 18107 20451
rect 18049 20411 18107 20417
rect 18138 20408 18144 20460
rect 18196 20448 18202 20460
rect 19260 20457 19288 20488
rect 20714 20476 20720 20488
rect 20772 20476 20778 20528
rect 34577 20519 34635 20525
rect 34577 20516 34589 20519
rect 33704 20488 34589 20516
rect 33704 20460 33732 20488
rect 34577 20485 34589 20488
rect 34623 20485 34635 20519
rect 34790 20516 34796 20528
rect 34751 20488 34796 20516
rect 34577 20479 34635 20485
rect 34790 20476 34796 20488
rect 34848 20476 34854 20528
rect 35342 20476 35348 20528
rect 35400 20516 35406 20528
rect 41506 20516 41512 20528
rect 35400 20488 41512 20516
rect 35400 20476 35406 20488
rect 41506 20476 41512 20488
rect 41564 20516 41570 20528
rect 41690 20516 41696 20528
rect 41564 20488 41696 20516
rect 41564 20476 41570 20488
rect 41690 20476 41696 20488
rect 41748 20476 41754 20528
rect 43548 20516 43576 20556
rect 43714 20544 43720 20556
rect 43772 20544 43778 20596
rect 43548 20488 44220 20516
rect 19245 20451 19303 20457
rect 18196 20420 18241 20448
rect 18196 20408 18202 20420
rect 19245 20417 19257 20451
rect 19291 20417 19303 20451
rect 19245 20411 19303 20417
rect 19334 20408 19340 20460
rect 19392 20448 19398 20460
rect 19501 20451 19559 20457
rect 19501 20448 19513 20451
rect 19392 20420 19513 20448
rect 19392 20408 19398 20420
rect 19501 20417 19513 20420
rect 19547 20417 19559 20451
rect 19501 20411 19559 20417
rect 22005 20451 22063 20457
rect 22005 20417 22017 20451
rect 22051 20448 22063 20451
rect 27614 20448 27620 20460
rect 22051 20420 27620 20448
rect 22051 20417 22063 20420
rect 22005 20411 22063 20417
rect 27614 20408 27620 20420
rect 27672 20408 27678 20460
rect 27706 20408 27712 20460
rect 27764 20448 27770 20460
rect 27801 20451 27859 20457
rect 27801 20448 27813 20451
rect 27764 20420 27813 20448
rect 27764 20408 27770 20420
rect 27801 20417 27813 20420
rect 27847 20417 27859 20451
rect 27801 20411 27859 20417
rect 28902 20408 28908 20460
rect 28960 20448 28966 20460
rect 29549 20451 29607 20457
rect 29549 20448 29561 20451
rect 28960 20420 29561 20448
rect 28960 20408 28966 20420
rect 29549 20417 29561 20420
rect 29595 20417 29607 20451
rect 33686 20448 33692 20460
rect 33647 20420 33692 20448
rect 29549 20411 29607 20417
rect 33686 20408 33692 20420
rect 33744 20408 33750 20460
rect 33965 20451 34023 20457
rect 33965 20417 33977 20451
rect 34011 20448 34023 20451
rect 34808 20448 34836 20476
rect 44192 20460 44220 20488
rect 35621 20451 35679 20457
rect 35621 20448 35633 20451
rect 34011 20420 34652 20448
rect 34808 20420 35633 20448
rect 34011 20417 34023 20420
rect 33965 20411 34023 20417
rect 17494 20340 17500 20392
rect 17552 20380 17558 20392
rect 18414 20380 18420 20392
rect 17552 20352 18420 20380
rect 17552 20340 17558 20352
rect 18414 20340 18420 20352
rect 18472 20340 18478 20392
rect 15948 20284 17080 20312
rect 12158 20204 12164 20256
rect 12216 20244 12222 20256
rect 12345 20247 12403 20253
rect 12345 20244 12357 20247
rect 12216 20216 12357 20244
rect 12216 20204 12222 20216
rect 12345 20213 12357 20216
rect 12391 20213 12403 20247
rect 12345 20207 12403 20213
rect 14277 20247 14335 20253
rect 14277 20213 14289 20247
rect 14323 20244 14335 20247
rect 14550 20244 14556 20256
rect 14323 20216 14556 20244
rect 14323 20213 14335 20216
rect 14277 20207 14335 20213
rect 14550 20204 14556 20216
rect 14608 20204 14614 20256
rect 15746 20244 15752 20256
rect 15707 20216 15752 20244
rect 15746 20204 15752 20216
rect 15804 20204 15810 20256
rect 16206 20244 16212 20256
rect 16167 20216 16212 20244
rect 16206 20204 16212 20216
rect 16264 20204 16270 20256
rect 17052 20244 17080 20284
rect 17218 20272 17224 20324
rect 17276 20272 17282 20324
rect 20254 20272 20260 20324
rect 20312 20312 20318 20324
rect 27985 20315 28043 20321
rect 20312 20284 22094 20312
rect 20312 20272 20318 20284
rect 17865 20247 17923 20253
rect 17865 20244 17877 20247
rect 17052 20216 17877 20244
rect 17865 20213 17877 20216
rect 17911 20213 17923 20247
rect 17865 20207 17923 20213
rect 17954 20204 17960 20256
rect 18012 20244 18018 20256
rect 20346 20244 20352 20256
rect 18012 20216 20352 20244
rect 18012 20204 18018 20216
rect 20346 20204 20352 20216
rect 20404 20244 20410 20256
rect 20625 20247 20683 20253
rect 20625 20244 20637 20247
rect 20404 20216 20637 20244
rect 20404 20204 20410 20216
rect 20625 20213 20637 20216
rect 20671 20213 20683 20247
rect 22066 20244 22094 20284
rect 27985 20281 27997 20315
rect 28031 20312 28043 20315
rect 29914 20312 29920 20324
rect 28031 20284 29920 20312
rect 28031 20281 28043 20284
rect 27985 20275 28043 20281
rect 29914 20272 29920 20284
rect 29972 20272 29978 20324
rect 22189 20247 22247 20253
rect 22189 20244 22201 20247
rect 22066 20216 22201 20244
rect 20625 20207 20683 20213
rect 22189 20213 22201 20216
rect 22235 20244 22247 20247
rect 22370 20244 22376 20256
rect 22235 20216 22376 20244
rect 22235 20213 22247 20216
rect 22189 20207 22247 20213
rect 22370 20204 22376 20216
rect 22428 20204 22434 20256
rect 33689 20247 33747 20253
rect 33689 20213 33701 20247
rect 33735 20244 33747 20247
rect 33778 20244 33784 20256
rect 33735 20216 33784 20244
rect 33735 20213 33747 20216
rect 33689 20207 33747 20213
rect 33778 20204 33784 20216
rect 33836 20204 33842 20256
rect 33870 20204 33876 20256
rect 33928 20244 33934 20256
rect 34624 20253 34652 20420
rect 35621 20417 35633 20420
rect 35667 20417 35679 20451
rect 35621 20411 35679 20417
rect 35894 20408 35900 20460
rect 35952 20448 35958 20460
rect 35989 20451 36047 20457
rect 35989 20448 36001 20451
rect 35952 20420 36001 20448
rect 35952 20408 35958 20420
rect 35989 20417 36001 20420
rect 36035 20448 36047 20451
rect 36538 20448 36544 20460
rect 36035 20420 36544 20448
rect 36035 20417 36047 20420
rect 35989 20411 36047 20417
rect 36538 20408 36544 20420
rect 36596 20408 36602 20460
rect 39384 20451 39442 20457
rect 39384 20417 39396 20451
rect 39430 20448 39442 20451
rect 39942 20448 39948 20460
rect 39430 20420 39948 20448
rect 39430 20417 39442 20420
rect 39384 20411 39442 20417
rect 39942 20408 39948 20420
rect 40000 20408 40006 20460
rect 41785 20451 41843 20457
rect 41785 20417 41797 20451
rect 41831 20448 41843 20451
rect 41874 20448 41880 20460
rect 41831 20420 41880 20448
rect 41831 20417 41843 20420
rect 41785 20411 41843 20417
rect 41874 20408 41880 20420
rect 41932 20408 41938 20460
rect 43993 20451 44051 20457
rect 43993 20417 44005 20451
rect 44039 20448 44051 20451
rect 44082 20448 44088 20460
rect 44039 20420 44088 20448
rect 44039 20417 44051 20420
rect 43993 20411 44051 20417
rect 44082 20408 44088 20420
rect 44140 20408 44146 20460
rect 44174 20408 44180 20460
rect 44232 20448 44238 20460
rect 44269 20451 44327 20457
rect 44269 20448 44281 20451
rect 44232 20420 44281 20448
rect 44232 20408 44238 20420
rect 44269 20417 44281 20420
rect 44315 20448 44327 20451
rect 45646 20448 45652 20460
rect 44315 20420 45652 20448
rect 44315 20417 44327 20420
rect 44269 20411 44327 20417
rect 45646 20408 45652 20420
rect 45704 20408 45710 20460
rect 46198 20448 46204 20460
rect 46159 20420 46204 20448
rect 46198 20408 46204 20420
rect 46256 20408 46262 20460
rect 37734 20340 37740 20392
rect 37792 20380 37798 20392
rect 39117 20383 39175 20389
rect 39117 20380 39129 20383
rect 37792 20352 39129 20380
rect 37792 20340 37798 20352
rect 39117 20349 39129 20352
rect 39163 20349 39175 20383
rect 39117 20343 39175 20349
rect 40126 20340 40132 20392
rect 40184 20380 40190 20392
rect 41049 20383 41107 20389
rect 41049 20380 41061 20383
rect 40184 20352 41061 20380
rect 40184 20340 40190 20352
rect 41049 20349 41061 20352
rect 41095 20380 41107 20383
rect 41322 20380 41328 20392
rect 41095 20352 41328 20380
rect 41095 20349 41107 20352
rect 41049 20343 41107 20349
rect 41322 20340 41328 20352
rect 41380 20340 41386 20392
rect 41509 20383 41567 20389
rect 41509 20349 41521 20383
rect 41555 20349 41567 20383
rect 43898 20380 43904 20392
rect 43859 20352 43904 20380
rect 41509 20343 41567 20349
rect 40497 20315 40555 20321
rect 40497 20281 40509 20315
rect 40543 20312 40555 20315
rect 40770 20312 40776 20324
rect 40543 20284 40776 20312
rect 40543 20281 40555 20284
rect 40497 20275 40555 20281
rect 40770 20272 40776 20284
rect 40828 20312 40834 20324
rect 41524 20312 41552 20343
rect 43898 20340 43904 20352
rect 43956 20340 43962 20392
rect 44361 20383 44419 20389
rect 44361 20349 44373 20383
rect 44407 20380 44419 20383
rect 44450 20380 44456 20392
rect 44407 20352 44456 20380
rect 44407 20349 44419 20352
rect 44361 20343 44419 20349
rect 44450 20340 44456 20352
rect 44508 20340 44514 20392
rect 40828 20284 41552 20312
rect 40828 20272 40834 20284
rect 34425 20247 34483 20253
rect 34425 20244 34437 20247
rect 33928 20216 34437 20244
rect 33928 20204 33934 20216
rect 34425 20213 34437 20216
rect 34471 20213 34483 20247
rect 34425 20207 34483 20213
rect 34609 20247 34667 20253
rect 34609 20213 34621 20247
rect 34655 20244 34667 20247
rect 34882 20244 34888 20256
rect 34655 20216 34888 20244
rect 34655 20213 34667 20216
rect 34609 20207 34667 20213
rect 34882 20204 34888 20216
rect 34940 20204 34946 20256
rect 35986 20244 35992 20256
rect 35947 20216 35992 20244
rect 35986 20204 35992 20216
rect 36044 20204 36050 20256
rect 36170 20244 36176 20256
rect 36131 20216 36176 20244
rect 36170 20204 36176 20216
rect 36228 20204 36234 20256
rect 46290 20244 46296 20256
rect 46251 20216 46296 20244
rect 46290 20204 46296 20216
rect 46348 20204 46354 20256
rect 46474 20204 46480 20256
rect 46532 20244 46538 20256
rect 46845 20247 46903 20253
rect 46845 20244 46857 20247
rect 46532 20216 46857 20244
rect 46532 20204 46538 20216
rect 46845 20213 46857 20216
rect 46891 20213 46903 20247
rect 46845 20207 46903 20213
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 2406 20040 2412 20052
rect 2367 20012 2412 20040
rect 2406 20000 2412 20012
rect 2464 20000 2470 20052
rect 12802 20000 12808 20052
rect 12860 20040 12866 20052
rect 12860 20012 15240 20040
rect 12860 20000 12866 20012
rect 15212 19972 15240 20012
rect 15286 20000 15292 20052
rect 15344 20040 15350 20052
rect 15657 20043 15715 20049
rect 15657 20040 15669 20043
rect 15344 20012 15669 20040
rect 15344 20000 15350 20012
rect 15657 20009 15669 20012
rect 15703 20009 15715 20043
rect 15657 20003 15715 20009
rect 17126 20000 17132 20052
rect 17184 20040 17190 20052
rect 17678 20040 17684 20052
rect 17184 20012 17684 20040
rect 17184 20000 17190 20012
rect 17678 20000 17684 20012
rect 17736 20040 17742 20052
rect 17865 20043 17923 20049
rect 17865 20040 17877 20043
rect 17736 20012 17877 20040
rect 17736 20000 17742 20012
rect 17865 20009 17877 20012
rect 17911 20009 17923 20043
rect 17865 20003 17923 20009
rect 19426 20000 19432 20052
rect 19484 20040 19490 20052
rect 19705 20043 19763 20049
rect 19705 20040 19717 20043
rect 19484 20012 19717 20040
rect 19484 20000 19490 20012
rect 19705 20009 19717 20012
rect 19751 20009 19763 20043
rect 19705 20003 19763 20009
rect 28902 20000 28908 20052
rect 28960 20040 28966 20052
rect 29089 20043 29147 20049
rect 29089 20040 29101 20043
rect 28960 20012 29101 20040
rect 28960 20000 28966 20012
rect 29089 20009 29101 20012
rect 29135 20009 29147 20043
rect 29089 20003 29147 20009
rect 33134 20000 33140 20052
rect 33192 20040 33198 20052
rect 35342 20040 35348 20052
rect 33192 20012 35348 20040
rect 33192 20000 33198 20012
rect 20438 19972 20444 19984
rect 15212 19944 20444 19972
rect 20438 19932 20444 19944
rect 20496 19932 20502 19984
rect 33612 19916 33640 20012
rect 35342 20000 35348 20012
rect 35400 20000 35406 20052
rect 35437 20043 35495 20049
rect 35437 20009 35449 20043
rect 35483 20040 35495 20043
rect 35894 20040 35900 20052
rect 35483 20012 35900 20040
rect 35483 20009 35495 20012
rect 35437 20003 35495 20009
rect 35894 20000 35900 20012
rect 35952 20000 35958 20052
rect 44082 20040 44088 20052
rect 39408 20012 41414 20040
rect 44043 20012 44088 20040
rect 33778 19972 33784 19984
rect 33739 19944 33784 19972
rect 33778 19932 33784 19944
rect 33836 19932 33842 19984
rect 16942 19864 16948 19916
rect 17000 19904 17006 19916
rect 26326 19904 26332 19916
rect 17000 19876 17908 19904
rect 17000 19864 17006 19876
rect 2498 19836 2504 19848
rect 2459 19808 2504 19836
rect 2498 19796 2504 19808
rect 2556 19836 2562 19848
rect 3142 19836 3148 19848
rect 2556 19808 3148 19836
rect 2556 19796 2562 19808
rect 3142 19796 3148 19808
rect 3200 19796 3206 19848
rect 11885 19839 11943 19845
rect 11885 19805 11897 19839
rect 11931 19836 11943 19839
rect 14277 19839 14335 19845
rect 14277 19836 14289 19839
rect 11931 19808 14289 19836
rect 11931 19805 11943 19808
rect 11885 19799 11943 19805
rect 12268 19780 12296 19808
rect 14277 19805 14289 19808
rect 14323 19836 14335 19839
rect 16298 19836 16304 19848
rect 14323 19808 15332 19836
rect 16259 19808 16304 19836
rect 14323 19805 14335 19808
rect 14277 19799 14335 19805
rect 12158 19777 12164 19780
rect 12152 19768 12164 19777
rect 12119 19740 12164 19768
rect 12152 19731 12164 19740
rect 12158 19728 12164 19731
rect 12216 19728 12222 19780
rect 12250 19728 12256 19780
rect 12308 19728 12314 19780
rect 14550 19777 14556 19780
rect 14544 19768 14556 19777
rect 14511 19740 14556 19768
rect 14544 19731 14556 19740
rect 14550 19728 14556 19731
rect 14608 19728 14614 19780
rect 15304 19768 15332 19808
rect 16298 19796 16304 19808
rect 16356 19796 16362 19848
rect 17678 19836 17684 19848
rect 17639 19808 17684 19836
rect 17678 19796 17684 19808
rect 17736 19796 17742 19848
rect 17880 19845 17908 19876
rect 25884 19876 26332 19904
rect 17865 19839 17923 19845
rect 17865 19805 17877 19839
rect 17911 19805 17923 19839
rect 17865 19799 17923 19805
rect 19889 19839 19947 19845
rect 19889 19805 19901 19839
rect 19935 19836 19947 19839
rect 19978 19836 19984 19848
rect 19935 19808 19984 19836
rect 19935 19805 19947 19808
rect 19889 19799 19947 19805
rect 19978 19796 19984 19808
rect 20036 19796 20042 19848
rect 20165 19839 20223 19845
rect 20165 19805 20177 19839
rect 20211 19805 20223 19839
rect 20346 19836 20352 19848
rect 20307 19808 20352 19836
rect 20165 19799 20223 19805
rect 17129 19771 17187 19777
rect 17129 19768 17141 19771
rect 15304 19740 17141 19768
rect 17129 19737 17141 19740
rect 17175 19768 17187 19771
rect 17494 19768 17500 19780
rect 17175 19740 17500 19768
rect 17175 19737 17187 19740
rect 17129 19731 17187 19737
rect 17494 19728 17500 19740
rect 17552 19728 17558 19780
rect 20180 19768 20208 19799
rect 20346 19796 20352 19808
rect 20404 19796 20410 19848
rect 21450 19796 21456 19848
rect 21508 19836 21514 19848
rect 21821 19839 21879 19845
rect 21821 19836 21833 19839
rect 21508 19808 21833 19836
rect 21508 19796 21514 19808
rect 21821 19805 21833 19808
rect 21867 19805 21879 19839
rect 22002 19836 22008 19848
rect 21915 19808 22008 19836
rect 21821 19799 21879 19805
rect 22002 19796 22008 19808
rect 22060 19796 22066 19848
rect 22094 19796 22100 19848
rect 22152 19836 22158 19848
rect 22281 19839 22339 19845
rect 22281 19836 22293 19839
rect 22152 19808 22293 19836
rect 22152 19796 22158 19808
rect 22281 19805 22293 19808
rect 22327 19805 22339 19839
rect 22281 19799 22339 19805
rect 25222 19796 25228 19848
rect 25280 19836 25286 19848
rect 25884 19845 25912 19876
rect 26326 19864 26332 19876
rect 26384 19864 26390 19916
rect 29733 19907 29791 19913
rect 29733 19904 29745 19907
rect 28920 19876 29745 19904
rect 28920 19845 28948 19876
rect 29733 19873 29745 19876
rect 29779 19873 29791 19907
rect 31662 19904 31668 19916
rect 31623 19876 31668 19904
rect 29733 19867 29791 19873
rect 31662 19864 31668 19876
rect 31720 19864 31726 19916
rect 33594 19904 33600 19916
rect 33507 19876 33600 19904
rect 33594 19864 33600 19876
rect 33652 19864 33658 19916
rect 33686 19864 33692 19916
rect 33744 19904 33750 19916
rect 33744 19876 35572 19904
rect 33744 19864 33750 19876
rect 25685 19839 25743 19845
rect 25685 19836 25697 19839
rect 25280 19808 25697 19836
rect 25280 19796 25286 19808
rect 25685 19805 25697 19808
rect 25731 19805 25743 19839
rect 25685 19799 25743 19805
rect 25869 19839 25927 19845
rect 25869 19805 25881 19839
rect 25915 19805 25927 19839
rect 25869 19799 25927 19805
rect 26145 19839 26203 19845
rect 26145 19805 26157 19839
rect 26191 19805 26203 19839
rect 26145 19799 26203 19805
rect 28905 19839 28963 19845
rect 28905 19805 28917 19839
rect 28951 19805 28963 19839
rect 28905 19799 28963 19805
rect 22020 19768 22048 19796
rect 26050 19768 26056 19780
rect 20180 19740 22048 19768
rect 25700 19740 26056 19768
rect 25700 19712 25728 19740
rect 26050 19728 26056 19740
rect 26108 19768 26114 19780
rect 26160 19768 26188 19799
rect 29178 19796 29184 19848
rect 29236 19836 29242 19848
rect 29914 19836 29920 19848
rect 29236 19808 29281 19836
rect 29875 19808 29920 19836
rect 29236 19796 29242 19808
rect 29914 19796 29920 19808
rect 29972 19796 29978 19848
rect 30190 19836 30196 19848
rect 30151 19808 30196 19836
rect 30190 19796 30196 19808
rect 30248 19796 30254 19848
rect 30374 19836 30380 19848
rect 30335 19808 30380 19836
rect 30374 19796 30380 19808
rect 30432 19796 30438 19848
rect 33870 19836 33876 19848
rect 33831 19808 33876 19836
rect 33870 19796 33876 19808
rect 33928 19796 33934 19848
rect 35345 19839 35403 19845
rect 35345 19805 35357 19839
rect 35391 19836 35403 19839
rect 35434 19836 35440 19848
rect 35391 19808 35440 19836
rect 35391 19805 35403 19808
rect 35345 19799 35403 19805
rect 35434 19796 35440 19808
rect 35492 19796 35498 19848
rect 35544 19845 35572 19876
rect 35529 19839 35587 19845
rect 35529 19805 35541 19839
rect 35575 19805 35587 19839
rect 39206 19836 39212 19848
rect 39167 19808 39212 19836
rect 35529 19799 35587 19805
rect 39206 19796 39212 19808
rect 39264 19796 39270 19848
rect 39301 19839 39359 19845
rect 39301 19805 39313 19839
rect 39347 19836 39359 19839
rect 39408 19836 39436 20012
rect 39485 19975 39543 19981
rect 39485 19941 39497 19975
rect 39531 19972 39543 19975
rect 39531 19944 40264 19972
rect 39531 19941 39543 19944
rect 39485 19935 39543 19941
rect 40236 19913 40264 19944
rect 40221 19907 40279 19913
rect 40221 19873 40233 19907
rect 40267 19873 40279 19907
rect 41141 19907 41199 19913
rect 41141 19904 41153 19907
rect 40221 19867 40279 19873
rect 40328 19876 41153 19904
rect 39347 19808 39436 19836
rect 39485 19839 39543 19845
rect 39347 19805 39359 19808
rect 39301 19799 39359 19805
rect 39485 19805 39497 19839
rect 39531 19836 39543 19839
rect 40126 19836 40132 19848
rect 39531 19808 40132 19836
rect 39531 19805 39543 19808
rect 39485 19799 39543 19805
rect 40126 19796 40132 19808
rect 40184 19796 40190 19848
rect 40328 19845 40356 19876
rect 41141 19873 41153 19876
rect 41187 19873 41199 19907
rect 41386 19904 41414 20012
rect 44082 20000 44088 20012
rect 44140 20000 44146 20052
rect 42260 19944 44588 19972
rect 41509 19907 41567 19913
rect 41509 19904 41521 19907
rect 41386 19876 41521 19904
rect 41141 19867 41199 19873
rect 41509 19873 41521 19876
rect 41555 19904 41567 19907
rect 41782 19904 41788 19916
rect 41555 19876 41788 19904
rect 41555 19873 41567 19876
rect 41509 19867 41567 19873
rect 41782 19864 41788 19876
rect 41840 19864 41846 19916
rect 40313 19839 40371 19845
rect 40313 19805 40325 19839
rect 40359 19805 40371 19839
rect 40313 19799 40371 19805
rect 40494 19796 40500 19848
rect 40552 19836 40558 19848
rect 40589 19839 40647 19845
rect 40589 19836 40601 19839
rect 40552 19808 40601 19836
rect 40552 19796 40558 19808
rect 40589 19805 40601 19808
rect 40635 19805 40647 19839
rect 40589 19799 40647 19805
rect 40681 19839 40739 19845
rect 40681 19805 40693 19839
rect 40727 19836 40739 19839
rect 40770 19836 40776 19848
rect 40727 19808 40776 19836
rect 40727 19805 40739 19808
rect 40681 19799 40739 19805
rect 40770 19796 40776 19808
rect 40828 19796 40834 19848
rect 41322 19836 41328 19848
rect 41283 19808 41328 19836
rect 41322 19796 41328 19808
rect 41380 19796 41386 19848
rect 41417 19839 41475 19845
rect 41417 19805 41429 19839
rect 41463 19805 41475 19839
rect 41417 19799 41475 19805
rect 41601 19839 41659 19845
rect 41601 19805 41613 19839
rect 41647 19836 41659 19839
rect 41690 19836 41696 19848
rect 41647 19808 41696 19836
rect 41647 19805 41659 19808
rect 41601 19799 41659 19805
rect 26108 19740 26188 19768
rect 31932 19771 31990 19777
rect 26108 19728 26114 19740
rect 31932 19737 31944 19771
rect 31978 19768 31990 19771
rect 32306 19768 32312 19780
rect 31978 19740 32312 19768
rect 31978 19737 31990 19740
rect 31932 19731 31990 19737
rect 32306 19728 32312 19740
rect 32364 19728 32370 19780
rect 33778 19768 33784 19780
rect 33060 19740 33784 19768
rect 13265 19703 13323 19709
rect 13265 19669 13277 19703
rect 13311 19700 13323 19703
rect 13446 19700 13452 19712
rect 13311 19672 13452 19700
rect 13311 19669 13323 19672
rect 13265 19663 13323 19669
rect 13446 19660 13452 19672
rect 13504 19700 13510 19712
rect 15102 19700 15108 19712
rect 13504 19672 15108 19700
rect 13504 19660 13510 19672
rect 15102 19660 15108 19672
rect 15160 19660 15166 19712
rect 22186 19660 22192 19712
rect 22244 19700 22250 19712
rect 22465 19703 22523 19709
rect 22465 19700 22477 19703
rect 22244 19672 22477 19700
rect 22244 19660 22250 19672
rect 22465 19669 22477 19672
rect 22511 19669 22523 19703
rect 22465 19663 22523 19669
rect 25682 19660 25688 19712
rect 25740 19660 25746 19712
rect 26329 19703 26387 19709
rect 26329 19669 26341 19703
rect 26375 19700 26387 19703
rect 27338 19700 27344 19712
rect 26375 19672 27344 19700
rect 26375 19669 26387 19672
rect 26329 19663 26387 19669
rect 27338 19660 27344 19672
rect 27396 19660 27402 19712
rect 28718 19700 28724 19712
rect 28679 19672 28724 19700
rect 28718 19660 28724 19672
rect 28776 19660 28782 19712
rect 32858 19660 32864 19712
rect 32916 19700 32922 19712
rect 33060 19709 33088 19740
rect 33778 19728 33784 19740
rect 33836 19728 33842 19780
rect 39942 19728 39948 19780
rect 40000 19768 40006 19780
rect 40000 19740 40080 19768
rect 40000 19728 40006 19740
rect 33045 19703 33103 19709
rect 33045 19700 33057 19703
rect 32916 19672 33057 19700
rect 32916 19660 32922 19672
rect 33045 19669 33057 19672
rect 33091 19669 33103 19703
rect 33045 19663 33103 19669
rect 33134 19660 33140 19712
rect 33192 19700 33198 19712
rect 40052 19709 40080 19740
rect 33873 19703 33931 19709
rect 33873 19700 33885 19703
rect 33192 19672 33885 19700
rect 33192 19660 33198 19672
rect 33873 19669 33885 19672
rect 33919 19669 33931 19703
rect 33873 19663 33931 19669
rect 40037 19703 40095 19709
rect 40037 19669 40049 19703
rect 40083 19669 40095 19703
rect 40037 19663 40095 19669
rect 40126 19660 40132 19712
rect 40184 19700 40190 19712
rect 41432 19700 41460 19799
rect 41690 19796 41696 19808
rect 41748 19836 41754 19848
rect 42260 19836 42288 19944
rect 43990 19864 43996 19916
rect 44048 19904 44054 19916
rect 44560 19913 44588 19944
rect 46290 19932 46296 19984
rect 46348 19972 46354 19984
rect 46348 19944 46704 19972
rect 46348 19932 46354 19944
rect 44269 19907 44327 19913
rect 44269 19904 44281 19907
rect 44048 19876 44281 19904
rect 44048 19864 44054 19876
rect 44269 19873 44281 19876
rect 44315 19873 44327 19907
rect 44269 19867 44327 19873
rect 44545 19907 44603 19913
rect 44545 19873 44557 19907
rect 44591 19873 44603 19907
rect 46474 19904 46480 19916
rect 46435 19876 46480 19904
rect 44545 19867 44603 19873
rect 46474 19864 46480 19876
rect 46532 19864 46538 19916
rect 46676 19913 46704 19944
rect 46661 19907 46719 19913
rect 46661 19873 46673 19907
rect 46707 19873 46719 19907
rect 48222 19904 48228 19916
rect 48183 19876 48228 19904
rect 46661 19867 46719 19873
rect 48222 19864 48228 19876
rect 48280 19864 48286 19916
rect 44358 19836 44364 19848
rect 41748 19808 42288 19836
rect 44319 19808 44364 19836
rect 41748 19796 41754 19808
rect 44358 19796 44364 19808
rect 44416 19796 44422 19848
rect 44453 19839 44511 19845
rect 44453 19805 44465 19839
rect 44499 19805 44511 19839
rect 44453 19799 44511 19805
rect 44266 19728 44272 19780
rect 44324 19768 44330 19780
rect 44468 19768 44496 19799
rect 44324 19740 44496 19768
rect 44324 19728 44330 19740
rect 40184 19672 41460 19700
rect 40184 19660 40190 19672
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 12526 19456 12532 19508
rect 12584 19496 12590 19508
rect 12805 19499 12863 19505
rect 12805 19496 12817 19499
rect 12584 19468 12817 19496
rect 12584 19456 12590 19468
rect 12805 19465 12817 19468
rect 12851 19465 12863 19499
rect 14642 19496 14648 19508
rect 14603 19468 14648 19496
rect 12805 19459 12863 19465
rect 14642 19456 14648 19468
rect 14700 19456 14706 19508
rect 15013 19499 15071 19505
rect 15013 19465 15025 19499
rect 15059 19496 15071 19499
rect 15746 19496 15752 19508
rect 15059 19468 15752 19496
rect 15059 19465 15071 19468
rect 15013 19459 15071 19465
rect 15746 19456 15752 19468
rect 15804 19456 15810 19508
rect 16209 19499 16267 19505
rect 16209 19465 16221 19499
rect 16255 19496 16267 19499
rect 17678 19496 17684 19508
rect 16255 19468 17684 19496
rect 16255 19465 16267 19468
rect 16209 19459 16267 19465
rect 17678 19456 17684 19468
rect 17736 19456 17742 19508
rect 25222 19496 25228 19508
rect 25183 19468 25228 19496
rect 25222 19456 25228 19468
rect 25280 19456 25286 19508
rect 27157 19499 27215 19505
rect 27157 19496 27169 19499
rect 26528 19468 27169 19496
rect 13354 19428 13360 19440
rect 13004 19400 13360 19428
rect 13004 19369 13032 19400
rect 13354 19388 13360 19400
rect 13412 19428 13418 19440
rect 14458 19428 14464 19440
rect 13412 19400 14464 19428
rect 13412 19388 13418 19400
rect 14458 19388 14464 19400
rect 14516 19388 14522 19440
rect 15105 19431 15163 19437
rect 15105 19397 15117 19431
rect 15151 19428 15163 19431
rect 15286 19428 15292 19440
rect 15151 19400 15292 19428
rect 15151 19397 15163 19400
rect 15105 19391 15163 19397
rect 15286 19388 15292 19400
rect 15344 19428 15350 19440
rect 15344 19400 16068 19428
rect 15344 19388 15350 19400
rect 12989 19363 13047 19369
rect 12989 19329 13001 19363
rect 13035 19329 13047 19363
rect 12989 19323 13047 19329
rect 13265 19363 13323 19369
rect 13265 19329 13277 19363
rect 13311 19329 13323 19363
rect 13446 19360 13452 19372
rect 13407 19332 13452 19360
rect 13265 19323 13323 19329
rect 13280 19292 13308 19323
rect 13446 19320 13452 19332
rect 13504 19320 13510 19372
rect 16040 19369 16068 19400
rect 16666 19388 16672 19440
rect 16724 19428 16730 19440
rect 16853 19431 16911 19437
rect 16853 19428 16865 19431
rect 16724 19400 16865 19428
rect 16724 19388 16730 19400
rect 16853 19397 16865 19400
rect 16899 19397 16911 19431
rect 17586 19428 17592 19440
rect 16853 19391 16911 19397
rect 17328 19400 17592 19428
rect 16025 19363 16083 19369
rect 15764 19332 15976 19360
rect 13538 19292 13544 19304
rect 13280 19264 13544 19292
rect 13538 19252 13544 19264
rect 13596 19292 13602 19304
rect 13814 19292 13820 19304
rect 13596 19264 13820 19292
rect 13596 19252 13602 19264
rect 13814 19252 13820 19264
rect 13872 19252 13878 19304
rect 14918 19252 14924 19304
rect 14976 19292 14982 19304
rect 15197 19295 15255 19301
rect 15197 19292 15209 19295
rect 14976 19264 15209 19292
rect 14976 19252 14982 19264
rect 15197 19261 15209 19264
rect 15243 19292 15255 19295
rect 15764 19292 15792 19332
rect 15243 19264 15792 19292
rect 15841 19295 15899 19301
rect 15243 19261 15255 19264
rect 15197 19255 15255 19261
rect 15841 19261 15853 19295
rect 15887 19261 15899 19295
rect 15948 19292 15976 19332
rect 16025 19329 16037 19363
rect 16071 19329 16083 19363
rect 16025 19323 16083 19329
rect 16942 19320 16948 19372
rect 17000 19360 17006 19372
rect 17083 19363 17141 19369
rect 17083 19360 17095 19363
rect 17000 19332 17095 19360
rect 17000 19320 17006 19332
rect 17083 19329 17095 19332
rect 17129 19329 17141 19363
rect 17218 19360 17224 19372
rect 17179 19332 17224 19360
rect 17083 19323 17141 19329
rect 17218 19320 17224 19332
rect 17276 19320 17282 19372
rect 17328 19369 17356 19400
rect 17586 19388 17592 19400
rect 17644 19388 17650 19440
rect 20070 19428 20076 19440
rect 19352 19400 20076 19428
rect 17313 19363 17371 19369
rect 17313 19329 17325 19363
rect 17359 19329 17371 19363
rect 17313 19323 17371 19329
rect 17402 19320 17408 19372
rect 17460 19360 17466 19372
rect 19352 19369 19380 19400
rect 20070 19388 20076 19400
rect 20128 19388 20134 19440
rect 20622 19428 20628 19440
rect 20583 19400 20628 19428
rect 20622 19388 20628 19400
rect 20680 19388 20686 19440
rect 21174 19388 21180 19440
rect 21232 19428 21238 19440
rect 21453 19431 21511 19437
rect 21453 19428 21465 19431
rect 21232 19400 21465 19428
rect 21232 19388 21238 19400
rect 21453 19397 21465 19400
rect 21499 19397 21511 19431
rect 21453 19391 21511 19397
rect 26360 19431 26418 19437
rect 26360 19397 26372 19431
rect 26406 19428 26418 19431
rect 26528 19428 26556 19468
rect 27157 19465 27169 19468
rect 27203 19465 27215 19499
rect 27157 19459 27215 19465
rect 29825 19499 29883 19505
rect 29825 19465 29837 19499
rect 29871 19496 29883 19499
rect 30374 19496 30380 19508
rect 29871 19468 30380 19496
rect 29871 19465 29883 19468
rect 29825 19459 29883 19465
rect 30374 19456 30380 19468
rect 30432 19496 30438 19508
rect 32306 19496 32312 19508
rect 30432 19468 31754 19496
rect 32267 19468 32312 19496
rect 30432 19456 30438 19468
rect 28718 19437 28724 19440
rect 28712 19428 28724 19437
rect 26406 19400 26556 19428
rect 26620 19400 28488 19428
rect 28679 19400 28724 19428
rect 26406 19397 26418 19400
rect 26360 19391 26418 19397
rect 17497 19363 17555 19369
rect 17497 19360 17509 19363
rect 17460 19332 17509 19360
rect 17460 19320 17466 19332
rect 17497 19329 17509 19332
rect 17543 19329 17555 19363
rect 17497 19323 17555 19329
rect 19337 19363 19395 19369
rect 19337 19329 19349 19363
rect 19383 19329 19395 19363
rect 19337 19323 19395 19329
rect 19521 19363 19579 19369
rect 19521 19329 19533 19363
rect 19567 19360 19579 19363
rect 19978 19360 19984 19372
rect 19567 19332 19984 19360
rect 19567 19329 19579 19332
rect 19521 19323 19579 19329
rect 19978 19320 19984 19332
rect 20036 19320 20042 19372
rect 22186 19360 22192 19372
rect 20548 19332 20760 19360
rect 22147 19332 22192 19360
rect 16482 19292 16488 19304
rect 15948 19264 16488 19292
rect 15841 19255 15899 19261
rect 15102 19184 15108 19236
rect 15160 19224 15166 19236
rect 15856 19224 15884 19255
rect 16482 19252 16488 19264
rect 16540 19252 16546 19304
rect 19242 19292 19248 19304
rect 19203 19264 19248 19292
rect 19242 19252 19248 19264
rect 19300 19252 19306 19304
rect 20548 19224 20576 19332
rect 20732 19292 20760 19332
rect 22186 19320 22192 19332
rect 22244 19320 22250 19372
rect 22370 19360 22376 19372
rect 22331 19332 22376 19360
rect 22370 19320 22376 19332
rect 22428 19320 22434 19372
rect 23652 19363 23710 19369
rect 23652 19329 23664 19363
rect 23698 19360 23710 19363
rect 25222 19360 25228 19372
rect 23698 19332 25228 19360
rect 23698 19329 23710 19332
rect 23652 19323 23710 19329
rect 25222 19320 25228 19332
rect 25280 19320 25286 19372
rect 26620 19369 26648 19400
rect 26605 19363 26663 19369
rect 26605 19329 26617 19363
rect 26651 19329 26663 19363
rect 27338 19360 27344 19372
rect 27299 19332 27344 19360
rect 26605 19323 26663 19329
rect 27338 19320 27344 19332
rect 27396 19320 27402 19372
rect 27430 19320 27436 19372
rect 27488 19360 27494 19372
rect 28460 19369 28488 19400
rect 28712 19391 28724 19400
rect 28718 19388 28724 19391
rect 28776 19388 28782 19440
rect 31726 19428 31754 19468
rect 32306 19456 32312 19468
rect 32364 19456 32370 19508
rect 32398 19456 32404 19508
rect 32456 19496 32462 19508
rect 33318 19496 33324 19508
rect 32456 19468 33324 19496
rect 32456 19456 32462 19468
rect 33318 19456 33324 19468
rect 33376 19456 33382 19508
rect 34517 19499 34575 19505
rect 34517 19496 34529 19499
rect 33612 19468 34529 19496
rect 32585 19431 32643 19437
rect 32585 19428 32597 19431
rect 31726 19400 32597 19428
rect 32585 19397 32597 19400
rect 32631 19397 32643 19431
rect 32585 19391 32643 19397
rect 32677 19431 32735 19437
rect 32677 19397 32689 19431
rect 32723 19428 32735 19431
rect 33410 19428 33416 19440
rect 32723 19400 33416 19428
rect 32723 19397 32735 19400
rect 32677 19391 32735 19397
rect 33410 19388 33416 19400
rect 33468 19388 33474 19440
rect 27525 19363 27583 19369
rect 27525 19360 27537 19363
rect 27488 19332 27537 19360
rect 27488 19320 27494 19332
rect 27525 19329 27537 19332
rect 27571 19329 27583 19363
rect 27525 19323 27583 19329
rect 28445 19363 28503 19369
rect 28445 19329 28457 19363
rect 28491 19360 28503 19363
rect 28534 19360 28540 19372
rect 28491 19332 28540 19360
rect 28491 19329 28503 19332
rect 28445 19323 28503 19329
rect 28534 19320 28540 19332
rect 28592 19320 28598 19372
rect 30650 19360 30656 19372
rect 30611 19332 30656 19360
rect 30650 19320 30656 19332
rect 30708 19320 30714 19372
rect 30834 19320 30840 19372
rect 30892 19360 30898 19372
rect 31294 19360 31300 19372
rect 30892 19332 31300 19360
rect 30892 19320 30898 19332
rect 31294 19320 31300 19332
rect 31352 19320 31358 19372
rect 31846 19320 31852 19372
rect 31904 19360 31910 19372
rect 32398 19360 32404 19372
rect 31904 19332 32404 19360
rect 31904 19320 31910 19332
rect 32398 19320 32404 19332
rect 32456 19369 32462 19372
rect 32456 19363 32505 19369
rect 32456 19329 32459 19363
rect 32493 19329 32505 19363
rect 32858 19360 32864 19372
rect 32819 19332 32864 19360
rect 32456 19323 32505 19329
rect 32456 19320 32462 19323
rect 32858 19320 32864 19332
rect 32916 19320 32922 19372
rect 32953 19363 33011 19369
rect 32953 19329 32965 19363
rect 32999 19360 33011 19363
rect 33134 19360 33140 19372
rect 32999 19332 33140 19360
rect 32999 19329 33011 19332
rect 32953 19323 33011 19329
rect 33134 19320 33140 19332
rect 33192 19320 33198 19372
rect 33612 19369 33640 19468
rect 34517 19465 34529 19468
rect 34563 19496 34575 19499
rect 34698 19496 34704 19508
rect 34563 19468 34704 19496
rect 34563 19465 34575 19468
rect 34517 19459 34575 19465
rect 34698 19456 34704 19468
rect 34756 19456 34762 19508
rect 39117 19499 39175 19505
rect 39117 19465 39129 19499
rect 39163 19496 39175 19499
rect 40218 19496 40224 19508
rect 39163 19468 40224 19496
rect 39163 19465 39175 19468
rect 39117 19459 39175 19465
rect 40218 19456 40224 19468
rect 40276 19456 40282 19508
rect 43898 19456 43904 19508
rect 43956 19496 43962 19508
rect 44183 19499 44241 19505
rect 44183 19496 44195 19499
rect 43956 19468 44195 19496
rect 43956 19456 43962 19468
rect 44183 19465 44195 19468
rect 44229 19465 44241 19499
rect 44183 19459 44241 19465
rect 33870 19388 33876 19440
rect 33928 19428 33934 19440
rect 39853 19431 39911 19437
rect 33928 19400 34744 19428
rect 33928 19388 33934 19400
rect 33597 19363 33655 19369
rect 33597 19334 33609 19363
rect 33428 19329 33609 19334
rect 33643 19329 33655 19363
rect 33778 19360 33784 19372
rect 33428 19323 33655 19329
rect 33704 19332 33784 19360
rect 33428 19306 33640 19323
rect 22465 19295 22523 19301
rect 22465 19292 22477 19295
rect 20732 19264 22477 19292
rect 22465 19261 22477 19264
rect 22511 19292 22523 19295
rect 23014 19292 23020 19304
rect 22511 19264 23020 19292
rect 22511 19261 22523 19264
rect 22465 19255 22523 19261
rect 23014 19252 23020 19264
rect 23072 19252 23078 19304
rect 23385 19295 23443 19301
rect 23385 19261 23397 19295
rect 23431 19261 23443 19295
rect 23385 19255 23443 19261
rect 27617 19295 27675 19301
rect 27617 19261 27629 19295
rect 27663 19261 27675 19295
rect 27617 19255 27675 19261
rect 30929 19295 30987 19301
rect 30929 19261 30941 19295
rect 30975 19292 30987 19295
rect 31570 19292 31576 19304
rect 30975 19264 31576 19292
rect 30975 19261 30987 19264
rect 30929 19255 30987 19261
rect 15160 19196 15884 19224
rect 15948 19196 20576 19224
rect 15160 19184 15166 19196
rect 12618 19116 12624 19168
rect 12676 19156 12682 19168
rect 15948 19156 15976 19196
rect 20622 19184 20628 19236
rect 20680 19224 20686 19236
rect 22830 19224 22836 19236
rect 20680 19196 22836 19224
rect 20680 19184 20686 19196
rect 22830 19184 22836 19196
rect 22888 19224 22894 19236
rect 23400 19224 23428 19255
rect 22888 19196 23428 19224
rect 22888 19184 22894 19196
rect 19702 19156 19708 19168
rect 12676 19128 15976 19156
rect 19663 19128 19708 19156
rect 12676 19116 12682 19128
rect 19702 19116 19708 19128
rect 19760 19116 19766 19168
rect 22002 19156 22008 19168
rect 21963 19128 22008 19156
rect 22002 19116 22008 19128
rect 22060 19116 22066 19168
rect 24762 19156 24768 19168
rect 24723 19128 24768 19156
rect 24762 19116 24768 19128
rect 24820 19116 24826 19168
rect 27632 19156 27660 19255
rect 31570 19252 31576 19264
rect 31628 19292 31634 19304
rect 33428 19292 33456 19306
rect 33704 19301 33732 19332
rect 33778 19320 33784 19332
rect 33836 19360 33842 19372
rect 34422 19360 34428 19372
rect 33836 19332 34428 19360
rect 33836 19320 33842 19332
rect 34422 19320 34428 19332
rect 34480 19320 34486 19372
rect 34716 19369 34744 19400
rect 39853 19397 39865 19431
rect 39899 19428 39911 19431
rect 40402 19428 40408 19440
rect 39899 19400 40408 19428
rect 39899 19397 39911 19400
rect 39853 19391 39911 19397
rect 40402 19388 40408 19400
rect 40460 19388 40466 19440
rect 43990 19388 43996 19440
rect 44048 19428 44054 19440
rect 44085 19431 44143 19437
rect 44085 19428 44097 19431
rect 44048 19400 44097 19428
rect 44048 19388 44054 19400
rect 44085 19397 44097 19400
rect 44131 19397 44143 19431
rect 44913 19431 44971 19437
rect 44913 19428 44925 19431
rect 44085 19391 44143 19397
rect 44284 19400 44925 19428
rect 34701 19363 34759 19369
rect 34701 19329 34713 19363
rect 34747 19329 34759 19363
rect 34701 19323 34759 19329
rect 38004 19363 38062 19369
rect 38004 19329 38016 19363
rect 38050 19360 38062 19363
rect 39577 19363 39635 19369
rect 39577 19360 39589 19363
rect 38050 19332 39589 19360
rect 38050 19329 38062 19332
rect 38004 19323 38062 19329
rect 39577 19329 39589 19332
rect 39623 19329 39635 19363
rect 39577 19323 39635 19329
rect 39761 19363 39819 19369
rect 39761 19329 39773 19363
rect 39807 19329 39819 19363
rect 39942 19360 39948 19372
rect 39903 19332 39948 19360
rect 39761 19323 39819 19329
rect 31628 19264 33456 19292
rect 33689 19295 33747 19301
rect 31628 19252 31634 19264
rect 33689 19261 33701 19295
rect 33735 19292 33747 19295
rect 37734 19292 37740 19304
rect 33735 19264 33769 19292
rect 37695 19264 37740 19292
rect 33735 19261 33747 19264
rect 33689 19255 33747 19261
rect 37734 19252 37740 19264
rect 37792 19252 37798 19304
rect 39776 19224 39804 19323
rect 39942 19320 39948 19332
rect 40000 19320 40006 19372
rect 40083 19363 40141 19369
rect 40083 19329 40095 19363
rect 40129 19360 40141 19363
rect 40586 19360 40592 19372
rect 40129 19332 40592 19360
rect 40129 19329 40141 19332
rect 40083 19323 40141 19329
rect 40586 19320 40592 19332
rect 40644 19320 40650 19372
rect 40954 19360 40960 19372
rect 40915 19332 40960 19360
rect 40954 19320 40960 19332
rect 41012 19320 41018 19372
rect 41782 19360 41788 19372
rect 41743 19332 41788 19360
rect 41782 19320 41788 19332
rect 41840 19320 41846 19372
rect 43438 19360 43444 19372
rect 43399 19332 43444 19360
rect 43438 19320 43444 19332
rect 43496 19320 43502 19372
rect 43625 19363 43683 19369
rect 43625 19329 43637 19363
rect 43671 19360 43683 19363
rect 44008 19360 44036 19388
rect 44284 19372 44312 19400
rect 44913 19397 44925 19400
rect 44959 19397 44971 19431
rect 44913 19391 44971 19397
rect 44266 19360 44272 19372
rect 43671 19332 44036 19360
rect 44227 19332 44272 19360
rect 43671 19329 43683 19332
rect 43625 19323 43683 19329
rect 44266 19320 44272 19332
rect 44324 19320 44330 19372
rect 44358 19320 44364 19372
rect 44416 19360 44422 19372
rect 44416 19332 44461 19360
rect 44416 19320 44422 19332
rect 44634 19320 44640 19372
rect 44692 19360 44698 19372
rect 44821 19363 44879 19369
rect 44821 19360 44833 19363
rect 44692 19332 44833 19360
rect 44692 19320 44698 19332
rect 44821 19329 44833 19332
rect 44867 19329 44879 19363
rect 44821 19323 44879 19329
rect 45005 19363 45063 19369
rect 45005 19329 45017 19363
rect 45051 19329 45063 19363
rect 47210 19360 47216 19372
rect 47123 19332 47216 19360
rect 45005 19323 45063 19329
rect 40218 19292 40224 19304
rect 40179 19264 40224 19292
rect 40218 19252 40224 19264
rect 40276 19292 40282 19304
rect 40681 19295 40739 19301
rect 40681 19292 40693 19295
rect 40276 19264 40693 19292
rect 40276 19252 40282 19264
rect 40681 19261 40693 19264
rect 40727 19261 40739 19295
rect 40681 19255 40739 19261
rect 40770 19252 40776 19304
rect 40828 19292 40834 19304
rect 41969 19295 42027 19301
rect 41969 19292 41981 19295
rect 40828 19264 41981 19292
rect 40828 19252 40834 19264
rect 41969 19261 41981 19264
rect 42015 19261 42027 19295
rect 41969 19255 42027 19261
rect 44542 19252 44548 19304
rect 44600 19292 44606 19304
rect 45020 19292 45048 19323
rect 47210 19320 47216 19332
rect 47268 19360 47274 19372
rect 47578 19360 47584 19372
rect 47268 19332 47584 19360
rect 47268 19320 47274 19332
rect 47578 19320 47584 19332
rect 47636 19320 47642 19372
rect 44600 19264 45048 19292
rect 44600 19252 44606 19264
rect 39942 19224 39948 19236
rect 39776 19196 39948 19224
rect 39942 19184 39948 19196
rect 40000 19184 40006 19236
rect 29178 19156 29184 19168
rect 27632 19128 29184 19156
rect 29178 19116 29184 19128
rect 29236 19116 29242 19168
rect 30466 19156 30472 19168
rect 30427 19128 30472 19156
rect 30466 19116 30472 19128
rect 30524 19116 30530 19168
rect 33686 19116 33692 19168
rect 33744 19156 33750 19168
rect 33965 19159 34023 19165
rect 33965 19156 33977 19159
rect 33744 19128 33977 19156
rect 33744 19116 33750 19128
rect 33965 19125 33977 19128
rect 34011 19125 34023 19159
rect 33965 19119 34023 19125
rect 34790 19116 34796 19168
rect 34848 19156 34854 19168
rect 34885 19159 34943 19165
rect 34885 19156 34897 19159
rect 34848 19128 34897 19156
rect 34848 19116 34854 19128
rect 34885 19125 34897 19128
rect 34931 19125 34943 19159
rect 34885 19119 34943 19125
rect 40773 19159 40831 19165
rect 40773 19125 40785 19159
rect 40819 19156 40831 19159
rect 40862 19156 40868 19168
rect 40819 19128 40868 19156
rect 40819 19125 40831 19128
rect 40773 19119 40831 19125
rect 40862 19116 40868 19128
rect 40920 19116 40926 19168
rect 41141 19159 41199 19165
rect 41141 19125 41153 19159
rect 41187 19156 41199 19159
rect 41230 19156 41236 19168
rect 41187 19128 41236 19156
rect 41187 19125 41199 19128
rect 41141 19119 41199 19125
rect 41230 19116 41236 19128
rect 41288 19116 41294 19168
rect 41598 19156 41604 19168
rect 41559 19128 41604 19156
rect 41598 19116 41604 19128
rect 41656 19116 41662 19168
rect 43625 19159 43683 19165
rect 43625 19125 43637 19159
rect 43671 19156 43683 19159
rect 44174 19156 44180 19168
rect 43671 19128 44180 19156
rect 43671 19125 43683 19128
rect 43625 19119 43683 19125
rect 44174 19116 44180 19128
rect 44232 19116 44238 19168
rect 47118 19156 47124 19168
rect 47079 19128 47124 19156
rect 47118 19116 47124 19128
rect 47176 19116 47182 19168
rect 47762 19156 47768 19168
rect 47723 19128 47768 19156
rect 47762 19116 47768 19128
rect 47820 19116 47826 19168
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 19242 18912 19248 18964
rect 19300 18952 19306 18964
rect 25038 18952 25044 18964
rect 19300 18924 25044 18952
rect 19300 18912 19306 18924
rect 25038 18912 25044 18924
rect 25096 18912 25102 18964
rect 25222 18952 25228 18964
rect 25183 18924 25228 18952
rect 25222 18912 25228 18924
rect 25280 18912 25286 18964
rect 31570 18952 31576 18964
rect 25332 18924 31156 18952
rect 31531 18924 31576 18952
rect 23014 18844 23020 18896
rect 23072 18884 23078 18896
rect 25332 18884 25360 18924
rect 28626 18884 28632 18896
rect 23072 18856 25360 18884
rect 28587 18856 28632 18884
rect 23072 18844 23078 18856
rect 28626 18844 28632 18856
rect 28684 18844 28690 18896
rect 31128 18884 31156 18924
rect 31570 18912 31576 18924
rect 31628 18912 31634 18964
rect 39206 18912 39212 18964
rect 39264 18952 39270 18964
rect 39393 18955 39451 18961
rect 39393 18952 39405 18955
rect 39264 18924 39405 18952
rect 39264 18912 39270 18924
rect 39393 18921 39405 18924
rect 39439 18952 39451 18955
rect 39942 18952 39948 18964
rect 39439 18924 39948 18952
rect 39439 18921 39451 18924
rect 39393 18915 39451 18921
rect 39942 18912 39948 18924
rect 40000 18912 40006 18964
rect 40770 18952 40776 18964
rect 40731 18924 40776 18952
rect 40770 18912 40776 18924
rect 40828 18912 40834 18964
rect 41233 18955 41291 18961
rect 41233 18921 41245 18955
rect 41279 18921 41291 18955
rect 41233 18915 41291 18921
rect 33502 18884 33508 18896
rect 31128 18856 33508 18884
rect 33502 18844 33508 18856
rect 33560 18844 33566 18896
rect 35529 18887 35587 18893
rect 35529 18853 35541 18887
rect 35575 18853 35587 18887
rect 35529 18847 35587 18853
rect 15102 18776 15108 18828
rect 15160 18816 15166 18828
rect 15160 18788 15700 18816
rect 15160 18776 15166 18788
rect 2038 18748 2044 18760
rect 1999 18720 2044 18748
rect 2038 18708 2044 18720
rect 2096 18708 2102 18760
rect 15286 18708 15292 18760
rect 15344 18748 15350 18760
rect 15672 18757 15700 18788
rect 16758 18776 16764 18828
rect 16816 18816 16822 18828
rect 22830 18816 22836 18828
rect 16816 18788 17356 18816
rect 22791 18788 22836 18816
rect 16816 18776 16822 18788
rect 15473 18751 15531 18757
rect 15473 18748 15485 18751
rect 15344 18720 15485 18748
rect 15344 18708 15350 18720
rect 15473 18717 15485 18720
rect 15519 18717 15531 18751
rect 15473 18711 15531 18717
rect 15657 18751 15715 18757
rect 15657 18717 15669 18751
rect 15703 18717 15715 18751
rect 15657 18711 15715 18717
rect 16942 18708 16948 18760
rect 17000 18748 17006 18760
rect 17328 18757 17356 18788
rect 22830 18776 22836 18788
rect 22888 18776 22894 18828
rect 27801 18819 27859 18825
rect 27801 18785 27813 18819
rect 27847 18816 27859 18819
rect 28534 18816 28540 18828
rect 27847 18788 28540 18816
rect 27847 18785 27859 18788
rect 27801 18779 27859 18785
rect 28534 18776 28540 18788
rect 28592 18816 28598 18828
rect 28592 18788 30236 18816
rect 28592 18776 28598 18788
rect 17037 18751 17095 18757
rect 17037 18748 17049 18751
rect 17000 18720 17049 18748
rect 17000 18708 17006 18720
rect 17037 18717 17049 18720
rect 17083 18717 17095 18751
rect 17037 18711 17095 18717
rect 17313 18751 17371 18757
rect 17313 18717 17325 18751
rect 17359 18717 17371 18751
rect 17313 18711 17371 18717
rect 19334 18708 19340 18760
rect 19392 18748 19398 18760
rect 19702 18757 19708 18760
rect 19429 18751 19487 18757
rect 19429 18748 19441 18751
rect 19392 18720 19441 18748
rect 19392 18708 19398 18720
rect 19429 18717 19441 18720
rect 19475 18717 19487 18751
rect 19696 18748 19708 18757
rect 19663 18720 19708 18748
rect 19429 18711 19487 18717
rect 19696 18711 19708 18720
rect 19702 18708 19708 18711
rect 19760 18708 19766 18760
rect 22002 18708 22008 18760
rect 22060 18748 22066 18760
rect 22566 18751 22624 18757
rect 22566 18748 22578 18751
rect 22060 18720 22578 18748
rect 22060 18708 22066 18720
rect 22566 18717 22578 18720
rect 22612 18717 22624 18751
rect 22566 18711 22624 18717
rect 23934 18708 23940 18760
rect 23992 18748 23998 18760
rect 24581 18751 24639 18757
rect 24581 18748 24593 18751
rect 23992 18720 24593 18748
rect 23992 18708 23998 18720
rect 24581 18717 24593 18720
rect 24627 18717 24639 18751
rect 24581 18711 24639 18717
rect 24674 18751 24732 18757
rect 24674 18717 24686 18751
rect 24720 18748 24732 18751
rect 24762 18748 24768 18760
rect 24720 18720 24768 18748
rect 24720 18717 24732 18720
rect 24674 18711 24732 18717
rect 15565 18683 15623 18689
rect 15565 18649 15577 18683
rect 15611 18680 15623 18683
rect 17221 18683 17279 18689
rect 17221 18680 17233 18683
rect 15611 18652 17233 18680
rect 15611 18649 15623 18652
rect 15565 18643 15623 18649
rect 17221 18649 17233 18652
rect 17267 18680 17279 18683
rect 17402 18680 17408 18692
rect 17267 18652 17408 18680
rect 17267 18649 17279 18652
rect 17221 18643 17279 18649
rect 17402 18640 17408 18652
rect 17460 18640 17466 18692
rect 23845 18683 23903 18689
rect 23845 18649 23857 18683
rect 23891 18649 23903 18683
rect 23845 18643 23903 18649
rect 24029 18683 24087 18689
rect 24029 18649 24041 18683
rect 24075 18680 24087 18683
rect 24688 18680 24716 18711
rect 24762 18708 24768 18720
rect 24820 18708 24826 18760
rect 25087 18751 25145 18757
rect 25087 18717 25099 18751
rect 25133 18748 25145 18751
rect 25222 18748 25228 18760
rect 25133 18720 25228 18748
rect 25133 18717 25145 18720
rect 25087 18711 25145 18717
rect 25222 18708 25228 18720
rect 25280 18748 25286 18760
rect 25590 18748 25596 18760
rect 25280 18720 25596 18748
rect 25280 18708 25286 18720
rect 25590 18708 25596 18720
rect 25648 18708 25654 18760
rect 28442 18748 28448 18760
rect 28403 18720 28448 18748
rect 28442 18708 28448 18720
rect 28500 18708 28506 18760
rect 28721 18751 28779 18757
rect 28721 18717 28733 18751
rect 28767 18748 28779 18751
rect 29178 18748 29184 18760
rect 28767 18720 29184 18748
rect 28767 18717 28779 18720
rect 28721 18711 28779 18717
rect 29178 18708 29184 18720
rect 29236 18748 29242 18760
rect 29822 18748 29828 18760
rect 29236 18720 29828 18748
rect 29236 18708 29242 18720
rect 29822 18708 29828 18720
rect 29880 18708 29886 18760
rect 30208 18757 30236 18788
rect 34790 18776 34796 18828
rect 34848 18816 34854 18828
rect 35069 18819 35127 18825
rect 35069 18816 35081 18819
rect 34848 18788 35081 18816
rect 34848 18776 34854 18788
rect 35069 18785 35081 18788
rect 35115 18785 35127 18819
rect 35069 18779 35127 18785
rect 30193 18751 30251 18757
rect 30193 18717 30205 18751
rect 30239 18748 30251 18751
rect 31662 18748 31668 18760
rect 30239 18720 31668 18748
rect 30239 18717 30251 18720
rect 30193 18711 30251 18717
rect 31662 18708 31668 18720
rect 31720 18748 31726 18760
rect 32769 18751 32827 18757
rect 32769 18748 32781 18751
rect 31720 18720 32781 18748
rect 31720 18708 31726 18720
rect 32769 18717 32781 18720
rect 32815 18717 32827 18751
rect 32769 18711 32827 18717
rect 35161 18751 35219 18757
rect 35161 18717 35173 18751
rect 35207 18748 35219 18751
rect 35434 18748 35440 18760
rect 35207 18720 35440 18748
rect 35207 18717 35219 18720
rect 35161 18711 35219 18717
rect 35434 18708 35440 18720
rect 35492 18708 35498 18760
rect 35544 18748 35572 18847
rect 40310 18844 40316 18896
rect 40368 18884 40374 18896
rect 41248 18884 41276 18915
rect 41782 18912 41788 18964
rect 41840 18952 41846 18964
rect 42153 18955 42211 18961
rect 42153 18952 42165 18955
rect 41840 18924 42165 18952
rect 41840 18912 41846 18924
rect 42153 18921 42165 18924
rect 42199 18921 42211 18955
rect 42153 18915 42211 18921
rect 40368 18856 41276 18884
rect 41601 18887 41659 18893
rect 40368 18844 40374 18856
rect 41601 18853 41613 18887
rect 41647 18884 41659 18887
rect 42886 18884 42892 18896
rect 41647 18856 42892 18884
rect 41647 18853 41659 18856
rect 41601 18847 41659 18853
rect 42886 18844 42892 18856
rect 42944 18844 42950 18896
rect 44542 18844 44548 18896
rect 44600 18884 44606 18896
rect 45462 18884 45468 18896
rect 44600 18856 45468 18884
rect 44600 18844 44606 18856
rect 45462 18844 45468 18856
rect 45520 18884 45526 18896
rect 47762 18884 47768 18896
rect 45520 18856 45876 18884
rect 45520 18844 45526 18856
rect 40218 18776 40224 18828
rect 40276 18816 40282 18828
rect 44266 18816 44272 18828
rect 40276 18788 42104 18816
rect 40276 18776 40282 18788
rect 36357 18751 36415 18757
rect 36357 18748 36369 18751
rect 35544 18720 36369 18748
rect 36357 18717 36369 18720
rect 36403 18717 36415 18751
rect 36357 18711 36415 18717
rect 36446 18708 36452 18760
rect 36504 18748 36510 18760
rect 36541 18751 36599 18757
rect 36541 18748 36553 18751
rect 36504 18720 36553 18748
rect 36504 18708 36510 18720
rect 36541 18717 36553 18720
rect 36587 18717 36599 18751
rect 36541 18711 36599 18717
rect 37734 18708 37740 18760
rect 37792 18748 37798 18760
rect 38381 18751 38439 18757
rect 38381 18748 38393 18751
rect 37792 18720 38393 18748
rect 37792 18708 37798 18720
rect 38381 18717 38393 18720
rect 38427 18717 38439 18751
rect 38381 18711 38439 18717
rect 39301 18751 39359 18757
rect 39301 18717 39313 18751
rect 39347 18717 39359 18751
rect 39301 18711 39359 18717
rect 39485 18751 39543 18757
rect 39485 18717 39497 18751
rect 39531 18748 39543 18751
rect 40034 18748 40040 18760
rect 39531 18720 40040 18748
rect 39531 18717 39543 18720
rect 39485 18711 39543 18717
rect 24854 18680 24860 18692
rect 24075 18652 24716 18680
rect 24815 18652 24860 18680
rect 24075 18649 24087 18652
rect 24029 18643 24087 18649
rect 16850 18612 16856 18624
rect 16811 18584 16856 18612
rect 16850 18572 16856 18584
rect 16908 18572 16914 18624
rect 20530 18572 20536 18624
rect 20588 18612 20594 18624
rect 20809 18615 20867 18621
rect 20809 18612 20821 18615
rect 20588 18584 20821 18612
rect 20588 18572 20594 18584
rect 20809 18581 20821 18584
rect 20855 18581 20867 18615
rect 21450 18612 21456 18624
rect 21411 18584 21456 18612
rect 20809 18575 20867 18581
rect 21450 18572 21456 18584
rect 21508 18572 21514 18624
rect 23661 18615 23719 18621
rect 23661 18581 23673 18615
rect 23707 18612 23719 18615
rect 23750 18612 23756 18624
rect 23707 18584 23756 18612
rect 23707 18581 23719 18584
rect 23661 18575 23719 18581
rect 23750 18572 23756 18584
rect 23808 18572 23814 18624
rect 23860 18612 23888 18643
rect 24854 18640 24860 18652
rect 24912 18640 24918 18692
rect 30466 18689 30472 18692
rect 24949 18683 25007 18689
rect 24949 18649 24961 18683
rect 24995 18680 25007 18683
rect 27556 18683 27614 18689
rect 24995 18652 26464 18680
rect 24995 18649 25007 18652
rect 24949 18643 25007 18649
rect 25130 18612 25136 18624
rect 23860 18584 25136 18612
rect 25130 18572 25136 18584
rect 25188 18572 25194 18624
rect 26436 18621 26464 18652
rect 27556 18649 27568 18683
rect 27602 18680 27614 18683
rect 28261 18683 28319 18689
rect 28261 18680 28273 18683
rect 27602 18652 28273 18680
rect 27602 18649 27614 18652
rect 27556 18643 27614 18649
rect 28261 18649 28273 18652
rect 28307 18649 28319 18683
rect 30460 18680 30472 18689
rect 30427 18652 30472 18680
rect 28261 18643 28319 18649
rect 30460 18643 30472 18652
rect 30466 18640 30472 18643
rect 30524 18640 30530 18692
rect 31754 18640 31760 18692
rect 31812 18680 31818 18692
rect 32033 18683 32091 18689
rect 32033 18680 32045 18683
rect 31812 18652 32045 18680
rect 31812 18640 31818 18652
rect 32033 18649 32045 18652
rect 32079 18680 32091 18683
rect 33042 18680 33048 18692
rect 32079 18652 33048 18680
rect 32079 18649 32091 18652
rect 32033 18643 32091 18649
rect 33042 18640 33048 18652
rect 33100 18680 33106 18692
rect 37645 18683 37703 18689
rect 37645 18680 37657 18683
rect 33100 18652 37657 18680
rect 33100 18640 33106 18652
rect 37645 18649 37657 18652
rect 37691 18649 37703 18683
rect 39316 18680 39344 18711
rect 40034 18708 40040 18720
rect 40092 18708 40098 18760
rect 40420 18757 40448 18788
rect 40405 18751 40463 18757
rect 40405 18717 40417 18751
rect 40451 18717 40463 18751
rect 41230 18748 41236 18760
rect 41191 18720 41236 18748
rect 40405 18711 40463 18717
rect 41230 18708 41236 18720
rect 41288 18708 41294 18760
rect 41414 18708 41420 18760
rect 41472 18748 41478 18760
rect 42076 18757 42104 18788
rect 43548 18788 44272 18816
rect 42061 18751 42119 18757
rect 41472 18720 41517 18748
rect 41472 18708 41478 18720
rect 42061 18717 42073 18751
rect 42107 18717 42119 18751
rect 42061 18711 42119 18717
rect 42245 18751 42303 18757
rect 42245 18717 42257 18751
rect 42291 18748 42303 18751
rect 42886 18748 42892 18760
rect 42291 18720 42892 18748
rect 42291 18717 42303 18720
rect 42245 18711 42303 18717
rect 40218 18680 40224 18692
rect 39316 18652 40224 18680
rect 37645 18643 37703 18649
rect 40218 18640 40224 18652
rect 40276 18640 40282 18692
rect 40586 18680 40592 18692
rect 40547 18652 40592 18680
rect 40586 18640 40592 18652
rect 40644 18640 40650 18692
rect 41874 18640 41880 18692
rect 41932 18680 41938 18692
rect 42260 18680 42288 18711
rect 42886 18708 42892 18720
rect 42944 18708 42950 18760
rect 43548 18757 43576 18788
rect 44266 18776 44272 18788
rect 44324 18776 44330 18828
rect 44358 18776 44364 18828
rect 44416 18816 44422 18828
rect 45848 18825 45876 18856
rect 46492 18856 47768 18884
rect 46492 18825 46520 18856
rect 47762 18844 47768 18856
rect 47820 18844 47826 18896
rect 45833 18819 45891 18825
rect 44416 18788 45508 18816
rect 44416 18776 44422 18788
rect 43533 18751 43591 18757
rect 43533 18717 43545 18751
rect 43579 18717 43591 18751
rect 43533 18711 43591 18717
rect 43717 18751 43775 18757
rect 43717 18717 43729 18751
rect 43763 18748 43775 18751
rect 44177 18751 44235 18757
rect 44177 18748 44189 18751
rect 43763 18720 44189 18748
rect 43763 18717 43775 18720
rect 43717 18711 43775 18717
rect 44177 18717 44189 18720
rect 44223 18717 44235 18751
rect 44634 18748 44640 18760
rect 44177 18711 44235 18717
rect 44376 18720 44640 18748
rect 41932 18652 42288 18680
rect 42904 18680 42932 18708
rect 44376 18689 44404 18720
rect 44634 18708 44640 18720
rect 44692 18708 44698 18760
rect 45370 18748 45376 18760
rect 45331 18720 45376 18748
rect 45370 18708 45376 18720
rect 45428 18708 45434 18760
rect 45480 18757 45508 18788
rect 45833 18785 45845 18819
rect 45879 18785 45891 18819
rect 45833 18779 45891 18785
rect 46477 18819 46535 18825
rect 46477 18785 46489 18819
rect 46523 18785 46535 18819
rect 46477 18779 46535 18785
rect 46661 18819 46719 18825
rect 46661 18785 46673 18819
rect 46707 18816 46719 18819
rect 47118 18816 47124 18828
rect 46707 18788 47124 18816
rect 46707 18785 46719 18788
rect 46661 18779 46719 18785
rect 47118 18776 47124 18788
rect 47176 18776 47182 18828
rect 48222 18816 48228 18828
rect 48183 18788 48228 18816
rect 48222 18776 48228 18788
rect 48280 18776 48286 18828
rect 45465 18751 45523 18757
rect 45465 18717 45477 18751
rect 45511 18717 45523 18751
rect 45465 18711 45523 18717
rect 44361 18683 44419 18689
rect 44361 18680 44373 18683
rect 42904 18652 44373 18680
rect 41932 18640 41938 18652
rect 44361 18649 44373 18652
rect 44407 18649 44419 18683
rect 44542 18680 44548 18692
rect 44503 18652 44548 18680
rect 44361 18643 44419 18649
rect 44542 18640 44548 18652
rect 44600 18640 44606 18692
rect 45554 18680 45560 18692
rect 45515 18652 45560 18680
rect 45554 18640 45560 18652
rect 45612 18640 45618 18692
rect 45646 18640 45652 18692
rect 45704 18689 45710 18692
rect 45704 18683 45753 18689
rect 45704 18649 45707 18683
rect 45741 18680 45753 18683
rect 46474 18680 46480 18692
rect 45741 18652 46480 18680
rect 45741 18649 45753 18652
rect 45704 18643 45753 18649
rect 45704 18640 45710 18643
rect 46474 18640 46480 18652
rect 46532 18640 46538 18692
rect 26421 18615 26479 18621
rect 26421 18581 26433 18615
rect 26467 18612 26479 18615
rect 27154 18612 27160 18624
rect 26467 18584 27160 18612
rect 26467 18581 26479 18584
rect 26421 18575 26479 18581
rect 27154 18572 27160 18584
rect 27212 18572 27218 18624
rect 36538 18612 36544 18624
rect 36499 18584 36544 18612
rect 36538 18572 36544 18584
rect 36596 18572 36602 18624
rect 43438 18572 43444 18624
rect 43496 18612 43502 18624
rect 43625 18615 43683 18621
rect 43625 18612 43637 18615
rect 43496 18584 43637 18612
rect 43496 18572 43502 18584
rect 43625 18581 43637 18584
rect 43671 18612 43683 18615
rect 43898 18612 43904 18624
rect 43671 18584 43904 18612
rect 43671 18581 43683 18584
rect 43625 18575 43683 18581
rect 43898 18572 43904 18584
rect 43956 18572 43962 18624
rect 45186 18612 45192 18624
rect 45147 18584 45192 18612
rect 45186 18572 45192 18584
rect 45244 18572 45250 18624
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 19978 18408 19984 18420
rect 19939 18380 19984 18408
rect 19978 18368 19984 18380
rect 20036 18368 20042 18420
rect 23934 18408 23940 18420
rect 23895 18380 23940 18408
rect 23934 18368 23940 18380
rect 23992 18368 23998 18420
rect 25038 18368 25044 18420
rect 25096 18408 25102 18420
rect 27801 18411 27859 18417
rect 25096 18380 27752 18408
rect 25096 18368 25102 18380
rect 18233 18343 18291 18349
rect 18233 18309 18245 18343
rect 18279 18340 18291 18343
rect 21450 18340 21456 18352
rect 18279 18312 21456 18340
rect 18279 18309 18291 18312
rect 18233 18303 18291 18309
rect 21450 18300 21456 18312
rect 21508 18300 21514 18352
rect 23566 18340 23572 18352
rect 23527 18312 23572 18340
rect 23566 18300 23572 18312
rect 23624 18300 23630 18352
rect 23658 18300 23664 18352
rect 23716 18340 23722 18352
rect 23769 18343 23827 18349
rect 23769 18340 23781 18343
rect 23716 18312 23781 18340
rect 23716 18300 23722 18312
rect 23769 18309 23781 18312
rect 23815 18309 23827 18343
rect 25130 18340 25136 18352
rect 23769 18303 23827 18309
rect 24412 18312 25136 18340
rect 2038 18272 2044 18284
rect 1999 18244 2044 18272
rect 2038 18232 2044 18244
rect 2096 18232 2102 18284
rect 12345 18275 12403 18281
rect 12345 18241 12357 18275
rect 12391 18272 12403 18275
rect 13081 18275 13139 18281
rect 13081 18272 13093 18275
rect 12391 18244 13093 18272
rect 12391 18241 12403 18244
rect 12345 18235 12403 18241
rect 13081 18241 13093 18244
rect 13127 18241 13139 18275
rect 13081 18235 13139 18241
rect 13265 18275 13323 18281
rect 13265 18241 13277 18275
rect 13311 18272 13323 18275
rect 13354 18272 13360 18284
rect 13311 18244 13360 18272
rect 13311 18241 13323 18244
rect 13265 18235 13323 18241
rect 13354 18232 13360 18244
rect 13412 18232 13418 18284
rect 13538 18272 13544 18284
rect 13499 18244 13544 18272
rect 13538 18232 13544 18244
rect 13596 18232 13602 18284
rect 13722 18272 13728 18284
rect 13683 18244 13728 18272
rect 13722 18232 13728 18244
rect 13780 18232 13786 18284
rect 16114 18272 16120 18284
rect 16075 18244 16120 18272
rect 16114 18232 16120 18244
rect 16172 18232 16178 18284
rect 16298 18272 16304 18284
rect 16259 18244 16304 18272
rect 16298 18232 16304 18244
rect 16356 18232 16362 18284
rect 17126 18232 17132 18284
rect 17184 18272 17190 18284
rect 17957 18275 18015 18281
rect 17957 18272 17969 18275
rect 17184 18244 17969 18272
rect 17184 18232 17190 18244
rect 17957 18241 17969 18244
rect 18003 18241 18015 18275
rect 17957 18235 18015 18241
rect 18141 18275 18199 18281
rect 18141 18241 18153 18275
rect 18187 18241 18199 18275
rect 18322 18272 18328 18284
rect 18283 18244 18328 18272
rect 18141 18235 18199 18241
rect 2222 18204 2228 18216
rect 2183 18176 2228 18204
rect 2222 18164 2228 18176
rect 2280 18164 2286 18216
rect 2774 18164 2780 18216
rect 2832 18204 2838 18216
rect 12161 18207 12219 18213
rect 2832 18176 2877 18204
rect 2832 18164 2838 18176
rect 12161 18173 12173 18207
rect 12207 18204 12219 18207
rect 12526 18204 12532 18216
rect 12207 18176 12532 18204
rect 12207 18173 12219 18176
rect 12161 18167 12219 18173
rect 12526 18164 12532 18176
rect 12584 18164 12590 18216
rect 12618 18164 12624 18216
rect 12676 18204 12682 18216
rect 13556 18204 13584 18232
rect 14734 18204 14740 18216
rect 12676 18176 12721 18204
rect 13556 18176 14740 18204
rect 12676 18164 12682 18176
rect 14734 18164 14740 18176
rect 14792 18164 14798 18216
rect 18156 18204 18184 18235
rect 18322 18232 18328 18244
rect 18380 18232 18386 18284
rect 20162 18272 20168 18284
rect 20123 18244 20168 18272
rect 20162 18232 20168 18244
rect 20220 18232 20226 18284
rect 20441 18275 20499 18281
rect 20441 18241 20453 18275
rect 20487 18241 20499 18275
rect 20441 18235 20499 18241
rect 20456 18204 20484 18235
rect 20530 18232 20536 18284
rect 20588 18272 20594 18284
rect 20625 18275 20683 18281
rect 20625 18272 20637 18275
rect 20588 18244 20637 18272
rect 20588 18232 20594 18244
rect 20625 18241 20637 18244
rect 20671 18241 20683 18275
rect 23584 18272 23612 18300
rect 24026 18272 24032 18284
rect 23584 18244 24032 18272
rect 20625 18235 20683 18241
rect 24026 18232 24032 18244
rect 24084 18232 24090 18284
rect 24412 18281 24440 18312
rect 25130 18300 25136 18312
rect 25188 18300 25194 18352
rect 27724 18340 27752 18380
rect 27801 18377 27813 18411
rect 27847 18408 27859 18411
rect 28442 18408 28448 18420
rect 27847 18380 28448 18408
rect 27847 18377 27859 18380
rect 27801 18371 27859 18377
rect 28442 18368 28448 18380
rect 28500 18368 28506 18420
rect 30650 18368 30656 18420
rect 30708 18408 30714 18420
rect 30929 18411 30987 18417
rect 30929 18408 30941 18411
rect 30708 18380 30941 18408
rect 30708 18368 30714 18380
rect 30929 18377 30941 18380
rect 30975 18377 30987 18411
rect 34790 18408 34796 18420
rect 30929 18371 30987 18377
rect 33980 18380 34796 18408
rect 29730 18340 29736 18352
rect 27724 18312 29736 18340
rect 29730 18300 29736 18312
rect 29788 18300 29794 18352
rect 24397 18275 24455 18281
rect 24397 18241 24409 18275
rect 24443 18241 24455 18275
rect 24397 18235 24455 18241
rect 24581 18275 24639 18281
rect 24581 18241 24593 18275
rect 24627 18272 24639 18275
rect 24762 18272 24768 18284
rect 24627 18244 24768 18272
rect 24627 18241 24639 18244
rect 24581 18235 24639 18241
rect 24762 18232 24768 18244
rect 24820 18232 24826 18284
rect 27154 18272 27160 18284
rect 27115 18244 27160 18272
rect 27154 18232 27160 18244
rect 27212 18232 27218 18284
rect 27246 18232 27252 18284
rect 27304 18272 27310 18284
rect 27341 18275 27399 18281
rect 27341 18272 27353 18275
rect 27304 18244 27353 18272
rect 27304 18232 27310 18244
rect 27341 18241 27353 18244
rect 27387 18272 27399 18275
rect 27522 18272 27528 18284
rect 27387 18244 27528 18272
rect 27387 18241 27399 18244
rect 27341 18235 27399 18241
rect 27522 18232 27528 18244
rect 27580 18232 27586 18284
rect 27617 18275 27675 18281
rect 27617 18241 27629 18275
rect 27663 18272 27675 18275
rect 27706 18272 27712 18284
rect 27663 18244 27712 18272
rect 27663 18241 27675 18244
rect 27617 18235 27675 18241
rect 27706 18232 27712 18244
rect 27764 18232 27770 18284
rect 29822 18232 29828 18284
rect 29880 18272 29886 18284
rect 30285 18275 30343 18281
rect 30285 18272 30297 18275
rect 29880 18244 30297 18272
rect 29880 18232 29886 18244
rect 30285 18241 30297 18244
rect 30331 18241 30343 18275
rect 30285 18235 30343 18241
rect 30469 18275 30527 18281
rect 30469 18241 30481 18275
rect 30515 18272 30527 18275
rect 30558 18272 30564 18284
rect 30515 18244 30564 18272
rect 30515 18241 30527 18244
rect 30469 18235 30527 18241
rect 30558 18232 30564 18244
rect 30616 18232 30622 18284
rect 30742 18272 30748 18284
rect 30703 18244 30748 18272
rect 30742 18232 30748 18244
rect 30800 18232 30806 18284
rect 33778 18272 33784 18284
rect 33739 18244 33784 18272
rect 33778 18232 33784 18244
rect 33836 18232 33842 18284
rect 33980 18281 34008 18380
rect 34790 18368 34796 18380
rect 34848 18408 34854 18420
rect 36909 18411 36967 18417
rect 34848 18380 36676 18408
rect 34848 18368 34854 18380
rect 34422 18300 34428 18352
rect 34480 18340 34486 18352
rect 34885 18343 34943 18349
rect 34480 18312 34744 18340
rect 34480 18300 34486 18312
rect 34716 18281 34744 18312
rect 34885 18309 34897 18343
rect 34931 18340 34943 18343
rect 35713 18343 35771 18349
rect 35713 18340 35725 18343
rect 34931 18312 35725 18340
rect 34931 18309 34943 18312
rect 34885 18303 34943 18309
rect 35713 18309 35725 18312
rect 35759 18309 35771 18343
rect 36538 18340 36544 18352
rect 36499 18312 36544 18340
rect 35713 18303 35771 18309
rect 36538 18300 36544 18312
rect 36596 18300 36602 18352
rect 36648 18349 36676 18380
rect 36909 18377 36921 18411
rect 36955 18377 36967 18411
rect 40402 18408 40408 18420
rect 40363 18380 40408 18408
rect 36909 18371 36967 18377
rect 36633 18343 36691 18349
rect 36633 18309 36645 18343
rect 36679 18309 36691 18343
rect 36633 18303 36691 18309
rect 33965 18275 34023 18281
rect 33965 18241 33977 18275
rect 34011 18241 34023 18275
rect 33965 18235 34023 18241
rect 34517 18275 34575 18281
rect 34517 18241 34529 18275
rect 34563 18241 34575 18275
rect 34517 18235 34575 18241
rect 34609 18275 34667 18281
rect 34609 18241 34621 18275
rect 34655 18241 34667 18275
rect 34609 18235 34667 18241
rect 34701 18275 34759 18281
rect 34701 18241 34713 18275
rect 34747 18241 34759 18275
rect 36354 18272 36360 18284
rect 36315 18244 36360 18272
rect 34701 18235 34759 18241
rect 21266 18204 21272 18216
rect 18156 18176 19334 18204
rect 20456 18176 21272 18204
rect 19306 18136 19334 18176
rect 21266 18164 21272 18176
rect 21324 18164 21330 18216
rect 21634 18136 21640 18148
rect 19306 18108 21640 18136
rect 21634 18096 21640 18108
rect 21692 18136 21698 18148
rect 24854 18136 24860 18148
rect 21692 18108 24860 18136
rect 21692 18096 21698 18108
rect 24854 18096 24860 18108
rect 24912 18096 24918 18148
rect 12529 18071 12587 18077
rect 12529 18037 12541 18071
rect 12575 18068 12587 18071
rect 12710 18068 12716 18080
rect 12575 18040 12716 18068
rect 12575 18037 12587 18040
rect 12529 18031 12587 18037
rect 12710 18028 12716 18040
rect 12768 18028 12774 18080
rect 16209 18071 16267 18077
rect 16209 18037 16221 18071
rect 16255 18068 16267 18071
rect 16574 18068 16580 18080
rect 16255 18040 16580 18068
rect 16255 18037 16267 18040
rect 16209 18031 16267 18037
rect 16574 18028 16580 18040
rect 16632 18028 16638 18080
rect 18322 18028 18328 18080
rect 18380 18068 18386 18080
rect 18509 18071 18567 18077
rect 18509 18068 18521 18071
rect 18380 18040 18521 18068
rect 18380 18028 18386 18040
rect 18509 18037 18521 18040
rect 18555 18037 18567 18071
rect 18509 18031 18567 18037
rect 23753 18071 23811 18077
rect 23753 18037 23765 18071
rect 23799 18068 23811 18071
rect 23842 18068 23848 18080
rect 23799 18040 23848 18068
rect 23799 18037 23811 18040
rect 23753 18031 23811 18037
rect 23842 18028 23848 18040
rect 23900 18028 23906 18080
rect 23934 18028 23940 18080
rect 23992 18068 23998 18080
rect 24489 18071 24547 18077
rect 24489 18068 24501 18071
rect 23992 18040 24501 18068
rect 23992 18028 23998 18040
rect 24489 18037 24501 18040
rect 24535 18037 24547 18071
rect 33962 18068 33968 18080
rect 33923 18040 33968 18068
rect 24489 18031 24547 18037
rect 33962 18028 33968 18040
rect 34020 18068 34026 18080
rect 34532 18068 34560 18235
rect 34624 18136 34652 18235
rect 36354 18232 36360 18244
rect 36412 18232 36418 18284
rect 34698 18136 34704 18148
rect 34624 18108 34704 18136
rect 34698 18096 34704 18108
rect 34756 18096 34762 18148
rect 35342 18136 35348 18148
rect 35303 18108 35348 18136
rect 35342 18096 35348 18108
rect 35400 18096 35406 18148
rect 36170 18136 36176 18148
rect 35728 18108 36176 18136
rect 35728 18077 35756 18108
rect 36170 18096 36176 18108
rect 36228 18096 36234 18148
rect 36648 18136 36676 18303
rect 36725 18275 36783 18281
rect 36725 18241 36737 18275
rect 36771 18241 36783 18275
rect 36924 18272 36952 18371
rect 40402 18368 40408 18380
rect 40460 18368 40466 18420
rect 43717 18411 43775 18417
rect 43717 18377 43729 18411
rect 43763 18408 43775 18411
rect 44358 18408 44364 18420
rect 43763 18380 44364 18408
rect 43763 18377 43775 18380
rect 43717 18371 43775 18377
rect 44358 18368 44364 18380
rect 44416 18368 44422 18420
rect 45462 18368 45468 18420
rect 45520 18408 45526 18420
rect 46017 18411 46075 18417
rect 46017 18408 46029 18411
rect 45520 18380 46029 18408
rect 45520 18368 45526 18380
rect 46017 18377 46029 18380
rect 46063 18377 46075 18411
rect 46017 18371 46075 18377
rect 37734 18300 37740 18352
rect 37792 18340 37798 18352
rect 40034 18340 40040 18352
rect 37792 18312 38884 18340
rect 39995 18312 40040 18340
rect 37792 18300 37798 18312
rect 38856 18281 38884 18312
rect 40034 18300 40040 18312
rect 40092 18300 40098 18352
rect 40218 18340 40224 18352
rect 40179 18312 40224 18340
rect 40218 18300 40224 18312
rect 40276 18340 40282 18352
rect 41598 18340 41604 18352
rect 40276 18312 41604 18340
rect 40276 18300 40282 18312
rect 41598 18300 41604 18312
rect 41656 18300 41662 18352
rect 44085 18343 44143 18349
rect 44085 18309 44097 18343
rect 44131 18340 44143 18343
rect 44266 18340 44272 18352
rect 44131 18312 44272 18340
rect 44131 18309 44143 18312
rect 44085 18303 44143 18309
rect 44266 18300 44272 18312
rect 44324 18300 44330 18352
rect 44904 18343 44962 18349
rect 44904 18309 44916 18343
rect 44950 18340 44962 18343
rect 45186 18340 45192 18352
rect 44950 18312 45192 18340
rect 44950 18309 44962 18312
rect 44904 18303 44962 18309
rect 45186 18300 45192 18312
rect 45244 18300 45250 18352
rect 38574 18275 38632 18281
rect 38574 18272 38586 18275
rect 36924 18244 38586 18272
rect 36725 18235 36783 18241
rect 38574 18241 38586 18244
rect 38620 18241 38632 18275
rect 38574 18235 38632 18241
rect 38841 18275 38899 18281
rect 38841 18241 38853 18275
rect 38887 18241 38899 18275
rect 41138 18272 41144 18284
rect 41099 18244 41144 18272
rect 38841 18235 38899 18241
rect 36740 18204 36768 18235
rect 38856 18204 38884 18235
rect 41138 18232 41144 18244
rect 41196 18232 41202 18284
rect 43898 18272 43904 18284
rect 43859 18244 43904 18272
rect 43898 18232 43904 18244
rect 43956 18232 43962 18284
rect 44177 18275 44235 18281
rect 44177 18241 44189 18275
rect 44223 18272 44235 18275
rect 45462 18272 45468 18284
rect 44223 18244 45468 18272
rect 44223 18241 44235 18244
rect 44177 18235 44235 18241
rect 45462 18232 45468 18244
rect 45520 18232 45526 18284
rect 44637 18207 44695 18213
rect 44637 18204 44649 18207
rect 36740 18176 37596 18204
rect 38856 18176 44649 18204
rect 37461 18139 37519 18145
rect 37461 18136 37473 18139
rect 36648 18108 37473 18136
rect 37461 18105 37473 18108
rect 37507 18105 37519 18139
rect 37461 18099 37519 18105
rect 34020 18040 34560 18068
rect 35713 18071 35771 18077
rect 34020 18028 34026 18040
rect 35713 18037 35725 18071
rect 35759 18037 35771 18071
rect 35713 18031 35771 18037
rect 35897 18071 35955 18077
rect 35897 18037 35909 18071
rect 35943 18068 35955 18071
rect 36078 18068 36084 18080
rect 35943 18040 36084 18068
rect 35943 18037 35955 18040
rect 35897 18031 35955 18037
rect 36078 18028 36084 18040
rect 36136 18028 36142 18080
rect 37568 18068 37596 18176
rect 44637 18173 44649 18176
rect 44683 18173 44695 18207
rect 44637 18167 44695 18173
rect 40678 18068 40684 18080
rect 37568 18040 40684 18068
rect 40678 18028 40684 18040
rect 40736 18028 40742 18080
rect 41322 18068 41328 18080
rect 41283 18040 41328 18068
rect 41322 18028 41328 18040
rect 41380 18028 41386 18080
rect 43898 18028 43904 18080
rect 43956 18068 43962 18080
rect 44634 18068 44640 18080
rect 43956 18040 44640 18068
rect 43956 18028 43962 18040
rect 44634 18028 44640 18040
rect 44692 18028 44698 18080
rect 47949 18071 48007 18077
rect 47949 18037 47961 18071
rect 47995 18068 48007 18071
rect 48314 18068 48320 18080
rect 47995 18040 48320 18068
rect 47995 18037 48007 18040
rect 47949 18031 48007 18037
rect 48314 18028 48320 18040
rect 48372 18028 48378 18080
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 2222 17824 2228 17876
rect 2280 17864 2286 17876
rect 2317 17867 2375 17873
rect 2317 17864 2329 17867
rect 2280 17836 2329 17864
rect 2280 17824 2286 17836
rect 2317 17833 2329 17836
rect 2363 17833 2375 17867
rect 2317 17827 2375 17833
rect 11425 17867 11483 17873
rect 11425 17833 11437 17867
rect 11471 17864 11483 17867
rect 12618 17864 12624 17876
rect 11471 17836 12624 17864
rect 11471 17833 11483 17836
rect 11425 17827 11483 17833
rect 12618 17824 12624 17836
rect 12676 17824 12682 17876
rect 13633 17867 13691 17873
rect 13633 17833 13645 17867
rect 13679 17864 13691 17867
rect 13722 17864 13728 17876
rect 13679 17836 13728 17864
rect 13679 17833 13691 17836
rect 13633 17827 13691 17833
rect 13722 17824 13728 17836
rect 13780 17824 13786 17876
rect 15473 17867 15531 17873
rect 15473 17833 15485 17867
rect 15519 17864 15531 17867
rect 15930 17864 15936 17876
rect 15519 17836 15936 17864
rect 15519 17833 15531 17836
rect 15473 17827 15531 17833
rect 15930 17824 15936 17836
rect 15988 17864 15994 17876
rect 16114 17864 16120 17876
rect 15988 17836 16120 17864
rect 15988 17824 15994 17836
rect 16114 17824 16120 17836
rect 16172 17824 16178 17876
rect 16209 17867 16267 17873
rect 16209 17833 16221 17867
rect 16255 17864 16267 17867
rect 16298 17864 16304 17876
rect 16255 17836 16304 17864
rect 16255 17833 16267 17836
rect 16209 17827 16267 17833
rect 16298 17824 16304 17836
rect 16356 17824 16362 17876
rect 17126 17864 17132 17876
rect 17087 17836 17132 17864
rect 17126 17824 17132 17836
rect 17184 17824 17190 17876
rect 19242 17864 19248 17876
rect 17512 17836 19248 17864
rect 17512 17796 17540 17836
rect 19242 17824 19248 17836
rect 19300 17824 19306 17876
rect 19521 17867 19579 17873
rect 19521 17833 19533 17867
rect 19567 17864 19579 17867
rect 21082 17864 21088 17876
rect 19567 17836 21088 17864
rect 19567 17833 19579 17836
rect 19521 17827 19579 17833
rect 21082 17824 21088 17836
rect 21140 17824 21146 17876
rect 23293 17867 23351 17873
rect 23293 17833 23305 17867
rect 23339 17864 23351 17867
rect 23658 17864 23664 17876
rect 23339 17836 23664 17864
rect 23339 17833 23351 17836
rect 23293 17827 23351 17833
rect 23658 17824 23664 17836
rect 23716 17824 23722 17876
rect 28813 17867 28871 17873
rect 28813 17833 28825 17867
rect 28859 17864 28871 17867
rect 28902 17864 28908 17876
rect 28859 17836 28908 17864
rect 28859 17833 28871 17836
rect 28813 17827 28871 17833
rect 28902 17824 28908 17836
rect 28960 17824 28966 17876
rect 31849 17867 31907 17873
rect 31849 17864 31861 17867
rect 31726 17836 31861 17864
rect 14292 17768 17540 17796
rect 11333 17731 11391 17737
rect 11333 17697 11345 17731
rect 11379 17697 11391 17731
rect 11333 17691 11391 17697
rect 2409 17663 2467 17669
rect 2409 17629 2421 17663
rect 2455 17660 2467 17663
rect 2590 17660 2596 17672
rect 2455 17632 2596 17660
rect 2455 17629 2467 17632
rect 2409 17623 2467 17629
rect 2590 17620 2596 17632
rect 2648 17660 2654 17672
rect 6730 17660 6736 17672
rect 2648 17632 6736 17660
rect 2648 17620 2654 17632
rect 6730 17620 6736 17632
rect 6788 17620 6794 17672
rect 11348 17592 11376 17691
rect 11609 17663 11667 17669
rect 11609 17629 11621 17663
rect 11655 17660 11667 17663
rect 12066 17660 12072 17672
rect 11655 17632 12072 17660
rect 11655 17629 11667 17632
rect 11609 17623 11667 17629
rect 12066 17620 12072 17632
rect 12124 17620 12130 17672
rect 12250 17620 12256 17672
rect 12308 17660 12314 17672
rect 12894 17660 12900 17672
rect 12308 17632 12353 17660
rect 12406 17632 12900 17660
rect 12308 17620 12314 17632
rect 12406 17592 12434 17632
rect 12894 17620 12900 17632
rect 12952 17660 12958 17672
rect 14292 17660 14320 17768
rect 16850 17728 16856 17740
rect 16408 17700 16856 17728
rect 14458 17660 14464 17672
rect 12952 17632 14320 17660
rect 14419 17632 14464 17660
rect 12952 17620 12958 17632
rect 14458 17620 14464 17632
rect 14516 17620 14522 17672
rect 14734 17660 14740 17672
rect 14695 17632 14740 17660
rect 14734 17620 14740 17632
rect 14792 17620 14798 17672
rect 14921 17663 14979 17669
rect 14921 17629 14933 17663
rect 14967 17629 14979 17663
rect 14921 17623 14979 17629
rect 12526 17601 12532 17604
rect 11348 17564 12434 17592
rect 12520 17555 12532 17601
rect 12584 17592 12590 17604
rect 14277 17595 14335 17601
rect 14277 17592 14289 17595
rect 12584 17564 12620 17592
rect 12728 17564 14289 17592
rect 12526 17552 12532 17555
rect 12584 17552 12590 17564
rect 11793 17527 11851 17533
rect 11793 17493 11805 17527
rect 11839 17524 11851 17527
rect 11974 17524 11980 17536
rect 11839 17496 11980 17524
rect 11839 17493 11851 17496
rect 11793 17487 11851 17493
rect 11974 17484 11980 17496
rect 12032 17484 12038 17536
rect 12066 17484 12072 17536
rect 12124 17524 12130 17536
rect 12728 17524 12756 17564
rect 14277 17561 14289 17564
rect 14323 17561 14335 17595
rect 14277 17555 14335 17561
rect 12124 17496 12756 17524
rect 12124 17484 12130 17496
rect 13262 17484 13268 17536
rect 13320 17524 13326 17536
rect 14936 17524 14964 17623
rect 15102 17620 15108 17672
rect 15160 17660 15166 17672
rect 16408 17669 16436 17700
rect 16850 17688 16856 17700
rect 16908 17688 16914 17740
rect 18509 17731 18567 17737
rect 18509 17697 18521 17731
rect 18555 17728 18567 17731
rect 19334 17728 19340 17740
rect 18555 17700 19340 17728
rect 18555 17697 18567 17700
rect 18509 17691 18567 17697
rect 19334 17688 19340 17700
rect 19392 17728 19398 17740
rect 23017 17731 23075 17737
rect 19392 17700 20392 17728
rect 19392 17688 19398 17700
rect 15381 17663 15439 17669
rect 15381 17660 15393 17663
rect 15160 17632 15393 17660
rect 15160 17620 15166 17632
rect 15381 17629 15393 17632
rect 15427 17629 15439 17663
rect 15381 17623 15439 17629
rect 15565 17663 15623 17669
rect 15565 17629 15577 17663
rect 15611 17629 15623 17663
rect 15565 17623 15623 17629
rect 16393 17663 16451 17669
rect 16393 17629 16405 17663
rect 16439 17629 16451 17663
rect 16666 17660 16672 17672
rect 16627 17632 16672 17660
rect 16393 17623 16451 17629
rect 15194 17552 15200 17604
rect 15252 17592 15258 17604
rect 15580 17592 15608 17623
rect 16666 17620 16672 17632
rect 16724 17620 16730 17672
rect 19426 17660 19432 17672
rect 19387 17632 19432 17660
rect 19426 17620 19432 17632
rect 19484 17620 19490 17672
rect 19705 17663 19763 17669
rect 19705 17629 19717 17663
rect 19751 17660 19763 17663
rect 20254 17660 20260 17672
rect 19751 17632 20260 17660
rect 19751 17629 19763 17632
rect 19705 17623 19763 17629
rect 20254 17620 20260 17632
rect 20312 17620 20318 17672
rect 20364 17669 20392 17700
rect 23017 17697 23029 17731
rect 23063 17728 23075 17731
rect 23198 17728 23204 17740
rect 23063 17700 23204 17728
rect 23063 17697 23075 17700
rect 23017 17691 23075 17697
rect 23198 17688 23204 17700
rect 23256 17688 23262 17740
rect 28721 17731 28779 17737
rect 28721 17697 28733 17731
rect 28767 17728 28779 17731
rect 29454 17728 29460 17740
rect 28767 17700 29460 17728
rect 28767 17697 28779 17700
rect 28721 17691 28779 17697
rect 29454 17688 29460 17700
rect 29512 17688 29518 17740
rect 31389 17731 31447 17737
rect 31389 17697 31401 17731
rect 31435 17728 31447 17731
rect 31726 17728 31754 17836
rect 31849 17833 31861 17836
rect 31895 17864 31907 17867
rect 33778 17864 33784 17876
rect 31895 17836 33784 17864
rect 31895 17833 31907 17836
rect 31849 17827 31907 17833
rect 33778 17824 33784 17836
rect 33836 17824 33842 17876
rect 35253 17867 35311 17873
rect 35253 17833 35265 17867
rect 35299 17864 35311 17867
rect 35342 17864 35348 17876
rect 35299 17836 35348 17864
rect 35299 17833 35311 17836
rect 35253 17827 35311 17833
rect 35342 17824 35348 17836
rect 35400 17824 35406 17876
rect 36354 17824 36360 17876
rect 36412 17864 36418 17876
rect 36633 17867 36691 17873
rect 36633 17864 36645 17867
rect 36412 17836 36645 17864
rect 36412 17824 36418 17836
rect 36633 17833 36645 17836
rect 36679 17833 36691 17867
rect 40034 17864 40040 17876
rect 39995 17836 40040 17864
rect 36633 17827 36691 17833
rect 40034 17824 40040 17836
rect 40092 17824 40098 17876
rect 43901 17867 43959 17873
rect 43901 17833 43913 17867
rect 43947 17864 43959 17867
rect 44542 17864 44548 17876
rect 43947 17836 44548 17864
rect 43947 17833 43959 17836
rect 43901 17827 43959 17833
rect 44542 17824 44548 17836
rect 44600 17824 44606 17876
rect 45370 17864 45376 17876
rect 45331 17836 45376 17864
rect 45370 17824 45376 17836
rect 45428 17824 45434 17876
rect 36265 17799 36323 17805
rect 36265 17765 36277 17799
rect 36311 17796 36323 17799
rect 36446 17796 36452 17808
rect 36311 17768 36452 17796
rect 36311 17765 36323 17768
rect 36265 17759 36323 17765
rect 36446 17756 36452 17768
rect 36504 17756 36510 17808
rect 43809 17799 43867 17805
rect 43809 17765 43821 17799
rect 43855 17796 43867 17799
rect 44358 17796 44364 17808
rect 43855 17768 44364 17796
rect 43855 17765 43867 17768
rect 43809 17759 43867 17765
rect 44358 17756 44364 17768
rect 44416 17756 44422 17808
rect 31435 17700 31754 17728
rect 33229 17731 33287 17737
rect 31435 17697 31447 17700
rect 31389 17691 31447 17697
rect 33229 17697 33241 17731
rect 33275 17728 33287 17731
rect 37734 17728 37740 17740
rect 33275 17700 37740 17728
rect 33275 17697 33287 17700
rect 33229 17691 33287 17697
rect 37734 17688 37740 17700
rect 37792 17688 37798 17740
rect 43993 17731 44051 17737
rect 43993 17697 44005 17731
rect 44039 17728 44051 17731
rect 44450 17728 44456 17740
rect 44039 17700 44456 17728
rect 44039 17697 44051 17700
rect 43993 17691 44051 17697
rect 44450 17688 44456 17700
rect 44508 17688 44514 17740
rect 46842 17728 46848 17740
rect 46803 17700 46848 17728
rect 46842 17688 46848 17700
rect 46900 17688 46906 17740
rect 48314 17728 48320 17740
rect 48275 17700 48320 17728
rect 48314 17688 48320 17700
rect 48372 17688 48378 17740
rect 20349 17663 20407 17669
rect 20349 17629 20361 17663
rect 20395 17660 20407 17663
rect 20438 17660 20444 17672
rect 20395 17632 20444 17660
rect 20395 17629 20407 17632
rect 20349 17623 20407 17629
rect 20438 17620 20444 17632
rect 20496 17620 20502 17672
rect 22925 17663 22983 17669
rect 22925 17629 22937 17663
rect 22971 17629 22983 17663
rect 23750 17660 23756 17672
rect 23711 17632 23756 17660
rect 22925 17623 22983 17629
rect 15252 17564 15608 17592
rect 18264 17595 18322 17601
rect 15252 17552 15258 17564
rect 18264 17561 18276 17595
rect 18310 17592 18322 17595
rect 18506 17592 18512 17604
rect 18310 17564 18512 17592
rect 18310 17561 18322 17564
rect 18264 17555 18322 17561
rect 18506 17552 18512 17564
rect 18564 17552 18570 17604
rect 19889 17595 19947 17601
rect 19889 17561 19901 17595
rect 19935 17592 19947 17595
rect 20594 17595 20652 17601
rect 20594 17592 20606 17595
rect 19935 17564 20606 17592
rect 19935 17561 19947 17564
rect 19889 17555 19947 17561
rect 20594 17561 20606 17564
rect 20640 17561 20652 17595
rect 22940 17592 22968 17623
rect 23750 17620 23756 17632
rect 23808 17620 23814 17672
rect 23934 17660 23940 17672
rect 23895 17632 23940 17660
rect 23934 17620 23940 17632
rect 23992 17620 23998 17672
rect 28997 17663 29055 17669
rect 28997 17629 29009 17663
rect 29043 17660 29055 17663
rect 29733 17663 29791 17669
rect 29733 17660 29745 17663
rect 29043 17632 29745 17660
rect 29043 17629 29055 17632
rect 28997 17623 29055 17629
rect 29733 17629 29745 17632
rect 29779 17629 29791 17663
rect 29733 17623 29791 17629
rect 29914 17620 29920 17672
rect 29972 17660 29978 17672
rect 30190 17660 30196 17672
rect 29972 17632 30065 17660
rect 30151 17632 30196 17660
rect 29972 17620 29978 17632
rect 30190 17620 30196 17632
rect 30248 17620 30254 17672
rect 30377 17663 30435 17669
rect 30377 17629 30389 17663
rect 30423 17629 30435 17663
rect 31110 17660 31116 17672
rect 31071 17632 31116 17660
rect 30377 17623 30435 17629
rect 23474 17592 23480 17604
rect 20594 17555 20652 17561
rect 21560 17564 22094 17592
rect 22940 17564 23480 17592
rect 13320 17496 14964 17524
rect 16577 17527 16635 17533
rect 13320 17484 13326 17496
rect 16577 17493 16589 17527
rect 16623 17524 16635 17527
rect 16942 17524 16948 17536
rect 16623 17496 16948 17524
rect 16623 17493 16635 17496
rect 16577 17487 16635 17493
rect 16942 17484 16948 17496
rect 17000 17484 17006 17536
rect 19426 17484 19432 17536
rect 19484 17524 19490 17536
rect 21560 17524 21588 17564
rect 21726 17524 21732 17536
rect 19484 17496 21588 17524
rect 21687 17496 21732 17524
rect 19484 17484 19490 17496
rect 21726 17484 21732 17496
rect 21784 17484 21790 17536
rect 22066 17524 22094 17564
rect 23474 17552 23480 17564
rect 23532 17592 23538 17604
rect 23845 17595 23903 17601
rect 23845 17592 23857 17595
rect 23532 17564 23857 17592
rect 23532 17552 23538 17564
rect 23845 17561 23857 17564
rect 23891 17561 23903 17595
rect 29932 17592 29960 17620
rect 30282 17592 30288 17604
rect 29932 17564 30288 17592
rect 23845 17555 23903 17561
rect 30282 17552 30288 17564
rect 30340 17552 30346 17604
rect 28994 17524 29000 17536
rect 22066 17496 29000 17524
rect 28994 17484 29000 17496
rect 29052 17484 29058 17536
rect 29178 17524 29184 17536
rect 29139 17496 29184 17524
rect 29178 17484 29184 17496
rect 29236 17484 29242 17536
rect 30098 17484 30104 17536
rect 30156 17524 30162 17536
rect 30392 17524 30420 17623
rect 31110 17620 31116 17632
rect 31168 17620 31174 17672
rect 31294 17620 31300 17672
rect 31352 17660 31358 17672
rect 31570 17660 31576 17672
rect 31352 17632 31576 17660
rect 31352 17620 31358 17632
rect 31570 17620 31576 17632
rect 31628 17620 31634 17672
rect 33778 17620 33784 17672
rect 33836 17660 33842 17672
rect 34885 17663 34943 17669
rect 34885 17660 34897 17663
rect 33836 17632 34897 17660
rect 33836 17620 33842 17632
rect 34885 17629 34897 17632
rect 34931 17629 34943 17663
rect 34885 17623 34943 17629
rect 35069 17663 35127 17669
rect 35069 17629 35081 17663
rect 35115 17629 35127 17663
rect 35069 17623 35127 17629
rect 36173 17663 36231 17669
rect 36173 17629 36185 17663
rect 36219 17629 36231 17663
rect 36173 17623 36231 17629
rect 30929 17595 30987 17601
rect 30929 17561 30941 17595
rect 30975 17592 30987 17595
rect 32962 17595 33020 17601
rect 32962 17592 32974 17595
rect 30975 17564 32974 17592
rect 30975 17561 30987 17564
rect 30929 17555 30987 17561
rect 32962 17561 32974 17564
rect 33008 17561 33020 17595
rect 32962 17555 33020 17561
rect 34790 17552 34796 17604
rect 34848 17592 34854 17604
rect 35084 17592 35112 17623
rect 34848 17564 35112 17592
rect 34848 17552 34854 17564
rect 36188 17524 36216 17623
rect 36354 17620 36360 17672
rect 36412 17660 36418 17672
rect 36449 17663 36507 17669
rect 36449 17660 36461 17663
rect 36412 17632 36461 17660
rect 36412 17620 36418 17632
rect 36449 17629 36461 17632
rect 36495 17629 36507 17663
rect 36449 17623 36507 17629
rect 40221 17663 40279 17669
rect 40221 17629 40233 17663
rect 40267 17660 40279 17663
rect 40310 17660 40316 17672
rect 40267 17632 40316 17660
rect 40267 17629 40279 17632
rect 40221 17623 40279 17629
rect 40310 17620 40316 17632
rect 40368 17620 40374 17672
rect 40497 17663 40555 17669
rect 40497 17629 40509 17663
rect 40543 17660 40555 17663
rect 41322 17660 41328 17672
rect 40543 17632 41184 17660
rect 41283 17632 41328 17660
rect 40543 17629 40555 17632
rect 40497 17623 40555 17629
rect 40954 17592 40960 17604
rect 40915 17564 40960 17592
rect 40954 17552 40960 17564
rect 41012 17552 41018 17604
rect 41156 17536 41184 17632
rect 41322 17620 41328 17632
rect 41380 17620 41386 17672
rect 43714 17660 43720 17672
rect 43675 17632 43720 17660
rect 43714 17620 43720 17632
rect 43772 17620 43778 17672
rect 44109 17663 44167 17669
rect 44109 17660 44121 17663
rect 44100 17629 44121 17660
rect 44155 17629 44167 17663
rect 44100 17623 44167 17629
rect 41233 17595 41291 17601
rect 41233 17561 41245 17595
rect 41279 17592 41291 17595
rect 41598 17592 41604 17604
rect 41279 17564 41604 17592
rect 41279 17561 41291 17564
rect 41233 17555 41291 17561
rect 41598 17552 41604 17564
rect 41656 17552 41662 17604
rect 30156 17496 36216 17524
rect 30156 17484 30162 17496
rect 40126 17484 40132 17536
rect 40184 17524 40190 17536
rect 40405 17527 40463 17533
rect 40405 17524 40417 17527
rect 40184 17496 40417 17524
rect 40184 17484 40190 17496
rect 40405 17493 40417 17496
rect 40451 17493 40463 17527
rect 41138 17524 41144 17536
rect 41099 17496 41144 17524
rect 40405 17487 40463 17493
rect 41138 17484 41144 17496
rect 41196 17484 41202 17536
rect 41506 17524 41512 17536
rect 41467 17496 41512 17524
rect 41506 17484 41512 17496
rect 41564 17484 41570 17536
rect 43346 17484 43352 17536
rect 43404 17524 43410 17536
rect 43441 17527 43499 17533
rect 43441 17524 43453 17527
rect 43404 17496 43453 17524
rect 43404 17484 43410 17496
rect 43441 17493 43453 17496
rect 43487 17493 43499 17527
rect 44100 17524 44128 17623
rect 44634 17620 44640 17672
rect 44692 17660 44698 17672
rect 45189 17663 45247 17669
rect 45189 17660 45201 17663
rect 44692 17632 45201 17660
rect 44692 17620 44698 17632
rect 45189 17629 45201 17632
rect 45235 17629 45247 17663
rect 45462 17660 45468 17672
rect 45423 17632 45468 17660
rect 45189 17623 45247 17629
rect 45462 17620 45468 17632
rect 45520 17620 45526 17672
rect 44266 17552 44272 17604
rect 44324 17592 44330 17604
rect 45281 17595 45339 17601
rect 45281 17592 45293 17595
rect 44324 17564 45293 17592
rect 44324 17552 44330 17564
rect 45281 17561 45293 17564
rect 45327 17561 45339 17595
rect 45281 17555 45339 17561
rect 47854 17552 47860 17604
rect 47912 17592 47918 17604
rect 48133 17595 48191 17601
rect 48133 17592 48145 17595
rect 47912 17564 48145 17592
rect 47912 17552 47918 17564
rect 48133 17561 48145 17564
rect 48179 17561 48191 17595
rect 48133 17555 48191 17561
rect 44542 17524 44548 17536
rect 44100 17496 44548 17524
rect 43441 17487 43499 17493
rect 44542 17484 44548 17496
rect 44600 17484 44606 17536
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 1946 17280 1952 17332
rect 2004 17320 2010 17332
rect 13262 17320 13268 17332
rect 2004 17292 12434 17320
rect 13223 17292 13268 17320
rect 2004 17280 2010 17292
rect 12250 17252 12256 17264
rect 11900 17224 12256 17252
rect 11900 17193 11928 17224
rect 12250 17212 12256 17224
rect 12308 17212 12314 17264
rect 11885 17187 11943 17193
rect 11885 17153 11897 17187
rect 11931 17153 11943 17187
rect 11885 17147 11943 17153
rect 11974 17144 11980 17196
rect 12032 17184 12038 17196
rect 12141 17187 12199 17193
rect 12141 17184 12153 17187
rect 12032 17156 12153 17184
rect 12032 17144 12038 17156
rect 12141 17153 12153 17156
rect 12187 17153 12199 17187
rect 12406 17184 12434 17292
rect 13262 17280 13268 17292
rect 13320 17280 13326 17332
rect 15102 17320 15108 17332
rect 15063 17292 15108 17320
rect 15102 17280 15108 17292
rect 15160 17280 15166 17332
rect 16942 17320 16948 17332
rect 16855 17292 16948 17320
rect 16942 17280 16948 17292
rect 17000 17320 17006 17332
rect 17770 17320 17776 17332
rect 17000 17292 17776 17320
rect 17000 17280 17006 17292
rect 17770 17280 17776 17292
rect 17828 17280 17834 17332
rect 18046 17280 18052 17332
rect 18104 17320 18110 17332
rect 18141 17323 18199 17329
rect 18141 17320 18153 17323
rect 18104 17292 18153 17320
rect 18104 17280 18110 17292
rect 18141 17289 18153 17292
rect 18187 17289 18199 17323
rect 18506 17320 18512 17332
rect 18467 17292 18512 17320
rect 18141 17283 18199 17289
rect 18506 17280 18512 17292
rect 18564 17280 18570 17332
rect 20254 17280 20260 17332
rect 20312 17320 20318 17332
rect 20809 17323 20867 17329
rect 20809 17320 20821 17323
rect 20312 17292 20821 17320
rect 20312 17280 20318 17292
rect 20809 17289 20821 17292
rect 20855 17289 20867 17323
rect 20809 17283 20867 17289
rect 21266 17280 21272 17332
rect 21324 17320 21330 17332
rect 22094 17320 22100 17332
rect 21324 17292 22100 17320
rect 21324 17280 21330 17292
rect 22094 17280 22100 17292
rect 22152 17280 22158 17332
rect 30098 17320 30104 17332
rect 30059 17292 30104 17320
rect 30098 17280 30104 17292
rect 30156 17280 30162 17332
rect 32490 17280 32496 17332
rect 32548 17320 32554 17332
rect 32677 17323 32735 17329
rect 32677 17320 32689 17323
rect 32548 17292 32689 17320
rect 32548 17280 32554 17292
rect 32677 17289 32689 17292
rect 32723 17320 32735 17323
rect 33042 17320 33048 17332
rect 32723 17292 33048 17320
rect 32723 17289 32735 17292
rect 32677 17283 32735 17289
rect 33042 17280 33048 17292
rect 33100 17320 33106 17332
rect 34977 17323 35035 17329
rect 33100 17292 34836 17320
rect 33100 17280 33106 17292
rect 13722 17212 13728 17264
rect 13780 17252 13786 17264
rect 14921 17255 14979 17261
rect 14921 17252 14933 17255
rect 13780 17224 14933 17252
rect 13780 17212 13786 17224
rect 14921 17221 14933 17224
rect 14967 17221 14979 17255
rect 15930 17252 15936 17264
rect 15891 17224 15936 17252
rect 14921 17215 14979 17221
rect 15930 17212 15936 17224
rect 15988 17212 15994 17264
rect 16117 17255 16175 17261
rect 16117 17221 16129 17255
rect 16163 17252 16175 17255
rect 16298 17252 16304 17264
rect 16163 17224 16304 17252
rect 16163 17221 16175 17224
rect 16117 17215 16175 17221
rect 16298 17212 16304 17224
rect 16356 17212 16362 17264
rect 17126 17252 17132 17264
rect 16408 17224 17132 17252
rect 14737 17187 14795 17193
rect 12406 17156 14688 17184
rect 12141 17147 12199 17153
rect 2038 17116 2044 17128
rect 1999 17088 2044 17116
rect 2038 17076 2044 17088
rect 2096 17076 2102 17128
rect 2225 17119 2283 17125
rect 2225 17085 2237 17119
rect 2271 17116 2283 17119
rect 2774 17116 2780 17128
rect 2271 17088 2780 17116
rect 2271 17085 2283 17088
rect 2225 17079 2283 17085
rect 2774 17076 2780 17088
rect 2832 17076 2838 17128
rect 2866 17076 2872 17128
rect 2924 17116 2930 17128
rect 14660 17116 14688 17156
rect 14737 17153 14749 17187
rect 14783 17184 14795 17187
rect 15010 17184 15016 17196
rect 14783 17156 15016 17184
rect 14783 17153 14795 17156
rect 14737 17147 14795 17153
rect 15010 17144 15016 17156
rect 15068 17184 15074 17196
rect 16408 17184 16436 17224
rect 17126 17212 17132 17224
rect 17184 17212 17190 17264
rect 19426 17252 19432 17264
rect 17880 17224 19432 17252
rect 15068 17156 16436 17184
rect 15068 17144 15074 17156
rect 16666 17144 16672 17196
rect 16724 17184 16730 17196
rect 16853 17187 16911 17193
rect 16853 17184 16865 17187
rect 16724 17156 16865 17184
rect 16724 17144 16730 17156
rect 16853 17153 16865 17156
rect 16899 17153 16911 17187
rect 17880 17184 17908 17224
rect 19426 17212 19432 17224
rect 19484 17212 19490 17264
rect 20162 17212 20168 17264
rect 20220 17252 20226 17264
rect 22002 17252 22008 17264
rect 20220 17224 22008 17252
rect 20220 17212 20226 17224
rect 18046 17184 18052 17196
rect 16853 17147 16911 17153
rect 17144 17156 17908 17184
rect 18007 17156 18052 17184
rect 17144 17116 17172 17156
rect 18046 17144 18052 17156
rect 18104 17144 18110 17196
rect 18322 17184 18328 17196
rect 18283 17156 18328 17184
rect 18322 17144 18328 17156
rect 18380 17144 18386 17196
rect 21008 17193 21036 17224
rect 22002 17212 22008 17224
rect 22060 17212 22066 17264
rect 28988 17255 29046 17261
rect 28988 17221 29000 17255
rect 29034 17252 29046 17255
rect 29178 17252 29184 17264
rect 29034 17224 29184 17252
rect 29034 17221 29046 17224
rect 28988 17215 29046 17221
rect 29178 17212 29184 17224
rect 29236 17212 29242 17264
rect 32766 17252 32772 17264
rect 32679 17224 32772 17252
rect 32766 17212 32772 17224
rect 32824 17252 32830 17264
rect 34698 17252 34704 17264
rect 32824 17224 34704 17252
rect 32824 17212 32830 17224
rect 34698 17212 34704 17224
rect 34756 17212 34762 17264
rect 34808 17252 34836 17292
rect 34977 17289 34989 17323
rect 35023 17320 35035 17323
rect 35434 17320 35440 17332
rect 35023 17292 35440 17320
rect 35023 17289 35035 17292
rect 34977 17283 35035 17289
rect 35434 17280 35440 17292
rect 35492 17280 35498 17332
rect 44266 17320 44272 17332
rect 44227 17292 44272 17320
rect 44266 17280 44272 17292
rect 44324 17280 44330 17332
rect 47854 17320 47860 17332
rect 47815 17292 47860 17320
rect 47854 17280 47860 17292
rect 47912 17280 47918 17332
rect 36446 17252 36452 17264
rect 34808 17224 36452 17252
rect 36446 17212 36452 17224
rect 36504 17212 36510 17264
rect 41064 17224 42656 17252
rect 20993 17187 21051 17193
rect 20993 17153 21005 17187
rect 21039 17153 21051 17187
rect 21266 17184 21272 17196
rect 21227 17156 21272 17184
rect 20993 17147 21051 17153
rect 21266 17144 21272 17156
rect 21324 17144 21330 17196
rect 21453 17187 21511 17193
rect 21453 17153 21465 17187
rect 21499 17184 21511 17187
rect 21542 17184 21548 17196
rect 21499 17156 21548 17184
rect 21499 17153 21511 17156
rect 21453 17147 21511 17153
rect 21542 17144 21548 17156
rect 21600 17184 21606 17196
rect 21726 17184 21732 17196
rect 21600 17156 21732 17184
rect 21600 17144 21606 17156
rect 21726 17144 21732 17156
rect 21784 17144 21790 17196
rect 23109 17187 23167 17193
rect 23109 17153 23121 17187
rect 23155 17184 23167 17187
rect 23474 17184 23480 17196
rect 23155 17156 23480 17184
rect 23155 17153 23167 17156
rect 23109 17147 23167 17153
rect 23474 17144 23480 17156
rect 23532 17144 23538 17196
rect 28534 17144 28540 17196
rect 28592 17184 28598 17196
rect 28721 17187 28779 17193
rect 28721 17184 28733 17187
rect 28592 17156 28733 17184
rect 28592 17144 28598 17156
rect 28721 17153 28733 17156
rect 28767 17153 28779 17187
rect 28721 17147 28779 17153
rect 33962 17144 33968 17196
rect 34020 17184 34026 17196
rect 34885 17187 34943 17193
rect 34885 17184 34897 17187
rect 34020 17156 34897 17184
rect 34020 17144 34026 17156
rect 34885 17153 34897 17156
rect 34931 17153 34943 17187
rect 34885 17147 34943 17153
rect 35069 17187 35127 17193
rect 35069 17153 35081 17187
rect 35115 17184 35127 17187
rect 35342 17184 35348 17196
rect 35115 17156 35348 17184
rect 35115 17153 35127 17156
rect 35069 17147 35127 17153
rect 35342 17144 35348 17156
rect 35400 17144 35406 17196
rect 40402 17144 40408 17196
rect 40460 17184 40466 17196
rect 40954 17184 40960 17196
rect 40460 17156 40960 17184
rect 40460 17144 40466 17156
rect 40954 17144 40960 17156
rect 41012 17184 41018 17196
rect 41064 17193 41092 17224
rect 41049 17187 41107 17193
rect 41049 17184 41061 17187
rect 41012 17156 41061 17184
rect 41012 17144 41018 17156
rect 41049 17153 41061 17156
rect 41095 17153 41107 17187
rect 41049 17147 41107 17153
rect 41325 17187 41383 17193
rect 41325 17153 41337 17187
rect 41371 17184 41383 17187
rect 41414 17184 41420 17196
rect 41371 17156 41420 17184
rect 41371 17153 41383 17156
rect 41325 17147 41383 17153
rect 41414 17144 41420 17156
rect 41472 17144 41478 17196
rect 42628 17193 42656 17224
rect 42613 17187 42671 17193
rect 42613 17153 42625 17187
rect 42659 17153 42671 17187
rect 42613 17147 42671 17153
rect 42978 17144 42984 17196
rect 43036 17184 43042 17196
rect 43073 17187 43131 17193
rect 43073 17184 43085 17187
rect 43036 17156 43085 17184
rect 43036 17144 43042 17156
rect 43073 17153 43085 17156
rect 43119 17153 43131 17187
rect 44450 17184 44456 17196
rect 44411 17156 44456 17184
rect 43073 17147 43131 17153
rect 44450 17144 44456 17156
rect 44508 17144 44514 17196
rect 44542 17144 44548 17196
rect 44600 17184 44606 17196
rect 44600 17156 44645 17184
rect 44600 17144 44606 17156
rect 47210 17144 47216 17196
rect 47268 17184 47274 17196
rect 47670 17184 47676 17196
rect 47268 17156 47676 17184
rect 47268 17144 47274 17156
rect 47670 17144 47676 17156
rect 47728 17184 47734 17196
rect 47765 17187 47823 17193
rect 47765 17184 47777 17187
rect 47728 17156 47777 17184
rect 47728 17144 47734 17156
rect 47765 17153 47777 17156
rect 47811 17153 47823 17187
rect 47765 17147 47823 17153
rect 2924 17088 2969 17116
rect 14660 17088 17172 17116
rect 17221 17119 17279 17125
rect 2924 17076 2930 17088
rect 17221 17085 17233 17119
rect 17267 17116 17279 17119
rect 23014 17116 23020 17128
rect 17267 17088 23020 17116
rect 17267 17085 17279 17088
rect 17221 17079 17279 17085
rect 23014 17076 23020 17088
rect 23072 17076 23078 17128
rect 23385 17119 23443 17125
rect 23385 17085 23397 17119
rect 23431 17116 23443 17119
rect 23934 17116 23940 17128
rect 23431 17088 23940 17116
rect 23431 17085 23443 17088
rect 23385 17079 23443 17085
rect 16850 17008 16856 17060
rect 16908 17048 16914 17060
rect 17129 17051 17187 17057
rect 17129 17048 17141 17051
rect 16908 17020 17141 17048
rect 16908 17008 16914 17020
rect 17129 17017 17141 17020
rect 17175 17017 17187 17051
rect 17129 17011 17187 17017
rect 18138 17008 18144 17060
rect 18196 17048 18202 17060
rect 20530 17048 20536 17060
rect 18196 17020 20536 17048
rect 18196 17008 18202 17020
rect 20530 17008 20536 17020
rect 20588 17008 20594 17060
rect 23106 17008 23112 17060
rect 23164 17048 23170 17060
rect 23400 17048 23428 17079
rect 23934 17076 23940 17088
rect 23992 17076 23998 17128
rect 42889 17119 42947 17125
rect 42889 17116 42901 17119
rect 41386 17088 42901 17116
rect 23164 17020 23428 17048
rect 41233 17051 41291 17057
rect 23164 17008 23170 17020
rect 41233 17017 41245 17051
rect 41279 17048 41291 17051
rect 41386 17048 41414 17088
rect 42889 17085 42901 17088
rect 42935 17116 42947 17119
rect 43438 17116 43444 17128
rect 42935 17088 43444 17116
rect 42935 17085 42947 17088
rect 42889 17079 42947 17085
rect 43438 17076 43444 17088
rect 43496 17076 43502 17128
rect 43714 17076 43720 17128
rect 43772 17116 43778 17128
rect 44269 17119 44327 17125
rect 44269 17116 44281 17119
rect 43772 17088 44281 17116
rect 43772 17076 43778 17088
rect 44269 17085 44281 17088
rect 44315 17116 44327 17119
rect 45278 17116 45284 17128
rect 44315 17088 45284 17116
rect 44315 17085 44327 17088
rect 44269 17079 44327 17085
rect 45278 17076 45284 17088
rect 45336 17076 45342 17128
rect 41279 17020 41414 17048
rect 41279 17017 41291 17020
rect 41233 17011 41291 17017
rect 41782 17008 41788 17060
rect 41840 17048 41846 17060
rect 42981 17051 43039 17057
rect 42981 17048 42993 17051
rect 41840 17020 42993 17048
rect 41840 17008 41846 17020
rect 42981 17017 42993 17020
rect 43027 17017 43039 17051
rect 42981 17011 43039 17017
rect 16298 16980 16304 16992
rect 16259 16952 16304 16980
rect 16298 16940 16304 16952
rect 16356 16940 16362 16992
rect 17310 16980 17316 16992
rect 17271 16952 17316 16980
rect 17310 16940 17316 16952
rect 17368 16940 17374 16992
rect 17589 16983 17647 16989
rect 17589 16949 17601 16983
rect 17635 16980 17647 16983
rect 20990 16980 20996 16992
rect 17635 16952 20996 16980
rect 17635 16949 17647 16952
rect 17589 16943 17647 16949
rect 20990 16940 20996 16952
rect 21048 16940 21054 16992
rect 23198 16980 23204 16992
rect 23159 16952 23204 16980
rect 23198 16940 23204 16952
rect 23256 16940 23262 16992
rect 23293 16983 23351 16989
rect 23293 16949 23305 16983
rect 23339 16980 23351 16983
rect 24026 16980 24032 16992
rect 23339 16952 24032 16980
rect 23339 16949 23351 16952
rect 23293 16943 23351 16949
rect 24026 16940 24032 16952
rect 24084 16940 24090 16992
rect 40126 16940 40132 16992
rect 40184 16980 40190 16992
rect 40865 16983 40923 16989
rect 40865 16980 40877 16983
rect 40184 16952 40877 16980
rect 40184 16940 40190 16952
rect 40865 16949 40877 16952
rect 40911 16949 40923 16983
rect 40865 16943 40923 16949
rect 41414 16940 41420 16992
rect 41472 16980 41478 16992
rect 42751 16983 42809 16989
rect 42751 16980 42763 16983
rect 41472 16952 42763 16980
rect 41472 16940 41478 16952
rect 42751 16949 42763 16952
rect 42797 16980 42809 16983
rect 43346 16980 43352 16992
rect 42797 16952 43352 16980
rect 42797 16949 42809 16952
rect 42751 16943 42809 16949
rect 43346 16940 43352 16952
rect 43404 16940 43410 16992
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 2038 16736 2044 16788
rect 2096 16776 2102 16788
rect 2133 16779 2191 16785
rect 2133 16776 2145 16779
rect 2096 16748 2145 16776
rect 2096 16736 2102 16748
rect 2133 16745 2145 16748
rect 2179 16745 2191 16779
rect 2133 16739 2191 16745
rect 16025 16779 16083 16785
rect 16025 16745 16037 16779
rect 16071 16776 16083 16779
rect 17310 16776 17316 16788
rect 16071 16748 17316 16776
rect 16071 16745 16083 16748
rect 16025 16739 16083 16745
rect 17310 16736 17316 16748
rect 17368 16736 17374 16788
rect 20622 16736 20628 16788
rect 20680 16776 20686 16788
rect 20680 16748 20852 16776
rect 20680 16736 20686 16748
rect 16853 16711 16911 16717
rect 16853 16677 16865 16711
rect 16899 16708 16911 16711
rect 18046 16708 18052 16720
rect 16899 16680 18052 16708
rect 16899 16677 16911 16680
rect 16853 16671 16911 16677
rect 18046 16668 18052 16680
rect 18104 16668 18110 16720
rect 13722 16600 13728 16652
rect 13780 16640 13786 16652
rect 13780 16612 14780 16640
rect 13780 16600 13786 16612
rect 2774 16532 2780 16584
rect 2832 16572 2838 16584
rect 2869 16575 2927 16581
rect 2869 16572 2881 16575
rect 2832 16544 2881 16572
rect 2832 16532 2838 16544
rect 2869 16541 2881 16544
rect 2915 16541 2927 16575
rect 2869 16535 2927 16541
rect 2958 16532 2964 16584
rect 3016 16572 3022 16584
rect 14752 16581 14780 16612
rect 16022 16600 16028 16652
rect 16080 16640 16086 16652
rect 16298 16640 16304 16652
rect 16080 16612 16304 16640
rect 16080 16600 16086 16612
rect 16298 16600 16304 16612
rect 16356 16640 16362 16652
rect 16485 16643 16543 16649
rect 16485 16640 16497 16643
rect 16356 16612 16497 16640
rect 16356 16600 16362 16612
rect 16485 16609 16497 16612
rect 16531 16609 16543 16643
rect 16485 16603 16543 16609
rect 16574 16600 16580 16652
rect 16632 16640 16638 16652
rect 20824 16649 20852 16748
rect 21560 16748 21772 16776
rect 20809 16643 20867 16649
rect 16632 16612 16712 16640
rect 16632 16600 16638 16612
rect 14737 16575 14795 16581
rect 3016 16544 3061 16572
rect 3016 16532 3022 16544
rect 14737 16541 14749 16575
rect 14783 16541 14795 16575
rect 14737 16535 14795 16541
rect 14921 16575 14979 16581
rect 14921 16541 14933 16575
rect 14967 16572 14979 16575
rect 15010 16572 15016 16584
rect 14967 16544 15016 16572
rect 14967 16541 14979 16544
rect 14921 16535 14979 16541
rect 15010 16532 15016 16544
rect 15068 16532 15074 16584
rect 15657 16575 15715 16581
rect 15657 16541 15669 16575
rect 15703 16572 15715 16575
rect 15930 16572 15936 16584
rect 15703 16544 15936 16572
rect 15703 16541 15715 16544
rect 15657 16535 15715 16541
rect 15930 16532 15936 16544
rect 15988 16532 15994 16584
rect 16684 16581 16712 16612
rect 20809 16609 20821 16643
rect 20855 16609 20867 16643
rect 20809 16603 20867 16609
rect 16669 16575 16727 16581
rect 16669 16541 16681 16575
rect 16715 16541 16727 16575
rect 21453 16575 21511 16581
rect 16669 16535 16727 16541
rect 20088 16544 21404 16572
rect 15838 16504 15844 16516
rect 15799 16476 15844 16504
rect 15838 16464 15844 16476
rect 15896 16464 15902 16516
rect 20088 16448 20116 16544
rect 20254 16464 20260 16516
rect 20312 16504 20318 16516
rect 20542 16507 20600 16513
rect 20542 16504 20554 16507
rect 20312 16476 20554 16504
rect 20312 16464 20318 16476
rect 20542 16473 20554 16476
rect 20588 16473 20600 16507
rect 20542 16467 20600 16473
rect 14829 16439 14887 16445
rect 14829 16405 14841 16439
rect 14875 16436 14887 16439
rect 15194 16436 15200 16448
rect 14875 16408 15200 16436
rect 14875 16405 14887 16408
rect 14829 16399 14887 16405
rect 15194 16396 15200 16408
rect 15252 16396 15258 16448
rect 19429 16439 19487 16445
rect 19429 16405 19441 16439
rect 19475 16436 19487 16439
rect 20070 16436 20076 16448
rect 19475 16408 20076 16436
rect 19475 16405 19487 16408
rect 19429 16399 19487 16405
rect 20070 16396 20076 16408
rect 20128 16396 20134 16448
rect 20438 16396 20444 16448
rect 20496 16436 20502 16448
rect 21269 16439 21327 16445
rect 21269 16436 21281 16439
rect 20496 16408 21281 16436
rect 20496 16396 20502 16408
rect 21269 16405 21281 16408
rect 21315 16405 21327 16439
rect 21376 16436 21404 16544
rect 21453 16541 21465 16575
rect 21499 16572 21511 16575
rect 21560 16572 21588 16748
rect 21744 16640 21772 16748
rect 23014 16736 23020 16788
rect 23072 16776 23078 16788
rect 23109 16779 23167 16785
rect 23109 16776 23121 16779
rect 23072 16748 23121 16776
rect 23072 16736 23078 16748
rect 23109 16745 23121 16748
rect 23155 16776 23167 16779
rect 23382 16776 23388 16788
rect 23155 16748 23388 16776
rect 23155 16745 23167 16748
rect 23109 16739 23167 16745
rect 23382 16736 23388 16748
rect 23440 16736 23446 16788
rect 30377 16779 30435 16785
rect 30377 16745 30389 16779
rect 30423 16776 30435 16779
rect 31110 16776 31116 16788
rect 30423 16748 31116 16776
rect 30423 16745 30435 16748
rect 30377 16739 30435 16745
rect 31110 16736 31116 16748
rect 31168 16736 31174 16788
rect 37550 16736 37556 16788
rect 37608 16736 37614 16788
rect 40218 16776 40224 16788
rect 38120 16748 40224 16776
rect 37568 16708 37596 16736
rect 36280 16680 37596 16708
rect 21744 16612 21956 16640
rect 21499 16544 21588 16572
rect 21499 16541 21511 16544
rect 21453 16535 21511 16541
rect 21634 16532 21640 16584
rect 21692 16572 21698 16584
rect 21821 16575 21879 16581
rect 21692 16544 21737 16572
rect 21692 16532 21698 16544
rect 21821 16541 21833 16575
rect 21867 16541 21879 16575
rect 21928 16572 21956 16612
rect 23308 16612 23612 16640
rect 23308 16572 23336 16612
rect 23474 16572 23480 16584
rect 21928 16544 23336 16572
rect 23435 16544 23480 16572
rect 21821 16535 21879 16541
rect 21542 16504 21548 16516
rect 21503 16476 21548 16504
rect 21542 16464 21548 16476
rect 21600 16464 21606 16516
rect 21836 16436 21864 16535
rect 23474 16532 23480 16544
rect 23532 16532 23538 16584
rect 23584 16572 23612 16612
rect 24854 16600 24860 16652
rect 24912 16640 24918 16652
rect 24912 16612 25452 16640
rect 24912 16600 24918 16612
rect 25222 16572 25228 16584
rect 23584 16544 25228 16572
rect 25222 16532 25228 16544
rect 25280 16532 25286 16584
rect 25424 16581 25452 16612
rect 25409 16575 25467 16581
rect 25409 16541 25421 16575
rect 25455 16541 25467 16575
rect 25590 16572 25596 16584
rect 25551 16544 25596 16572
rect 25409 16535 25467 16541
rect 25590 16532 25596 16544
rect 25648 16532 25654 16584
rect 29454 16532 29460 16584
rect 29512 16572 29518 16584
rect 29733 16575 29791 16581
rect 29733 16572 29745 16575
rect 29512 16544 29745 16572
rect 29512 16532 29518 16544
rect 29733 16541 29745 16544
rect 29779 16541 29791 16575
rect 29733 16535 29791 16541
rect 29917 16575 29975 16581
rect 29917 16541 29929 16575
rect 29963 16541 29975 16575
rect 29917 16535 29975 16541
rect 30193 16575 30251 16581
rect 30193 16541 30205 16575
rect 30239 16572 30251 16575
rect 30742 16572 30748 16584
rect 30239 16544 30748 16572
rect 30239 16541 30251 16544
rect 30193 16535 30251 16541
rect 23290 16504 23296 16516
rect 23251 16476 23296 16504
rect 23290 16464 23296 16476
rect 23348 16464 23354 16516
rect 25317 16507 25375 16513
rect 25317 16473 25329 16507
rect 25363 16473 25375 16507
rect 29932 16504 29960 16535
rect 30742 16532 30748 16544
rect 30800 16532 30806 16584
rect 36078 16572 36084 16584
rect 36039 16544 36084 16572
rect 36078 16532 36084 16544
rect 36136 16532 36142 16584
rect 36280 16581 36308 16680
rect 37274 16600 37280 16652
rect 37332 16640 37338 16652
rect 38120 16649 38148 16748
rect 40218 16736 40224 16748
rect 40276 16736 40282 16788
rect 43438 16776 43444 16788
rect 43399 16748 43444 16776
rect 43438 16736 43444 16748
rect 43496 16736 43502 16788
rect 45281 16779 45339 16785
rect 45281 16745 45293 16779
rect 45327 16776 45339 16779
rect 45462 16776 45468 16788
rect 45327 16748 45468 16776
rect 45327 16745 45339 16748
rect 45281 16739 45339 16745
rect 45462 16736 45468 16748
rect 45520 16736 45526 16788
rect 37553 16643 37611 16649
rect 37553 16640 37565 16643
rect 37332 16612 37565 16640
rect 37332 16600 37338 16612
rect 37553 16609 37565 16612
rect 37599 16640 37611 16643
rect 38105 16643 38163 16649
rect 38105 16640 38117 16643
rect 37599 16612 38117 16640
rect 37599 16609 37611 16612
rect 37553 16603 37611 16609
rect 38105 16609 38117 16612
rect 38151 16609 38163 16643
rect 38105 16603 38163 16609
rect 40034 16600 40040 16652
rect 40092 16640 40098 16652
rect 40681 16643 40739 16649
rect 40681 16640 40693 16643
rect 40092 16612 40693 16640
rect 40092 16600 40098 16612
rect 40681 16609 40693 16612
rect 40727 16609 40739 16643
rect 40681 16603 40739 16609
rect 41506 16600 41512 16652
rect 41564 16640 41570 16652
rect 42334 16640 42340 16652
rect 41564 16612 41920 16640
rect 41564 16600 41570 16612
rect 36265 16575 36323 16581
rect 36265 16541 36277 16575
rect 36311 16541 36323 16575
rect 36265 16535 36323 16541
rect 40126 16532 40132 16584
rect 40184 16572 40190 16584
rect 40221 16575 40279 16581
rect 40221 16572 40233 16575
rect 40184 16544 40233 16572
rect 40184 16532 40190 16544
rect 40221 16541 40233 16544
rect 40267 16541 40279 16575
rect 40221 16535 40279 16541
rect 40313 16575 40371 16581
rect 40313 16541 40325 16575
rect 40359 16572 40371 16575
rect 41782 16572 41788 16584
rect 40359 16544 41788 16572
rect 40359 16541 40371 16544
rect 40313 16535 40371 16541
rect 41782 16532 41788 16544
rect 41840 16532 41846 16584
rect 41892 16581 41920 16612
rect 42168 16612 42340 16640
rect 42168 16581 42196 16612
rect 42334 16600 42340 16612
rect 42392 16600 42398 16652
rect 42981 16643 43039 16649
rect 42981 16609 42993 16643
rect 43027 16609 43039 16643
rect 46106 16640 46112 16652
rect 46067 16612 46112 16640
rect 42981 16603 43039 16609
rect 41877 16575 41935 16581
rect 41877 16541 41889 16575
rect 41923 16541 41935 16575
rect 41877 16535 41935 16541
rect 42061 16575 42119 16581
rect 42061 16541 42073 16575
rect 42107 16541 42119 16575
rect 42061 16535 42119 16541
rect 42153 16575 42211 16581
rect 42153 16541 42165 16575
rect 42199 16541 42211 16575
rect 42153 16535 42211 16541
rect 30558 16504 30564 16516
rect 29932 16476 30564 16504
rect 25317 16467 25375 16473
rect 21376 16408 21864 16436
rect 25041 16439 25099 16445
rect 21269 16399 21327 16405
rect 25041 16405 25053 16439
rect 25087 16436 25099 16439
rect 25222 16436 25228 16448
rect 25087 16408 25228 16436
rect 25087 16405 25099 16408
rect 25041 16399 25099 16405
rect 25222 16396 25228 16408
rect 25280 16396 25286 16448
rect 25332 16436 25360 16467
rect 30558 16464 30564 16476
rect 30616 16464 30622 16516
rect 31754 16464 31760 16516
rect 31812 16504 31818 16516
rect 36725 16507 36783 16513
rect 36725 16504 36737 16507
rect 31812 16476 36737 16504
rect 31812 16464 31818 16476
rect 36725 16473 36737 16476
rect 36771 16473 36783 16507
rect 36725 16467 36783 16473
rect 38372 16507 38430 16513
rect 38372 16473 38384 16507
rect 38418 16504 38430 16507
rect 40589 16507 40647 16513
rect 38418 16476 40080 16504
rect 38418 16473 38430 16476
rect 38372 16467 38430 16473
rect 27798 16436 27804 16448
rect 25332 16408 27804 16436
rect 27798 16396 27804 16408
rect 27856 16396 27862 16448
rect 34146 16396 34152 16448
rect 34204 16436 34210 16448
rect 36170 16436 36176 16448
rect 34204 16408 36176 16436
rect 34204 16396 34210 16408
rect 36170 16396 36176 16408
rect 36228 16396 36234 16448
rect 36265 16439 36323 16445
rect 36265 16405 36277 16439
rect 36311 16436 36323 16439
rect 36446 16436 36452 16448
rect 36311 16408 36452 16436
rect 36311 16405 36323 16408
rect 36265 16399 36323 16405
rect 36446 16396 36452 16408
rect 36504 16396 36510 16448
rect 39485 16439 39543 16445
rect 39485 16405 39497 16439
rect 39531 16436 39543 16439
rect 39942 16436 39948 16448
rect 39531 16408 39948 16436
rect 39531 16405 39543 16408
rect 39485 16399 39543 16405
rect 39942 16396 39948 16408
rect 40000 16396 40006 16448
rect 40052 16445 40080 16476
rect 40589 16473 40601 16507
rect 40635 16504 40647 16507
rect 40678 16504 40684 16516
rect 40635 16476 40684 16504
rect 40635 16473 40647 16476
rect 40589 16467 40647 16473
rect 40678 16464 40684 16476
rect 40736 16464 40742 16516
rect 42076 16504 42104 16535
rect 42242 16532 42248 16584
rect 42300 16572 42306 16584
rect 42996 16572 43024 16603
rect 46106 16600 46112 16612
rect 46164 16600 46170 16652
rect 42300 16544 43024 16572
rect 42300 16532 42306 16544
rect 43070 16532 43076 16584
rect 43128 16572 43134 16584
rect 43128 16544 43173 16572
rect 43128 16532 43134 16544
rect 43254 16532 43260 16584
rect 43312 16572 43318 16584
rect 45186 16572 45192 16584
rect 43312 16544 43357 16572
rect 45147 16544 45192 16572
rect 43312 16532 43318 16544
rect 45186 16532 45192 16544
rect 45244 16532 45250 16584
rect 45373 16575 45431 16581
rect 45373 16541 45385 16575
rect 45419 16572 45431 16575
rect 45462 16572 45468 16584
rect 45419 16544 45468 16572
rect 45419 16541 45431 16544
rect 45373 16535 45431 16541
rect 45462 16532 45468 16544
rect 45520 16532 45526 16584
rect 43272 16504 43300 16532
rect 42076 16476 43300 16504
rect 46376 16507 46434 16513
rect 46376 16473 46388 16507
rect 46422 16504 46434 16507
rect 46658 16504 46664 16516
rect 46422 16476 46664 16504
rect 46422 16473 46434 16476
rect 46376 16467 46434 16473
rect 46658 16464 46664 16476
rect 46716 16464 46722 16516
rect 40037 16439 40095 16445
rect 40037 16405 40049 16439
rect 40083 16405 40095 16439
rect 40037 16399 40095 16405
rect 42521 16439 42579 16445
rect 42521 16405 42533 16439
rect 42567 16436 42579 16439
rect 42794 16436 42800 16448
rect 42567 16408 42800 16436
rect 42567 16405 42579 16408
rect 42521 16399 42579 16405
rect 42794 16396 42800 16408
rect 42852 16396 42858 16448
rect 47394 16396 47400 16448
rect 47452 16436 47458 16448
rect 47489 16439 47547 16445
rect 47489 16436 47501 16439
rect 47452 16408 47501 16436
rect 47452 16396 47458 16408
rect 47489 16405 47501 16408
rect 47535 16405 47547 16439
rect 47489 16399 47547 16405
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 16298 16192 16304 16244
rect 16356 16232 16362 16244
rect 20254 16232 20260 16244
rect 16356 16204 17080 16232
rect 20215 16204 20260 16232
rect 16356 16192 16362 16204
rect 15194 16164 15200 16176
rect 14568 16136 15200 16164
rect 14568 16105 14596 16136
rect 15194 16124 15200 16136
rect 15252 16164 15258 16176
rect 15252 16136 16252 16164
rect 15252 16124 15258 16136
rect 14553 16099 14611 16105
rect 14553 16065 14565 16099
rect 14599 16065 14611 16099
rect 14553 16059 14611 16065
rect 14642 16056 14648 16108
rect 14700 16096 14706 16108
rect 14700 16068 14745 16096
rect 14700 16056 14706 16068
rect 14826 16056 14832 16108
rect 14884 16096 14890 16108
rect 15933 16099 15991 16105
rect 14884 16068 14929 16096
rect 14884 16056 14890 16068
rect 15933 16065 15945 16099
rect 15979 16096 15991 16099
rect 16022 16096 16028 16108
rect 15979 16068 16028 16096
rect 15979 16065 15991 16068
rect 15933 16059 15991 16065
rect 16022 16056 16028 16068
rect 16080 16056 16086 16108
rect 16117 16099 16175 16105
rect 16117 16065 16129 16099
rect 16163 16065 16175 16099
rect 16224 16096 16252 16136
rect 17052 16105 17080 16204
rect 20254 16192 20260 16204
rect 20312 16192 20318 16244
rect 20530 16192 20536 16244
rect 20588 16232 20594 16244
rect 20625 16235 20683 16241
rect 20625 16232 20637 16235
rect 20588 16204 20637 16232
rect 20588 16192 20594 16204
rect 20625 16201 20637 16204
rect 20671 16232 20683 16235
rect 24489 16235 24547 16241
rect 20671 16204 22094 16232
rect 20671 16201 20683 16204
rect 20625 16195 20683 16201
rect 22066 16164 22094 16204
rect 24489 16201 24501 16235
rect 24535 16201 24547 16235
rect 24489 16195 24547 16201
rect 22066 16136 24256 16164
rect 16853 16099 16911 16105
rect 16853 16096 16865 16099
rect 16224 16068 16865 16096
rect 16117 16059 16175 16065
rect 16853 16065 16865 16068
rect 16899 16065 16911 16099
rect 16853 16059 16911 16065
rect 17037 16099 17095 16105
rect 17037 16065 17049 16099
rect 17083 16065 17095 16099
rect 20438 16096 20444 16108
rect 20399 16068 20444 16096
rect 17037 16059 17095 16065
rect 15838 16028 15844 16040
rect 15799 16000 15844 16028
rect 15838 15988 15844 16000
rect 15896 15988 15902 16040
rect 16132 16028 16160 16059
rect 20438 16056 20444 16068
rect 20496 16056 20502 16108
rect 20717 16099 20775 16105
rect 20717 16065 20729 16099
rect 20763 16096 20775 16099
rect 21450 16096 21456 16108
rect 20763 16068 21456 16096
rect 20763 16065 20775 16068
rect 20717 16059 20775 16065
rect 21450 16056 21456 16068
rect 21508 16056 21514 16108
rect 22830 16056 22836 16108
rect 22888 16096 22894 16108
rect 22925 16099 22983 16105
rect 22925 16096 22937 16099
rect 22888 16068 22937 16096
rect 22888 16056 22894 16068
rect 22925 16065 22937 16068
rect 22971 16065 22983 16099
rect 23201 16099 23259 16105
rect 23201 16096 23213 16099
rect 22925 16059 22983 16065
rect 23032 16068 23213 16096
rect 23032 16028 23060 16068
rect 23201 16065 23213 16068
rect 23247 16065 23259 16099
rect 23201 16059 23259 16065
rect 23293 16099 23351 16105
rect 23293 16065 23305 16099
rect 23339 16096 23351 16099
rect 23382 16096 23388 16108
rect 23339 16068 23388 16096
rect 23339 16065 23351 16068
rect 23293 16059 23351 16065
rect 23382 16056 23388 16068
rect 23440 16056 23446 16108
rect 23474 16056 23480 16108
rect 23532 16096 23538 16108
rect 24121 16099 24179 16105
rect 23532 16068 23577 16096
rect 23532 16056 23538 16068
rect 24121 16065 24133 16099
rect 24167 16065 24179 16099
rect 24121 16059 24179 16065
rect 16132 16000 23060 16028
rect 15013 15963 15071 15969
rect 15013 15929 15025 15963
rect 15059 15960 15071 15963
rect 16132 15960 16160 16000
rect 23106 15988 23112 16040
rect 23164 16028 23170 16040
rect 24026 16028 24032 16040
rect 23164 16000 23209 16028
rect 23987 16000 24032 16028
rect 23164 15988 23170 16000
rect 24026 15988 24032 16000
rect 24084 15988 24090 16040
rect 15059 15932 16160 15960
rect 16301 15963 16359 15969
rect 15059 15929 15071 15932
rect 15013 15923 15071 15929
rect 16301 15929 16313 15963
rect 16347 15960 16359 15963
rect 23198 15960 23204 15972
rect 16347 15932 23204 15960
rect 16347 15929 16359 15932
rect 16301 15923 16359 15929
rect 23198 15920 23204 15932
rect 23256 15920 23262 15972
rect 23290 15920 23296 15972
rect 23348 15960 23354 15972
rect 24136 15960 24164 16059
rect 24228 16028 24256 16136
rect 24504 16096 24532 16195
rect 26510 16192 26516 16244
rect 26568 16232 26574 16244
rect 28626 16232 28632 16244
rect 26568 16204 28632 16232
rect 26568 16192 26574 16204
rect 28626 16192 28632 16204
rect 28684 16192 28690 16244
rect 36078 16192 36084 16244
rect 36136 16232 36142 16244
rect 36136 16204 37504 16232
rect 36136 16192 36142 16204
rect 27706 16164 27712 16176
rect 27356 16136 27712 16164
rect 27356 16108 27384 16136
rect 27706 16124 27712 16136
rect 27764 16124 27770 16176
rect 28718 16164 28724 16176
rect 28368 16136 28724 16164
rect 24949 16099 25007 16105
rect 24949 16096 24961 16099
rect 24504 16068 24961 16096
rect 24949 16065 24961 16068
rect 24995 16065 25007 16099
rect 24949 16059 25007 16065
rect 25041 16099 25099 16105
rect 25041 16065 25053 16099
rect 25087 16065 25099 16099
rect 25222 16096 25228 16108
rect 25183 16068 25228 16096
rect 25041 16059 25099 16065
rect 25056 16028 25084 16059
rect 25222 16056 25228 16068
rect 25280 16056 25286 16108
rect 26329 16099 26387 16105
rect 26329 16065 26341 16099
rect 26375 16096 26387 16099
rect 27157 16099 27215 16105
rect 27157 16096 27169 16099
rect 26375 16068 27169 16096
rect 26375 16065 26387 16068
rect 26329 16059 26387 16065
rect 27157 16065 27169 16068
rect 27203 16065 27215 16099
rect 27157 16059 27215 16065
rect 27338 16056 27344 16108
rect 27396 16096 27402 16108
rect 27614 16096 27620 16108
rect 27396 16068 27489 16096
rect 27575 16068 27620 16096
rect 27396 16056 27402 16068
rect 27614 16056 27620 16068
rect 27672 16056 27678 16108
rect 27798 16096 27804 16108
rect 27759 16068 27804 16096
rect 27798 16056 27804 16068
rect 27856 16056 27862 16108
rect 28368 16105 28396 16136
rect 28718 16124 28724 16136
rect 28776 16164 28782 16176
rect 30929 16167 30987 16173
rect 30929 16164 30941 16167
rect 28776 16136 30941 16164
rect 28776 16124 28782 16136
rect 30929 16133 30941 16136
rect 30975 16133 30987 16167
rect 30929 16127 30987 16133
rect 31754 16124 31760 16176
rect 31812 16164 31818 16176
rect 37274 16164 37280 16176
rect 31812 16136 31857 16164
rect 32324 16136 37280 16164
rect 31812 16124 31818 16136
rect 32324 16108 32352 16136
rect 28626 16105 28632 16108
rect 28353 16099 28411 16105
rect 28353 16065 28365 16099
rect 28399 16065 28411 16099
rect 28353 16059 28411 16065
rect 28620 16059 28632 16105
rect 28684 16096 28690 16108
rect 32306 16096 32312 16108
rect 28684 16068 28720 16096
rect 32219 16068 32312 16096
rect 28626 16056 28632 16059
rect 28684 16056 28690 16068
rect 32306 16056 32312 16068
rect 32364 16056 32370 16108
rect 32398 16056 32404 16108
rect 32456 16096 32462 16108
rect 34164 16105 34192 16136
rect 37274 16124 37280 16136
rect 37332 16124 37338 16176
rect 32565 16099 32623 16105
rect 32565 16096 32577 16099
rect 32456 16068 32577 16096
rect 32456 16056 32462 16068
rect 32565 16065 32577 16068
rect 32611 16065 32623 16099
rect 32565 16059 32623 16065
rect 34149 16099 34207 16105
rect 34149 16065 34161 16099
rect 34195 16065 34207 16099
rect 34149 16059 34207 16065
rect 34238 16056 34244 16108
rect 34296 16096 34302 16108
rect 34405 16099 34463 16105
rect 34405 16096 34417 16099
rect 34296 16068 34417 16096
rect 34296 16056 34302 16068
rect 34405 16065 34417 16068
rect 34451 16065 34463 16099
rect 34405 16059 34463 16065
rect 35989 16099 36047 16105
rect 35989 16065 36001 16099
rect 36035 16065 36047 16099
rect 36170 16096 36176 16108
rect 36131 16068 36176 16096
rect 35989 16059 36047 16065
rect 26510 16028 26516 16040
rect 24228 16000 25084 16028
rect 26471 16000 26516 16028
rect 26510 15988 26516 16000
rect 26568 15988 26574 16040
rect 26605 16031 26663 16037
rect 26605 15997 26617 16031
rect 26651 15997 26663 16031
rect 36004 16028 36032 16059
rect 36170 16056 36176 16068
rect 36228 16056 36234 16108
rect 37476 16105 37504 16204
rect 37550 16192 37556 16244
rect 37608 16232 37614 16244
rect 37608 16204 37653 16232
rect 37608 16192 37614 16204
rect 40310 16192 40316 16244
rect 40368 16232 40374 16244
rect 41325 16235 41383 16241
rect 41325 16232 41337 16235
rect 40368 16204 41337 16232
rect 40368 16192 40374 16204
rect 41325 16201 41337 16204
rect 41371 16201 41383 16235
rect 41325 16195 41383 16201
rect 42334 16192 42340 16244
rect 42392 16232 42398 16244
rect 43070 16232 43076 16244
rect 42392 16204 43076 16232
rect 42392 16192 42398 16204
rect 43070 16192 43076 16204
rect 43128 16192 43134 16244
rect 45278 16232 45284 16244
rect 43640 16204 45284 16232
rect 41046 16164 41052 16176
rect 40052 16136 41052 16164
rect 37461 16099 37519 16105
rect 37461 16065 37473 16099
rect 37507 16065 37519 16099
rect 37734 16096 37740 16108
rect 37695 16068 37740 16096
rect 37461 16059 37519 16065
rect 37734 16056 37740 16068
rect 37792 16056 37798 16108
rect 40052 16105 40080 16136
rect 40328 16108 40356 16136
rect 41046 16124 41052 16136
rect 41104 16164 41110 16176
rect 43640 16164 43668 16204
rect 45278 16192 45284 16204
rect 45336 16192 45342 16244
rect 45649 16235 45707 16241
rect 45649 16201 45661 16235
rect 45695 16201 45707 16235
rect 46658 16232 46664 16244
rect 46619 16204 46664 16232
rect 45649 16195 45707 16201
rect 41104 16136 43668 16164
rect 41104 16124 41110 16136
rect 40037 16099 40095 16105
rect 40037 16065 40049 16099
rect 40083 16065 40095 16099
rect 40037 16059 40095 16065
rect 40310 16056 40316 16108
rect 40368 16056 40374 16108
rect 41156 16105 41184 16136
rect 44450 16124 44456 16176
rect 44508 16164 44514 16176
rect 45664 16164 45692 16195
rect 46658 16192 46664 16204
rect 46716 16192 46722 16244
rect 46293 16167 46351 16173
rect 46293 16164 46305 16167
rect 44508 16136 45416 16164
rect 45664 16136 46305 16164
rect 44508 16124 44514 16136
rect 41141 16099 41199 16105
rect 41141 16065 41153 16099
rect 41187 16096 41199 16099
rect 41187 16068 41221 16096
rect 41187 16065 41199 16068
rect 41141 16059 41199 16065
rect 42886 16056 42892 16108
rect 42944 16096 42950 16108
rect 44269 16099 44327 16105
rect 44269 16096 44281 16099
rect 42944 16068 44281 16096
rect 42944 16056 42950 16068
rect 44269 16065 44281 16068
rect 44315 16065 44327 16099
rect 45186 16096 45192 16108
rect 44269 16059 44327 16065
rect 44652 16068 45192 16096
rect 39942 16028 39948 16040
rect 26605 15991 26663 15997
rect 35544 16000 36032 16028
rect 39903 16000 39948 16028
rect 23348 15932 24164 15960
rect 23348 15920 23354 15932
rect 26620 15904 26648 15991
rect 16942 15892 16948 15904
rect 16903 15864 16948 15892
rect 16942 15852 16948 15864
rect 17000 15852 17006 15904
rect 20806 15852 20812 15904
rect 20864 15892 20870 15904
rect 22741 15895 22799 15901
rect 22741 15892 22753 15895
rect 20864 15864 22753 15892
rect 20864 15852 20870 15864
rect 22741 15861 22753 15864
rect 22787 15861 22799 15895
rect 25406 15892 25412 15904
rect 25367 15864 25412 15892
rect 22741 15855 22799 15861
rect 25406 15852 25412 15864
rect 25464 15852 25470 15904
rect 26142 15892 26148 15904
rect 26103 15864 26148 15892
rect 26142 15852 26148 15864
rect 26200 15852 26206 15904
rect 26602 15852 26608 15904
rect 26660 15892 26666 15904
rect 29454 15892 29460 15904
rect 26660 15864 29460 15892
rect 26660 15852 26666 15864
rect 29454 15852 29460 15864
rect 29512 15852 29518 15904
rect 29733 15895 29791 15901
rect 29733 15861 29745 15895
rect 29779 15892 29791 15895
rect 30834 15892 30840 15904
rect 29779 15864 30840 15892
rect 29779 15861 29791 15864
rect 29733 15855 29791 15861
rect 30834 15852 30840 15864
rect 30892 15852 30898 15904
rect 31754 15852 31760 15904
rect 31812 15892 31818 15904
rect 33686 15892 33692 15904
rect 31812 15864 33692 15892
rect 31812 15852 31818 15864
rect 33686 15852 33692 15864
rect 33744 15852 33750 15904
rect 35434 15852 35440 15904
rect 35492 15892 35498 15904
rect 35544 15901 35572 16000
rect 39942 15988 39948 16000
rect 40000 16028 40006 16040
rect 40865 16031 40923 16037
rect 40865 16028 40877 16031
rect 40000 16000 40877 16028
rect 40000 15988 40006 16000
rect 40865 15997 40877 16000
rect 40911 15997 40923 16031
rect 40865 15991 40923 15997
rect 44361 16031 44419 16037
rect 44361 15997 44373 16031
rect 44407 16028 44419 16031
rect 44450 16028 44456 16040
rect 44407 16000 44456 16028
rect 44407 15997 44419 16000
rect 44361 15991 44419 15997
rect 44450 15988 44456 16000
rect 44508 15988 44514 16040
rect 37737 15963 37795 15969
rect 37737 15929 37749 15963
rect 37783 15960 37795 15963
rect 42242 15960 42248 15972
rect 37783 15932 42248 15960
rect 37783 15929 37795 15932
rect 37737 15923 37795 15929
rect 42242 15920 42248 15932
rect 42300 15920 42306 15972
rect 44652 15904 44680 16068
rect 45186 16056 45192 16068
rect 45244 16096 45250 16108
rect 45281 16099 45339 16105
rect 45281 16096 45293 16099
rect 45244 16068 45293 16096
rect 45244 16056 45250 16068
rect 45281 16065 45293 16068
rect 45327 16065 45339 16099
rect 45388 16096 45416 16136
rect 46293 16133 46305 16136
rect 46339 16133 46351 16167
rect 47394 16164 47400 16176
rect 46293 16127 46351 16133
rect 46400 16136 47400 16164
rect 45388 16068 45508 16096
rect 45281 16059 45339 16065
rect 45370 16028 45376 16040
rect 45331 16000 45376 16028
rect 45370 15988 45376 16000
rect 45428 15988 45434 16040
rect 45480 15960 45508 16068
rect 45554 16056 45560 16108
rect 45612 16096 45618 16108
rect 46400 16105 46428 16136
rect 47394 16124 47400 16136
rect 47452 16124 47458 16176
rect 46109 16099 46167 16105
rect 46109 16096 46121 16099
rect 45612 16068 46121 16096
rect 45612 16056 45618 16068
rect 46109 16065 46121 16068
rect 46155 16065 46167 16099
rect 46109 16059 46167 16065
rect 46385 16099 46443 16105
rect 46385 16065 46397 16099
rect 46431 16065 46443 16099
rect 46385 16059 46443 16065
rect 46400 15960 46428 16059
rect 46474 16056 46480 16108
rect 46532 16096 46538 16108
rect 46532 16068 46577 16096
rect 46532 16056 46538 16068
rect 45480 15932 46428 15960
rect 35529 15895 35587 15901
rect 35529 15892 35541 15895
rect 35492 15864 35541 15892
rect 35492 15852 35498 15864
rect 35529 15861 35541 15864
rect 35575 15861 35587 15895
rect 36354 15892 36360 15904
rect 36315 15864 36360 15892
rect 35529 15855 35587 15861
rect 36354 15852 36360 15864
rect 36412 15852 36418 15904
rect 40402 15892 40408 15904
rect 40363 15864 40408 15892
rect 40402 15852 40408 15864
rect 40460 15852 40466 15904
rect 40954 15892 40960 15904
rect 40915 15864 40960 15892
rect 40954 15852 40960 15864
rect 41012 15852 41018 15904
rect 44634 15892 44640 15904
rect 44595 15864 44640 15892
rect 44634 15852 44640 15864
rect 44692 15852 44698 15904
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 14274 15648 14280 15700
rect 14332 15688 14338 15700
rect 14645 15691 14703 15697
rect 14645 15688 14657 15691
rect 14332 15660 14657 15688
rect 14332 15648 14338 15660
rect 14645 15657 14657 15660
rect 14691 15688 14703 15691
rect 14826 15688 14832 15700
rect 14691 15660 14832 15688
rect 14691 15657 14703 15660
rect 14645 15651 14703 15657
rect 14826 15648 14832 15660
rect 14884 15648 14890 15700
rect 21450 15688 21456 15700
rect 21411 15660 21456 15688
rect 21450 15648 21456 15660
rect 21508 15648 21514 15700
rect 23290 15688 23296 15700
rect 23251 15660 23296 15688
rect 23290 15648 23296 15660
rect 23348 15648 23354 15700
rect 23661 15691 23719 15697
rect 23661 15657 23673 15691
rect 23707 15688 23719 15691
rect 24581 15691 24639 15697
rect 24581 15688 24593 15691
rect 23707 15660 24593 15688
rect 23707 15657 23719 15660
rect 23661 15651 23719 15657
rect 24581 15657 24593 15660
rect 24627 15657 24639 15691
rect 24581 15651 24639 15657
rect 27433 15691 27491 15697
rect 27433 15657 27445 15691
rect 27479 15688 27491 15691
rect 27798 15688 27804 15700
rect 27479 15660 27804 15688
rect 27479 15657 27491 15660
rect 27433 15651 27491 15657
rect 22830 15580 22836 15632
rect 22888 15620 22894 15632
rect 23676 15620 23704 15651
rect 27798 15648 27804 15660
rect 27856 15648 27862 15700
rect 28626 15648 28632 15700
rect 28684 15688 28690 15700
rect 28721 15691 28779 15697
rect 28721 15688 28733 15691
rect 28684 15660 28733 15688
rect 28684 15648 28690 15660
rect 28721 15657 28733 15660
rect 28767 15657 28779 15691
rect 28721 15651 28779 15657
rect 28902 15648 28908 15700
rect 28960 15688 28966 15700
rect 29089 15691 29147 15697
rect 29089 15688 29101 15691
rect 28960 15660 29101 15688
rect 28960 15648 28966 15660
rect 29089 15657 29101 15660
rect 29135 15688 29147 15691
rect 30006 15688 30012 15700
rect 29135 15660 30012 15688
rect 29135 15657 29147 15660
rect 29089 15651 29147 15657
rect 30006 15648 30012 15660
rect 30064 15648 30070 15700
rect 31297 15691 31355 15697
rect 31297 15657 31309 15691
rect 31343 15688 31355 15691
rect 32398 15688 32404 15700
rect 31343 15660 32404 15688
rect 31343 15657 31355 15660
rect 31297 15651 31355 15657
rect 32398 15648 32404 15660
rect 32456 15648 32462 15700
rect 33597 15691 33655 15697
rect 33597 15657 33609 15691
rect 33643 15688 33655 15691
rect 34238 15688 34244 15700
rect 33643 15660 34244 15688
rect 33643 15657 33655 15660
rect 33597 15651 33655 15657
rect 34238 15648 34244 15660
rect 34296 15648 34302 15700
rect 35621 15691 35679 15697
rect 35621 15657 35633 15691
rect 35667 15688 35679 15691
rect 36814 15688 36820 15700
rect 35667 15660 36820 15688
rect 35667 15657 35679 15660
rect 35621 15651 35679 15657
rect 36814 15648 36820 15660
rect 36872 15648 36878 15700
rect 43254 15648 43260 15700
rect 43312 15688 43318 15700
rect 43993 15691 44051 15697
rect 43993 15688 44005 15691
rect 43312 15660 44005 15688
rect 43312 15648 43318 15660
rect 43993 15657 44005 15660
rect 44039 15657 44051 15691
rect 43993 15651 44051 15657
rect 44177 15691 44235 15697
rect 44177 15657 44189 15691
rect 44223 15688 44235 15691
rect 44634 15688 44640 15700
rect 44223 15660 44640 15688
rect 44223 15657 44235 15660
rect 44177 15651 44235 15657
rect 44634 15648 44640 15660
rect 44692 15648 44698 15700
rect 45370 15648 45376 15700
rect 45428 15688 45434 15700
rect 45465 15691 45523 15697
rect 45465 15688 45477 15691
rect 45428 15660 45477 15688
rect 45428 15648 45434 15660
rect 45465 15657 45477 15660
rect 45511 15657 45523 15691
rect 45465 15651 45523 15657
rect 25590 15620 25596 15632
rect 22888 15592 23704 15620
rect 24596 15592 25596 15620
rect 22888 15580 22894 15592
rect 13633 15555 13691 15561
rect 13633 15521 13645 15555
rect 13679 15552 13691 15555
rect 14642 15552 14648 15564
rect 13679 15524 14648 15552
rect 13679 15521 13691 15524
rect 13633 15515 13691 15521
rect 4709 15487 4767 15493
rect 4709 15453 4721 15487
rect 4755 15484 4767 15487
rect 5994 15484 6000 15496
rect 4755 15456 6000 15484
rect 4755 15453 4767 15456
rect 4709 15447 4767 15453
rect 5994 15444 6000 15456
rect 6052 15444 6058 15496
rect 13262 15444 13268 15496
rect 13320 15484 13326 15496
rect 13541 15487 13599 15493
rect 13541 15484 13553 15487
rect 13320 15456 13553 15484
rect 13320 15444 13326 15456
rect 13541 15453 13553 15456
rect 13587 15453 13599 15487
rect 13541 15447 13599 15453
rect 13725 15487 13783 15493
rect 13725 15453 13737 15487
rect 13771 15484 13783 15487
rect 14366 15484 14372 15496
rect 13771 15456 14372 15484
rect 13771 15453 13783 15456
rect 13725 15447 13783 15453
rect 14366 15444 14372 15456
rect 14424 15444 14430 15496
rect 14568 15493 14596 15524
rect 14642 15512 14648 15524
rect 14700 15512 14706 15564
rect 15013 15555 15071 15561
rect 15013 15521 15025 15555
rect 15059 15521 15071 15555
rect 15013 15515 15071 15521
rect 15749 15555 15807 15561
rect 15749 15521 15761 15555
rect 15795 15552 15807 15555
rect 16942 15552 16948 15564
rect 15795 15524 16948 15552
rect 15795 15521 15807 15524
rect 15749 15515 15807 15521
rect 14553 15487 14611 15493
rect 14553 15453 14565 15487
rect 14599 15453 14611 15487
rect 15028 15484 15056 15515
rect 16942 15512 16948 15524
rect 17000 15512 17006 15564
rect 18325 15555 18383 15561
rect 18325 15521 18337 15555
rect 18371 15552 18383 15555
rect 19426 15552 19432 15564
rect 18371 15524 19432 15552
rect 18371 15521 18383 15524
rect 18325 15515 18383 15521
rect 19426 15512 19432 15524
rect 19484 15512 19490 15564
rect 20990 15552 20996 15564
rect 20951 15524 20996 15552
rect 20990 15512 20996 15524
rect 21048 15512 21054 15564
rect 15657 15487 15715 15493
rect 15657 15484 15669 15487
rect 15028 15456 15669 15484
rect 14553 15447 14611 15453
rect 15657 15453 15669 15456
rect 15703 15484 15715 15487
rect 15838 15484 15844 15496
rect 15703 15456 15844 15484
rect 15703 15453 15715 15456
rect 15657 15447 15715 15453
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 18046 15484 18052 15496
rect 18007 15456 18052 15484
rect 18046 15444 18052 15456
rect 18104 15444 18110 15496
rect 18230 15484 18236 15496
rect 18191 15456 18236 15484
rect 18230 15444 18236 15456
rect 18288 15444 18294 15496
rect 20438 15484 20444 15496
rect 20399 15456 20444 15484
rect 20438 15444 20444 15456
rect 20496 15444 20502 15496
rect 20806 15484 20812 15496
rect 20767 15456 20812 15484
rect 20806 15444 20812 15456
rect 20864 15444 20870 15496
rect 21450 15484 21456 15496
rect 21411 15456 21456 15484
rect 21450 15444 21456 15456
rect 21508 15444 21514 15496
rect 21637 15487 21695 15493
rect 21637 15453 21649 15487
rect 21683 15453 21695 15487
rect 21637 15447 21695 15453
rect 16022 15348 16028 15360
rect 15983 15320 16028 15348
rect 16022 15308 16028 15320
rect 16080 15308 16086 15360
rect 17862 15348 17868 15360
rect 17823 15320 17868 15348
rect 17862 15308 17868 15320
rect 17920 15308 17926 15360
rect 20254 15308 20260 15360
rect 20312 15348 20318 15360
rect 20809 15351 20867 15357
rect 20809 15348 20821 15351
rect 20312 15320 20821 15348
rect 20312 15308 20318 15320
rect 20809 15317 20821 15320
rect 20855 15348 20867 15351
rect 21652 15348 21680 15447
rect 23474 15444 23480 15496
rect 23532 15484 23538 15496
rect 24596 15493 24624 15592
rect 25590 15580 25596 15592
rect 25648 15580 25654 15632
rect 30558 15620 30564 15632
rect 29196 15592 30564 15620
rect 25498 15552 25504 15564
rect 25240 15524 25504 15552
rect 25240 15493 25268 15524
rect 25498 15512 25504 15524
rect 25556 15512 25562 15564
rect 28994 15512 29000 15564
rect 29052 15552 29058 15564
rect 29196 15561 29224 15592
rect 30558 15580 30564 15592
rect 30616 15580 30622 15632
rect 33686 15580 33692 15632
rect 33744 15620 33750 15632
rect 36170 15620 36176 15632
rect 33744 15592 36176 15620
rect 33744 15580 33750 15592
rect 29181 15555 29239 15561
rect 29181 15552 29193 15555
rect 29052 15524 29193 15552
rect 29052 15512 29058 15524
rect 29181 15521 29193 15524
rect 29227 15521 29239 15555
rect 29181 15515 29239 15521
rect 30098 15512 30104 15564
rect 30156 15552 30162 15564
rect 34057 15555 34115 15561
rect 30156 15524 30696 15552
rect 30156 15512 30162 15524
rect 23753 15487 23811 15493
rect 23753 15484 23765 15487
rect 23532 15456 23765 15484
rect 23532 15444 23538 15456
rect 23753 15453 23765 15456
rect 23799 15453 23811 15487
rect 23753 15447 23811 15453
rect 24581 15487 24639 15493
rect 24581 15453 24593 15487
rect 24627 15453 24639 15487
rect 24581 15447 24639 15453
rect 24765 15487 24823 15493
rect 24765 15453 24777 15487
rect 24811 15484 24823 15487
rect 25225 15487 25283 15493
rect 25225 15484 25237 15487
rect 24811 15456 25237 15484
rect 24811 15453 24823 15456
rect 24765 15447 24823 15453
rect 25225 15453 25237 15456
rect 25271 15453 25283 15487
rect 25225 15447 25283 15453
rect 25409 15487 25467 15493
rect 25409 15453 25421 15487
rect 25455 15484 25467 15487
rect 25590 15484 25596 15496
rect 25455 15456 25596 15484
rect 25455 15453 25467 15456
rect 25409 15447 25467 15453
rect 23768 15416 23796 15447
rect 25590 15444 25596 15456
rect 25648 15444 25654 15496
rect 26053 15487 26111 15493
rect 26053 15453 26065 15487
rect 26099 15484 26111 15487
rect 28718 15484 28724 15496
rect 26099 15456 28724 15484
rect 26099 15453 26111 15456
rect 26053 15447 26111 15453
rect 28718 15444 28724 15456
rect 28776 15444 28782 15496
rect 28905 15487 28963 15493
rect 28905 15453 28917 15487
rect 28951 15453 28963 15487
rect 28905 15447 28963 15453
rect 25317 15419 25375 15425
rect 25317 15416 25329 15419
rect 23768 15388 25329 15416
rect 25317 15385 25329 15388
rect 25363 15385 25375 15419
rect 25317 15379 25375 15385
rect 26142 15376 26148 15428
rect 26200 15416 26206 15428
rect 26298 15419 26356 15425
rect 26298 15416 26310 15419
rect 26200 15388 26310 15416
rect 26200 15376 26206 15388
rect 26298 15385 26310 15388
rect 26344 15385 26356 15419
rect 28920 15416 28948 15447
rect 30282 15444 30288 15496
rect 30340 15484 30346 15496
rect 30668 15493 30696 15524
rect 30852 15524 33824 15552
rect 30852 15496 30880 15524
rect 30377 15487 30435 15493
rect 30377 15484 30389 15487
rect 30340 15456 30389 15484
rect 30340 15444 30346 15456
rect 30377 15453 30389 15456
rect 30423 15453 30435 15487
rect 30377 15447 30435 15453
rect 30653 15487 30711 15493
rect 30653 15453 30665 15487
rect 30699 15453 30711 15487
rect 30834 15484 30840 15496
rect 30795 15456 30840 15484
rect 30653 15447 30711 15453
rect 30834 15444 30840 15456
rect 30892 15444 30898 15496
rect 31478 15484 31484 15496
rect 31439 15456 31484 15484
rect 31478 15444 31484 15456
rect 31536 15444 31542 15496
rect 31570 15444 31576 15496
rect 31628 15484 31634 15496
rect 31665 15487 31723 15493
rect 31665 15484 31677 15487
rect 31628 15456 31677 15484
rect 31628 15444 31634 15456
rect 31665 15453 31677 15456
rect 31711 15453 31723 15487
rect 31665 15447 31723 15453
rect 31754 15444 31760 15496
rect 31812 15484 31818 15496
rect 33796 15493 33824 15524
rect 34057 15521 34069 15555
rect 34103 15552 34115 15555
rect 35434 15552 35440 15564
rect 34103 15524 35440 15552
rect 34103 15521 34115 15524
rect 34057 15515 34115 15521
rect 35434 15512 35440 15524
rect 35492 15512 35498 15564
rect 32401 15487 32459 15493
rect 32401 15484 32413 15487
rect 31812 15456 31857 15484
rect 32048 15456 32413 15484
rect 31812 15444 31818 15456
rect 30193 15419 30251 15425
rect 30193 15416 30205 15419
rect 28920 15388 30205 15416
rect 26298 15379 26356 15385
rect 30193 15385 30205 15388
rect 30239 15385 30251 15419
rect 30193 15379 30251 15385
rect 30466 15376 30472 15428
rect 30524 15416 30530 15428
rect 32048 15416 32076 15456
rect 32401 15453 32413 15456
rect 32447 15453 32459 15487
rect 32401 15447 32459 15453
rect 33781 15487 33839 15493
rect 33781 15453 33793 15487
rect 33827 15453 33839 15487
rect 33781 15447 33839 15453
rect 33965 15487 34023 15493
rect 33965 15453 33977 15487
rect 34011 15453 34023 15487
rect 34146 15484 34152 15496
rect 34107 15456 34152 15484
rect 33965 15447 34023 15453
rect 30524 15388 32076 15416
rect 32217 15419 32275 15425
rect 30524 15376 30530 15388
rect 32217 15385 32229 15419
rect 32263 15416 32275 15419
rect 33042 15416 33048 15428
rect 32263 15388 33048 15416
rect 32263 15385 32275 15388
rect 32217 15379 32275 15385
rect 33042 15376 33048 15388
rect 33100 15416 33106 15428
rect 33980 15416 34008 15447
rect 34146 15444 34152 15456
rect 34204 15444 34210 15496
rect 34333 15487 34391 15493
rect 34333 15453 34345 15487
rect 34379 15453 34391 15487
rect 35452 15484 35480 15512
rect 35728 15493 35756 15592
rect 36170 15580 36176 15592
rect 36228 15580 36234 15632
rect 40313 15623 40371 15629
rect 40313 15589 40325 15623
rect 40359 15620 40371 15623
rect 40402 15620 40408 15632
rect 40359 15592 40408 15620
rect 40359 15589 40371 15592
rect 40313 15583 40371 15589
rect 40402 15580 40408 15592
rect 40460 15580 40466 15632
rect 36354 15552 36360 15564
rect 36315 15524 36360 15552
rect 36354 15512 36360 15524
rect 36412 15512 36418 15564
rect 36446 15512 36452 15564
rect 36504 15552 36510 15564
rect 36504 15524 37504 15552
rect 36504 15512 36510 15524
rect 37476 15493 37504 15524
rect 37550 15512 37556 15564
rect 37608 15552 37614 15564
rect 37829 15555 37887 15561
rect 37608 15524 37653 15552
rect 37608 15512 37614 15524
rect 37829 15521 37841 15555
rect 37875 15521 37887 15555
rect 37829 15515 37887 15521
rect 35529 15487 35587 15493
rect 35529 15484 35541 15487
rect 35452 15456 35541 15484
rect 34333 15447 34391 15453
rect 35529 15453 35541 15456
rect 35575 15453 35587 15487
rect 35529 15447 35587 15453
rect 35713 15487 35771 15493
rect 35713 15453 35725 15487
rect 35759 15453 35771 15487
rect 35713 15447 35771 15453
rect 37461 15487 37519 15493
rect 37461 15453 37473 15487
rect 37507 15453 37519 15487
rect 37844 15484 37872 15515
rect 42978 15512 42984 15564
rect 43036 15552 43042 15564
rect 43533 15555 43591 15561
rect 43533 15552 43545 15555
rect 43036 15524 43545 15552
rect 43036 15512 43042 15524
rect 43533 15521 43545 15524
rect 43579 15552 43591 15555
rect 45554 15552 45560 15564
rect 43579 15524 45560 15552
rect 43579 15521 43591 15524
rect 43533 15515 43591 15521
rect 45554 15512 45560 15524
rect 45612 15512 45618 15564
rect 38289 15487 38347 15493
rect 38289 15484 38301 15487
rect 37844 15456 38301 15484
rect 37461 15447 37519 15453
rect 38289 15453 38301 15456
rect 38335 15453 38347 15487
rect 38289 15447 38347 15453
rect 33100 15388 34008 15416
rect 34348 15416 34376 15447
rect 38470 15444 38476 15496
rect 38528 15484 38534 15496
rect 39850 15484 39856 15496
rect 38528 15456 39856 15484
rect 38528 15444 38534 15456
rect 39850 15444 39856 15456
rect 39908 15444 39914 15496
rect 40034 15484 40040 15496
rect 39995 15456 40040 15484
rect 40034 15444 40040 15456
rect 40092 15444 40098 15496
rect 40126 15444 40132 15496
rect 40184 15484 40190 15496
rect 40313 15487 40371 15493
rect 40313 15484 40325 15487
rect 40184 15456 40325 15484
rect 40184 15444 40190 15456
rect 40313 15453 40325 15456
rect 40359 15453 40371 15487
rect 40313 15447 40371 15453
rect 42242 15444 42248 15496
rect 42300 15484 42306 15496
rect 42521 15487 42579 15493
rect 42521 15484 42533 15487
rect 42300 15456 42533 15484
rect 42300 15444 42306 15456
rect 42521 15453 42533 15456
rect 42567 15453 42579 15487
rect 42521 15447 42579 15453
rect 42705 15487 42763 15493
rect 42705 15453 42717 15487
rect 42751 15484 42763 15487
rect 43254 15484 43260 15496
rect 42751 15456 43260 15484
rect 42751 15453 42763 15456
rect 42705 15447 42763 15453
rect 43254 15444 43260 15456
rect 43312 15444 43318 15496
rect 43346 15444 43352 15496
rect 43404 15484 43410 15496
rect 43404 15456 44404 15484
rect 43404 15444 43410 15456
rect 38381 15419 38439 15425
rect 38381 15416 38393 15419
rect 34348 15388 38393 15416
rect 33100 15376 33106 15388
rect 38381 15385 38393 15388
rect 38427 15385 38439 15419
rect 42334 15416 42340 15428
rect 42295 15388 42340 15416
rect 38381 15379 38439 15385
rect 42334 15376 42340 15388
rect 42392 15376 42398 15428
rect 44174 15425 44180 15428
rect 44161 15419 44180 15425
rect 44161 15385 44173 15419
rect 44161 15379 44180 15385
rect 44174 15376 44180 15379
rect 44232 15376 44238 15428
rect 44376 15425 44404 15456
rect 44450 15444 44456 15496
rect 44508 15484 44514 15496
rect 45189 15487 45247 15493
rect 45189 15484 45201 15487
rect 44508 15456 45201 15484
rect 44508 15444 44514 15456
rect 45189 15453 45201 15456
rect 45235 15453 45247 15487
rect 45189 15447 45247 15453
rect 45278 15444 45284 15496
rect 45336 15484 45342 15496
rect 47673 15487 47731 15493
rect 45336 15456 45381 15484
rect 45336 15444 45342 15456
rect 47673 15453 47685 15487
rect 47719 15484 47731 15487
rect 48314 15484 48320 15496
rect 47719 15456 48320 15484
rect 47719 15453 47731 15456
rect 47673 15447 47731 15453
rect 48314 15444 48320 15456
rect 48372 15444 48378 15496
rect 44361 15419 44419 15425
rect 44361 15385 44373 15419
rect 44407 15416 44419 15419
rect 45002 15416 45008 15428
rect 44407 15388 45008 15416
rect 44407 15385 44419 15388
rect 44361 15379 44419 15385
rect 45002 15376 45008 15388
rect 45060 15376 45066 15428
rect 45462 15416 45468 15428
rect 45423 15388 45468 15416
rect 45462 15376 45468 15388
rect 45520 15376 45526 15428
rect 20855 15320 21680 15348
rect 32585 15351 32643 15357
rect 20855 15317 20867 15320
rect 20809 15311 20867 15317
rect 32585 15317 32597 15351
rect 32631 15348 32643 15351
rect 33318 15348 33324 15360
rect 32631 15320 33324 15348
rect 32631 15317 32643 15320
rect 32585 15311 32643 15317
rect 33318 15308 33324 15320
rect 33376 15308 33382 15360
rect 36170 15348 36176 15360
rect 36131 15320 36176 15348
rect 36170 15308 36176 15320
rect 36228 15308 36234 15360
rect 36814 15348 36820 15360
rect 36775 15320 36820 15348
rect 36814 15308 36820 15320
rect 36872 15308 36878 15360
rect 40129 15351 40187 15357
rect 40129 15317 40141 15351
rect 40175 15348 40187 15351
rect 40310 15348 40316 15360
rect 40175 15320 40316 15348
rect 40175 15317 40187 15320
rect 40129 15311 40187 15317
rect 40310 15308 40316 15320
rect 40368 15308 40374 15360
rect 43530 15348 43536 15360
rect 43491 15320 43536 15348
rect 43530 15308 43536 15320
rect 43588 15308 43594 15360
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 14274 15144 14280 15156
rect 14235 15116 14280 15144
rect 14274 15104 14280 15116
rect 14332 15104 14338 15156
rect 19981 15147 20039 15153
rect 19981 15113 19993 15147
rect 20027 15144 20039 15147
rect 20438 15144 20444 15156
rect 20027 15116 20444 15144
rect 20027 15113 20039 15116
rect 19981 15107 20039 15113
rect 20438 15104 20444 15116
rect 20496 15144 20502 15156
rect 20733 15147 20791 15153
rect 20733 15144 20745 15147
rect 20496 15116 20745 15144
rect 20496 15104 20502 15116
rect 20733 15113 20745 15116
rect 20779 15113 20791 15147
rect 20733 15107 20791 15113
rect 20901 15147 20959 15153
rect 20901 15113 20913 15147
rect 20947 15144 20959 15147
rect 21450 15144 21456 15156
rect 20947 15116 21456 15144
rect 20947 15113 20959 15116
rect 20901 15107 20959 15113
rect 21450 15104 21456 15116
rect 21508 15104 21514 15156
rect 30101 15147 30159 15153
rect 30101 15113 30113 15147
rect 30147 15144 30159 15147
rect 30466 15144 30472 15156
rect 30147 15116 30472 15144
rect 30147 15113 30159 15116
rect 30101 15107 30159 15113
rect 30466 15104 30472 15116
rect 30524 15104 30530 15156
rect 31205 15147 31263 15153
rect 31205 15113 31217 15147
rect 31251 15144 31263 15147
rect 31478 15144 31484 15156
rect 31251 15116 31484 15144
rect 31251 15113 31263 15116
rect 31205 15107 31263 15113
rect 31478 15104 31484 15116
rect 31536 15104 31542 15156
rect 37734 15104 37740 15156
rect 37792 15144 37798 15156
rect 37829 15147 37887 15153
rect 37829 15144 37841 15147
rect 37792 15116 37841 15144
rect 37792 15104 37798 15116
rect 37829 15113 37841 15116
rect 37875 15113 37887 15147
rect 37829 15107 37887 15113
rect 3418 15036 3424 15088
rect 3476 15076 3482 15088
rect 4157 15079 4215 15085
rect 4157 15076 4169 15079
rect 3476 15048 4169 15076
rect 3476 15036 3482 15048
rect 4157 15045 4169 15048
rect 4203 15045 4215 15079
rect 4157 15039 4215 15045
rect 17764 15079 17822 15085
rect 17764 15045 17776 15079
rect 17810 15076 17822 15079
rect 17862 15076 17868 15088
rect 17810 15048 17868 15076
rect 17810 15045 17822 15048
rect 17764 15039 17822 15045
rect 17862 15036 17868 15048
rect 17920 15036 17926 15088
rect 20533 15079 20591 15085
rect 20533 15045 20545 15079
rect 20579 15076 20591 15079
rect 24296 15079 24354 15085
rect 20579 15048 20852 15076
rect 20579 15045 20591 15048
rect 20533 15039 20591 15045
rect 20824 15020 20852 15048
rect 24296 15045 24308 15079
rect 24342 15076 24354 15079
rect 25406 15076 25412 15088
rect 24342 15048 25412 15076
rect 24342 15045 24354 15048
rect 24296 15039 24354 15045
rect 25406 15036 25412 15048
rect 25464 15036 25470 15088
rect 30650 15036 30656 15088
rect 30708 15076 30714 15088
rect 30708 15048 30788 15076
rect 30708 15036 30714 15048
rect 5994 14968 6000 15020
rect 6052 15008 6058 15020
rect 6052 14980 6097 15008
rect 6052 14968 6058 14980
rect 13262 14968 13268 15020
rect 13320 15008 13326 15020
rect 14185 15011 14243 15017
rect 14185 15008 14197 15011
rect 13320 14980 14197 15008
rect 13320 14968 13326 14980
rect 14185 14977 14197 14980
rect 14231 14977 14243 15011
rect 14366 15008 14372 15020
rect 14327 14980 14372 15008
rect 14185 14971 14243 14977
rect 14366 14968 14372 14980
rect 14424 14968 14430 15020
rect 17494 15008 17500 15020
rect 17455 14980 17500 15008
rect 17494 14968 17500 14980
rect 17552 14968 17558 15020
rect 19426 14968 19432 15020
rect 19484 15008 19490 15020
rect 19889 15011 19947 15017
rect 19889 15008 19901 15011
rect 19484 14980 19901 15008
rect 19484 14968 19490 14980
rect 19889 14977 19901 14980
rect 19935 14977 19947 15011
rect 19889 14971 19947 14977
rect 20073 15011 20131 15017
rect 20073 14977 20085 15011
rect 20119 15008 20131 15011
rect 20162 15008 20168 15020
rect 20119 14980 20168 15008
rect 20119 14977 20131 14980
rect 20073 14971 20131 14977
rect 20162 14968 20168 14980
rect 20220 14968 20226 15020
rect 20806 14968 20812 15020
rect 20864 14968 20870 15020
rect 25774 14968 25780 15020
rect 25832 15008 25838 15020
rect 26145 15011 26203 15017
rect 26145 15008 26157 15011
rect 25832 14980 26157 15008
rect 25832 14968 25838 14980
rect 26145 14977 26157 14980
rect 26191 14977 26203 15011
rect 26145 14971 26203 14977
rect 26329 15011 26387 15017
rect 26329 14977 26341 15011
rect 26375 15008 26387 15011
rect 26510 15008 26516 15020
rect 26375 14980 26516 15008
rect 26375 14977 26387 14980
rect 26329 14971 26387 14977
rect 26510 14968 26516 14980
rect 26568 15008 26574 15020
rect 27430 15008 27436 15020
rect 26568 14980 27436 15008
rect 26568 14968 26574 14980
rect 27430 14968 27436 14980
rect 27488 14968 27494 15020
rect 28718 15008 28724 15020
rect 28679 14980 28724 15008
rect 28718 14968 28724 14980
rect 28776 14968 28782 15020
rect 28988 15011 29046 15017
rect 28988 14977 29000 15011
rect 29034 15008 29046 15011
rect 30466 15008 30472 15020
rect 29034 14980 30472 15008
rect 29034 14977 29046 14980
rect 28988 14971 29046 14977
rect 30466 14968 30472 14980
rect 30524 14968 30530 15020
rect 30558 14968 30564 15020
rect 30616 15008 30622 15020
rect 30760 15017 30788 15048
rect 43254 15036 43260 15088
rect 43312 15076 43318 15088
rect 43312 15048 44864 15076
rect 43312 15036 43318 15048
rect 30745 15011 30803 15017
rect 30616 14980 30661 15008
rect 30616 14968 30622 14980
rect 30745 14977 30757 15011
rect 30791 14977 30803 15011
rect 30745 14971 30803 14977
rect 30834 14968 30840 15020
rect 30892 15008 30898 15020
rect 31021 15011 31079 15017
rect 31021 15008 31033 15011
rect 30892 14980 31033 15008
rect 30892 14968 30898 14980
rect 31021 14977 31033 14980
rect 31067 14977 31079 15011
rect 32306 15008 32312 15020
rect 32267 14980 32312 15008
rect 31021 14971 31079 14977
rect 32306 14968 32312 14980
rect 32364 14968 32370 15020
rect 32582 15017 32588 15020
rect 32576 14971 32588 15017
rect 32640 15008 32646 15020
rect 35437 15011 35495 15017
rect 32640 14980 32676 15008
rect 32582 14968 32588 14971
rect 32640 14968 32646 14980
rect 35437 14977 35449 15011
rect 35483 15008 35495 15011
rect 36170 15008 36176 15020
rect 35483 14980 36176 15008
rect 35483 14977 35495 14980
rect 35437 14971 35495 14977
rect 36170 14968 36176 14980
rect 36228 14968 36234 15020
rect 36354 14968 36360 15020
rect 36412 15008 36418 15020
rect 36633 15011 36691 15017
rect 36633 15008 36645 15011
rect 36412 14980 36645 15008
rect 36412 14968 36418 14980
rect 36633 14977 36645 14980
rect 36679 14977 36691 15011
rect 36814 15008 36820 15020
rect 36775 14980 36820 15008
rect 36633 14971 36691 14977
rect 36814 14968 36820 14980
rect 36872 14968 36878 15020
rect 36906 14968 36912 15020
rect 36964 15008 36970 15020
rect 37461 15011 37519 15017
rect 37461 15008 37473 15011
rect 36964 14980 37473 15008
rect 36964 14968 36970 14980
rect 37461 14977 37473 14980
rect 37507 14977 37519 15011
rect 37461 14971 37519 14977
rect 40313 15011 40371 15017
rect 40313 14977 40325 15011
rect 40359 15008 40371 15011
rect 41509 15011 41567 15017
rect 40359 14980 40816 15008
rect 40359 14977 40371 14980
rect 40313 14971 40371 14977
rect 5074 14900 5080 14952
rect 5132 14940 5138 14952
rect 5813 14943 5871 14949
rect 5813 14940 5825 14943
rect 5132 14912 5825 14940
rect 5132 14900 5138 14912
rect 5813 14909 5825 14912
rect 5859 14909 5871 14943
rect 5813 14903 5871 14909
rect 22646 14900 22652 14952
rect 22704 14940 22710 14952
rect 24029 14943 24087 14949
rect 24029 14940 24041 14943
rect 22704 14912 24041 14940
rect 22704 14900 22710 14912
rect 24029 14909 24041 14912
rect 24075 14909 24087 14943
rect 24029 14903 24087 14909
rect 26421 14943 26479 14949
rect 26421 14909 26433 14943
rect 26467 14940 26479 14943
rect 26602 14940 26608 14952
rect 26467 14912 26608 14940
rect 26467 14909 26479 14912
rect 26421 14903 26479 14909
rect 26602 14900 26608 14912
rect 26660 14900 26666 14952
rect 35529 14943 35587 14949
rect 35529 14909 35541 14943
rect 35575 14909 35587 14943
rect 35529 14903 35587 14909
rect 36725 14943 36783 14949
rect 36725 14909 36737 14943
rect 36771 14940 36783 14943
rect 37550 14940 37556 14952
rect 36771 14912 37556 14940
rect 36771 14909 36783 14912
rect 36725 14903 36783 14909
rect 25409 14875 25467 14881
rect 25409 14841 25421 14875
rect 25455 14872 25467 14875
rect 25590 14872 25596 14884
rect 25455 14844 25596 14872
rect 25455 14841 25467 14844
rect 25409 14835 25467 14841
rect 25590 14832 25596 14844
rect 25648 14832 25654 14884
rect 33689 14875 33747 14881
rect 33689 14841 33701 14875
rect 33735 14872 33747 14875
rect 33962 14872 33968 14884
rect 33735 14844 33968 14872
rect 33735 14841 33747 14844
rect 33689 14835 33747 14841
rect 33962 14832 33968 14844
rect 34020 14832 34026 14884
rect 35434 14832 35440 14884
rect 35492 14872 35498 14884
rect 35544 14872 35572 14903
rect 37550 14900 37556 14912
rect 37608 14900 37614 14952
rect 40402 14940 40408 14952
rect 40363 14912 40408 14940
rect 40402 14900 40408 14912
rect 40460 14900 40466 14952
rect 40788 14872 40816 14980
rect 41509 14977 41521 15011
rect 41555 15008 41567 15011
rect 42886 15008 42892 15020
rect 41555 14980 42892 15008
rect 41555 14977 41567 14980
rect 41509 14971 41567 14977
rect 42886 14968 42892 14980
rect 42944 14968 42950 15020
rect 43530 14968 43536 15020
rect 43588 15008 43594 15020
rect 44836 15017 44864 15048
rect 43993 15011 44051 15017
rect 43993 15008 44005 15011
rect 43588 14980 44005 15008
rect 43588 14968 43594 14980
rect 43993 14977 44005 14980
rect 44039 14977 44051 15011
rect 43993 14971 44051 14977
rect 44821 15011 44879 15017
rect 44821 14977 44833 15011
rect 44867 14977 44879 15011
rect 45002 15008 45008 15020
rect 44963 14980 45008 15008
rect 44821 14971 44879 14977
rect 45002 14968 45008 14980
rect 45060 14968 45066 15020
rect 47486 14968 47492 15020
rect 47544 15008 47550 15020
rect 47765 15011 47823 15017
rect 47765 15008 47777 15011
rect 47544 14980 47777 15008
rect 47544 14968 47550 14980
rect 47765 14977 47777 14980
rect 47811 14977 47823 15011
rect 47765 14971 47823 14977
rect 40954 14900 40960 14952
rect 41012 14940 41018 14952
rect 41417 14943 41475 14949
rect 41417 14940 41429 14943
rect 41012 14912 41429 14940
rect 41012 14900 41018 14912
rect 41417 14909 41429 14912
rect 41463 14909 41475 14943
rect 41417 14903 41475 14909
rect 42981 14943 43039 14949
rect 42981 14909 42993 14943
rect 43027 14909 43039 14943
rect 42981 14903 43039 14909
rect 43257 14943 43315 14949
rect 43257 14909 43269 14943
rect 43303 14940 43315 14943
rect 43346 14940 43352 14952
rect 43303 14912 43352 14940
rect 43303 14909 43315 14912
rect 43257 14903 43315 14909
rect 41138 14872 41144 14884
rect 35492 14844 37504 14872
rect 40788 14844 41144 14872
rect 35492 14832 35498 14844
rect 2317 14807 2375 14813
rect 2317 14773 2329 14807
rect 2363 14804 2375 14807
rect 3418 14804 3424 14816
rect 2363 14776 3424 14804
rect 2363 14773 2375 14776
rect 2317 14767 2375 14773
rect 3418 14764 3424 14776
rect 3476 14764 3482 14816
rect 18782 14764 18788 14816
rect 18840 14804 18846 14816
rect 18877 14807 18935 14813
rect 18877 14804 18889 14807
rect 18840 14776 18889 14804
rect 18840 14764 18846 14776
rect 18877 14773 18889 14776
rect 18923 14773 18935 14807
rect 18877 14767 18935 14773
rect 20717 14807 20775 14813
rect 20717 14773 20729 14807
rect 20763 14804 20775 14807
rect 20990 14804 20996 14816
rect 20763 14776 20996 14804
rect 20763 14773 20775 14776
rect 20717 14767 20775 14773
rect 20990 14764 20996 14776
rect 21048 14764 21054 14816
rect 25961 14807 26019 14813
rect 25961 14773 25973 14807
rect 26007 14804 26019 14807
rect 26234 14804 26240 14816
rect 26007 14776 26240 14804
rect 26007 14773 26019 14776
rect 25961 14767 26019 14773
rect 26234 14764 26240 14776
rect 26292 14764 26298 14816
rect 33870 14764 33876 14816
rect 33928 14804 33934 14816
rect 37476 14813 37504 14844
rect 41138 14832 41144 14844
rect 41196 14832 41202 14884
rect 42996 14872 43024 14903
rect 43346 14900 43352 14912
rect 43404 14900 43410 14952
rect 43901 14943 43959 14949
rect 43901 14909 43913 14943
rect 43947 14909 43959 14943
rect 44266 14940 44272 14952
rect 44227 14912 44272 14940
rect 43901 14903 43959 14909
rect 43916 14872 43944 14903
rect 44266 14900 44272 14912
rect 44324 14900 44330 14952
rect 44358 14900 44364 14952
rect 44416 14940 44422 14952
rect 44416 14912 44461 14940
rect 44416 14900 44422 14912
rect 45189 14875 45247 14881
rect 45189 14872 45201 14875
rect 42996 14844 43852 14872
rect 43916 14844 45201 14872
rect 35161 14807 35219 14813
rect 35161 14804 35173 14807
rect 33928 14776 35173 14804
rect 33928 14764 33934 14776
rect 35161 14773 35173 14776
rect 35207 14773 35219 14807
rect 35161 14767 35219 14773
rect 37461 14807 37519 14813
rect 37461 14773 37473 14807
rect 37507 14773 37519 14807
rect 37461 14767 37519 14773
rect 40589 14807 40647 14813
rect 40589 14773 40601 14807
rect 40635 14804 40647 14807
rect 40862 14804 40868 14816
rect 40635 14776 40868 14804
rect 40635 14773 40647 14776
rect 40589 14767 40647 14773
rect 40862 14764 40868 14776
rect 40920 14764 40926 14816
rect 43714 14804 43720 14816
rect 43675 14776 43720 14804
rect 43714 14764 43720 14776
rect 43772 14764 43778 14816
rect 43824 14804 43852 14844
rect 45189 14841 45201 14844
rect 45235 14872 45247 14875
rect 45462 14872 45468 14884
rect 45235 14844 45468 14872
rect 45235 14841 45247 14844
rect 45189 14835 45247 14841
rect 45462 14832 45468 14844
rect 45520 14832 45526 14884
rect 44358 14804 44364 14816
rect 43824 14776 44364 14804
rect 44358 14764 44364 14776
rect 44416 14764 44422 14816
rect 47857 14807 47915 14813
rect 47857 14773 47869 14807
rect 47903 14804 47915 14807
rect 48130 14804 48136 14816
rect 47903 14776 48136 14804
rect 47903 14773 47915 14776
rect 47857 14767 47915 14773
rect 48130 14764 48136 14776
rect 48188 14764 48194 14816
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 5074 14600 5080 14612
rect 5035 14572 5080 14600
rect 5074 14560 5080 14572
rect 5132 14560 5138 14612
rect 18046 14560 18052 14612
rect 18104 14600 18110 14612
rect 18141 14603 18199 14609
rect 18141 14600 18153 14603
rect 18104 14572 18153 14600
rect 18104 14560 18110 14572
rect 18141 14569 18153 14572
rect 18187 14569 18199 14603
rect 20162 14600 20168 14612
rect 20123 14572 20168 14600
rect 18141 14563 18199 14569
rect 20162 14560 20168 14572
rect 20220 14560 20226 14612
rect 21082 14560 21088 14612
rect 21140 14600 21146 14612
rect 21269 14603 21327 14609
rect 21269 14600 21281 14603
rect 21140 14572 21281 14600
rect 21140 14560 21146 14572
rect 21269 14569 21281 14572
rect 21315 14569 21327 14603
rect 21269 14563 21327 14569
rect 30466 14560 30472 14612
rect 30524 14600 30530 14612
rect 31297 14603 31355 14609
rect 31297 14600 31309 14603
rect 30524 14572 31309 14600
rect 30524 14560 30530 14572
rect 31297 14569 31309 14572
rect 31343 14569 31355 14603
rect 32582 14600 32588 14612
rect 32543 14572 32588 14600
rect 31297 14563 31355 14569
rect 32582 14560 32588 14572
rect 32640 14560 32646 14612
rect 33594 14600 33600 14612
rect 32876 14572 33600 14600
rect 20438 14532 20444 14544
rect 16776 14504 20444 14532
rect 3418 14464 3424 14476
rect 3379 14436 3424 14464
rect 3418 14424 3424 14436
rect 3476 14424 3482 14476
rect 14366 14424 14372 14476
rect 14424 14464 14430 14476
rect 14829 14467 14887 14473
rect 14829 14464 14841 14467
rect 14424 14436 14841 14464
rect 14424 14424 14430 14436
rect 14829 14433 14841 14436
rect 14875 14433 14887 14467
rect 14829 14427 14887 14433
rect 14918 14424 14924 14476
rect 14976 14464 14982 14476
rect 15013 14467 15071 14473
rect 15013 14464 15025 14467
rect 14976 14436 15025 14464
rect 14976 14424 14982 14436
rect 15013 14433 15025 14436
rect 15059 14433 15071 14467
rect 15013 14427 15071 14433
rect 1578 14396 1584 14408
rect 1539 14368 1584 14396
rect 1578 14356 1584 14368
rect 1636 14356 1642 14408
rect 5169 14399 5227 14405
rect 5169 14365 5181 14399
rect 5215 14396 5227 14399
rect 5810 14396 5816 14408
rect 5215 14368 5816 14396
rect 5215 14365 5227 14368
rect 5169 14359 5227 14365
rect 5810 14356 5816 14368
rect 5868 14356 5874 14408
rect 13725 14399 13783 14405
rect 13725 14365 13737 14399
rect 13771 14396 13783 14399
rect 15028 14396 15056 14427
rect 16022 14424 16028 14476
rect 16080 14464 16086 14476
rect 16776 14473 16804 14504
rect 20438 14492 20444 14504
rect 20496 14492 20502 14544
rect 30006 14492 30012 14544
rect 30064 14532 30070 14544
rect 30929 14535 30987 14541
rect 30929 14532 30941 14535
rect 30064 14504 30941 14532
rect 30064 14492 30070 14504
rect 30929 14501 30941 14504
rect 30975 14501 30987 14535
rect 30929 14495 30987 14501
rect 16577 14467 16635 14473
rect 16577 14464 16589 14467
rect 16080 14436 16589 14464
rect 16080 14424 16086 14436
rect 16577 14433 16589 14436
rect 16623 14433 16635 14467
rect 16577 14427 16635 14433
rect 16761 14467 16819 14473
rect 16761 14433 16773 14467
rect 16807 14433 16819 14467
rect 25682 14464 25688 14476
rect 16761 14427 16819 14433
rect 18340 14436 25688 14464
rect 18340 14408 18368 14436
rect 25682 14424 25688 14436
rect 25740 14424 25746 14476
rect 30377 14467 30435 14473
rect 30377 14433 30389 14467
rect 30423 14464 30435 14467
rect 30423 14436 31156 14464
rect 30423 14433 30435 14436
rect 30377 14427 30435 14433
rect 17494 14396 17500 14408
rect 13771 14368 14412 14396
rect 15028 14368 17500 14396
rect 13771 14365 13783 14368
rect 13725 14359 13783 14365
rect 2406 14288 2412 14340
rect 2464 14328 2470 14340
rect 3237 14331 3295 14337
rect 3237 14328 3249 14331
rect 2464 14300 3249 14328
rect 2464 14288 2470 14300
rect 3237 14297 3249 14300
rect 3283 14297 3295 14331
rect 3237 14291 3295 14297
rect 13446 14220 13452 14272
rect 13504 14260 13510 14272
rect 14384 14269 14412 14368
rect 17494 14356 17500 14368
rect 17552 14356 17558 14408
rect 18322 14396 18328 14408
rect 18235 14368 18328 14396
rect 18322 14356 18328 14368
rect 18380 14356 18386 14408
rect 18506 14356 18512 14408
rect 18564 14396 18570 14408
rect 18601 14399 18659 14405
rect 18601 14396 18613 14399
rect 18564 14368 18613 14396
rect 18564 14356 18570 14368
rect 18601 14365 18613 14368
rect 18647 14365 18659 14399
rect 18782 14396 18788 14408
rect 18743 14368 18788 14396
rect 18601 14359 18659 14365
rect 18782 14356 18788 14368
rect 18840 14396 18846 14408
rect 19978 14396 19984 14408
rect 18840 14368 19984 14396
rect 18840 14356 18846 14368
rect 19978 14356 19984 14368
rect 20036 14356 20042 14408
rect 21082 14396 21088 14408
rect 21043 14368 21088 14396
rect 21082 14356 21088 14368
rect 21140 14356 21146 14408
rect 21358 14396 21364 14408
rect 21319 14368 21364 14396
rect 21358 14356 21364 14368
rect 21416 14356 21422 14408
rect 26234 14356 26240 14408
rect 26292 14396 26298 14408
rect 26614 14399 26672 14405
rect 26614 14396 26626 14399
rect 26292 14368 26626 14396
rect 26292 14356 26298 14368
rect 26614 14365 26626 14368
rect 26660 14365 26672 14399
rect 26614 14359 26672 14365
rect 26881 14399 26939 14405
rect 26881 14365 26893 14399
rect 26927 14396 26939 14399
rect 28718 14396 28724 14408
rect 26927 14368 28724 14396
rect 26927 14365 26939 14368
rect 26881 14359 26939 14365
rect 28718 14356 28724 14368
rect 28776 14356 28782 14408
rect 29733 14399 29791 14405
rect 29733 14365 29745 14399
rect 29779 14365 29791 14399
rect 29733 14359 29791 14365
rect 29917 14399 29975 14405
rect 29917 14365 29929 14399
rect 29963 14396 29975 14399
rect 30098 14396 30104 14408
rect 29963 14368 30104 14396
rect 29963 14365 29975 14368
rect 29917 14359 29975 14365
rect 14737 14331 14795 14337
rect 14737 14297 14749 14331
rect 14783 14328 14795 14331
rect 19797 14331 19855 14337
rect 14783 14300 16160 14328
rect 14783 14297 14795 14300
rect 14737 14291 14795 14297
rect 16132 14269 16160 14300
rect 19797 14297 19809 14331
rect 19843 14328 19855 14331
rect 20070 14328 20076 14340
rect 19843 14300 20076 14328
rect 19843 14297 19855 14300
rect 19797 14291 19855 14297
rect 20070 14288 20076 14300
rect 20128 14288 20134 14340
rect 21376 14328 21404 14356
rect 29748 14328 29776 14359
rect 30098 14356 30104 14368
rect 30156 14356 30162 14408
rect 30193 14399 30251 14405
rect 30193 14365 30205 14399
rect 30239 14396 30251 14399
rect 30282 14396 30288 14408
rect 30239 14368 30288 14396
rect 30239 14365 30251 14368
rect 30193 14359 30251 14365
rect 30282 14356 30288 14368
rect 30340 14356 30346 14408
rect 31128 14405 31156 14436
rect 30837 14399 30895 14405
rect 30837 14365 30849 14399
rect 30883 14365 30895 14399
rect 30837 14359 30895 14365
rect 31113 14399 31171 14405
rect 31113 14365 31125 14399
rect 31159 14365 31171 14399
rect 31113 14359 31171 14365
rect 32769 14399 32827 14405
rect 32769 14365 32781 14399
rect 32815 14365 32827 14399
rect 32876 14396 32904 14572
rect 33594 14560 33600 14572
rect 33652 14560 33658 14612
rect 33965 14603 34023 14609
rect 33965 14569 33977 14603
rect 34011 14600 34023 14603
rect 35069 14603 35127 14609
rect 35069 14600 35081 14603
rect 34011 14572 35081 14600
rect 34011 14569 34023 14572
rect 33965 14563 34023 14569
rect 35069 14569 35081 14572
rect 35115 14569 35127 14603
rect 35434 14600 35440 14612
rect 35395 14572 35440 14600
rect 35069 14563 35127 14569
rect 34146 14532 34152 14544
rect 32968 14504 34152 14532
rect 32968 14473 32996 14504
rect 34146 14492 34152 14504
rect 34204 14492 34210 14544
rect 32953 14467 33011 14473
rect 32953 14433 32965 14467
rect 32999 14433 33011 14467
rect 33870 14464 33876 14476
rect 32953 14427 33011 14433
rect 33152 14436 33876 14464
rect 33152 14405 33180 14436
rect 33870 14424 33876 14436
rect 33928 14424 33934 14476
rect 33045 14399 33103 14405
rect 33045 14396 33057 14399
rect 32876 14368 33057 14396
rect 32769 14359 32827 14365
rect 33045 14365 33057 14368
rect 33091 14365 33103 14399
rect 33045 14359 33103 14365
rect 33137 14399 33195 14405
rect 33137 14365 33149 14399
rect 33183 14365 33195 14399
rect 33318 14396 33324 14408
rect 33279 14368 33324 14396
rect 33137 14359 33195 14365
rect 30374 14328 30380 14340
rect 21376 14300 29684 14328
rect 29748 14300 30380 14328
rect 13541 14263 13599 14269
rect 13541 14260 13553 14263
rect 13504 14232 13553 14260
rect 13504 14220 13510 14232
rect 13541 14229 13553 14232
rect 13587 14229 13599 14263
rect 13541 14223 13599 14229
rect 14369 14263 14427 14269
rect 14369 14229 14381 14263
rect 14415 14229 14427 14263
rect 14369 14223 14427 14229
rect 16117 14263 16175 14269
rect 16117 14229 16129 14263
rect 16163 14229 16175 14263
rect 16117 14223 16175 14229
rect 16485 14263 16543 14269
rect 16485 14229 16497 14263
rect 16531 14260 16543 14263
rect 20346 14260 20352 14272
rect 16531 14232 20352 14260
rect 16531 14229 16543 14232
rect 16485 14223 16543 14229
rect 20346 14220 20352 14232
rect 20404 14220 20410 14272
rect 20898 14260 20904 14272
rect 20859 14232 20904 14260
rect 20898 14220 20904 14232
rect 20956 14220 20962 14272
rect 25498 14260 25504 14272
rect 25459 14232 25504 14260
rect 25498 14220 25504 14232
rect 25556 14220 25562 14272
rect 29656 14260 29684 14300
rect 30374 14288 30380 14300
rect 30432 14288 30438 14340
rect 29914 14260 29920 14272
rect 29656 14232 29920 14260
rect 29914 14220 29920 14232
rect 29972 14260 29978 14272
rect 30852 14260 30880 14359
rect 32784 14328 32812 14359
rect 33318 14356 33324 14368
rect 33376 14356 33382 14408
rect 33410 14356 33416 14408
rect 33468 14396 33474 14408
rect 33781 14399 33839 14405
rect 33781 14396 33793 14399
rect 33468 14368 33793 14396
rect 33468 14356 33474 14368
rect 33781 14365 33793 14368
rect 33827 14365 33839 14399
rect 33962 14396 33968 14408
rect 33923 14368 33968 14396
rect 33781 14359 33839 14365
rect 33962 14356 33968 14368
rect 34020 14356 34026 14408
rect 34974 14396 34980 14408
rect 34935 14368 34980 14396
rect 34974 14356 34980 14368
rect 35032 14356 35038 14408
rect 35084 14396 35112 14563
rect 35434 14560 35440 14572
rect 35492 14560 35498 14612
rect 40954 14560 40960 14612
rect 41012 14600 41018 14612
rect 41601 14603 41659 14609
rect 41601 14600 41613 14603
rect 41012 14572 41613 14600
rect 41012 14560 41018 14572
rect 41601 14569 41613 14572
rect 41647 14569 41659 14603
rect 41601 14563 41659 14569
rect 44358 14560 44364 14612
rect 44416 14600 44422 14612
rect 44637 14603 44695 14609
rect 44637 14600 44649 14603
rect 44416 14572 44649 14600
rect 44416 14560 44422 14572
rect 44637 14569 44649 14572
rect 44683 14569 44695 14603
rect 44637 14563 44695 14569
rect 36354 14492 36360 14544
rect 36412 14532 36418 14544
rect 36449 14535 36507 14541
rect 36449 14532 36461 14535
rect 36412 14504 36461 14532
rect 36412 14492 36418 14504
rect 36449 14501 36461 14504
rect 36495 14501 36507 14535
rect 36449 14495 36507 14501
rect 36630 14464 36636 14476
rect 36591 14436 36636 14464
rect 36630 14424 36636 14436
rect 36688 14424 36694 14476
rect 46842 14464 46848 14476
rect 46803 14436 46848 14464
rect 46842 14424 46848 14436
rect 46900 14424 46906 14476
rect 48130 14464 48136 14476
rect 48091 14436 48136 14464
rect 48130 14424 48136 14436
rect 48188 14424 48194 14476
rect 48314 14464 48320 14476
rect 48275 14436 48320 14464
rect 48314 14424 48320 14436
rect 48372 14424 48378 14476
rect 36357 14399 36415 14405
rect 36357 14396 36369 14399
rect 35084 14368 36369 14396
rect 36357 14365 36369 14368
rect 36403 14396 36415 14399
rect 36446 14396 36452 14408
rect 36403 14368 36452 14396
rect 36403 14365 36415 14368
rect 36357 14359 36415 14365
rect 36446 14356 36452 14368
rect 36504 14356 36510 14408
rect 40218 14396 40224 14408
rect 40131 14368 40224 14396
rect 40218 14356 40224 14368
rect 40276 14396 40282 14408
rect 43257 14399 43315 14405
rect 43257 14396 43269 14399
rect 40276 14368 43269 14396
rect 40276 14356 40282 14368
rect 43257 14365 43269 14368
rect 43303 14396 43315 14399
rect 46106 14396 46112 14408
rect 43303 14368 46112 14396
rect 43303 14365 43315 14368
rect 43257 14359 43315 14365
rect 46106 14356 46112 14368
rect 46164 14356 46170 14408
rect 33980 14328 34008 14356
rect 40494 14337 40500 14340
rect 32784 14300 34008 14328
rect 33060 14272 33088 14300
rect 40488 14291 40500 14337
rect 40552 14328 40558 14340
rect 43524 14331 43582 14337
rect 40552 14300 40588 14328
rect 40494 14288 40500 14291
rect 40552 14288 40558 14300
rect 43524 14297 43536 14331
rect 43570 14328 43582 14331
rect 43714 14328 43720 14340
rect 43570 14300 43720 14328
rect 43570 14297 43582 14300
rect 43524 14291 43582 14297
rect 43714 14288 43720 14300
rect 43772 14288 43778 14340
rect 29972 14232 30880 14260
rect 29972 14220 29978 14232
rect 33042 14220 33048 14272
rect 33100 14220 33106 14272
rect 36633 14263 36691 14269
rect 36633 14229 36645 14263
rect 36679 14260 36691 14263
rect 37642 14260 37648 14272
rect 36679 14232 37648 14260
rect 36679 14229 36691 14232
rect 36633 14223 36691 14229
rect 37642 14220 37648 14232
rect 37700 14220 37706 14272
rect 40678 14220 40684 14272
rect 40736 14260 40742 14272
rect 44266 14260 44272 14272
rect 40736 14232 44272 14260
rect 40736 14220 40742 14232
rect 44266 14220 44272 14232
rect 44324 14220 44330 14272
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 2406 14056 2412 14068
rect 2367 14028 2412 14056
rect 2406 14016 2412 14028
rect 2464 14016 2470 14068
rect 14366 14016 14372 14068
rect 14424 14056 14430 14068
rect 14553 14059 14611 14065
rect 14553 14056 14565 14059
rect 14424 14028 14565 14056
rect 14424 14016 14430 14028
rect 14553 14025 14565 14028
rect 14599 14025 14611 14059
rect 14553 14019 14611 14025
rect 19426 14016 19432 14068
rect 19484 14056 19490 14068
rect 19521 14059 19579 14065
rect 19521 14056 19533 14059
rect 19484 14028 19533 14056
rect 19484 14016 19490 14028
rect 19521 14025 19533 14028
rect 19567 14025 19579 14059
rect 20070 14056 20076 14068
rect 19521 14019 19579 14025
rect 19904 14028 20076 14056
rect 19904 14000 19932 14028
rect 20070 14016 20076 14028
rect 20128 14016 20134 14068
rect 21174 14016 21180 14068
rect 21232 14056 21238 14068
rect 25774 14056 25780 14068
rect 21232 14028 23612 14056
rect 25735 14028 25780 14056
rect 21232 14016 21238 14028
rect 16206 13988 16212 14000
rect 13188 13960 16212 13988
rect 2498 13920 2504 13932
rect 2459 13892 2504 13920
rect 2498 13880 2504 13892
rect 2556 13920 2562 13932
rect 5166 13920 5172 13932
rect 2556 13892 5172 13920
rect 2556 13880 2562 13892
rect 5166 13880 5172 13892
rect 5224 13880 5230 13932
rect 12250 13880 12256 13932
rect 12308 13920 12314 13932
rect 13188 13929 13216 13960
rect 16206 13948 16212 13960
rect 16264 13948 16270 14000
rect 19886 13988 19892 14000
rect 19444 13960 19892 13988
rect 13446 13929 13452 13932
rect 13173 13923 13231 13929
rect 13173 13920 13185 13923
rect 12308 13892 13185 13920
rect 12308 13880 12314 13892
rect 13173 13889 13185 13892
rect 13219 13889 13231 13923
rect 13440 13920 13452 13929
rect 13407 13892 13452 13920
rect 13173 13883 13231 13889
rect 13440 13883 13452 13892
rect 13446 13880 13452 13883
rect 13504 13880 13510 13932
rect 19444 13929 19472 13960
rect 19886 13948 19892 13960
rect 19944 13948 19950 14000
rect 20622 13988 20628 14000
rect 20088 13960 20628 13988
rect 19429 13923 19487 13929
rect 19429 13889 19441 13923
rect 19475 13889 19487 13923
rect 19429 13883 19487 13889
rect 19613 13923 19671 13929
rect 19613 13889 19625 13923
rect 19659 13920 19671 13923
rect 19978 13920 19984 13932
rect 19659 13892 19984 13920
rect 19659 13889 19671 13892
rect 19613 13883 19671 13889
rect 19978 13880 19984 13892
rect 20036 13880 20042 13932
rect 19334 13812 19340 13864
rect 19392 13852 19398 13864
rect 20088 13861 20116 13960
rect 20622 13948 20628 13960
rect 20680 13988 20686 14000
rect 22646 13988 22652 14000
rect 20680 13960 22652 13988
rect 20680 13948 20686 13960
rect 22646 13948 22652 13960
rect 22704 13948 22710 14000
rect 20340 13923 20398 13929
rect 20340 13889 20352 13923
rect 20386 13920 20398 13923
rect 20898 13920 20904 13932
rect 20386 13892 20904 13920
rect 20386 13889 20398 13892
rect 20340 13883 20398 13889
rect 20898 13880 20904 13892
rect 20956 13880 20962 13932
rect 23382 13920 23388 13932
rect 23343 13892 23388 13920
rect 23382 13880 23388 13892
rect 23440 13880 23446 13932
rect 23584 13929 23612 14028
rect 25774 14016 25780 14028
rect 25832 14016 25838 14068
rect 33229 14059 33287 14065
rect 33229 14025 33241 14059
rect 33275 14056 33287 14059
rect 34974 14056 34980 14068
rect 33275 14028 34980 14056
rect 33275 14025 33287 14028
rect 33229 14019 33287 14025
rect 34974 14016 34980 14028
rect 35032 14016 35038 14068
rect 40494 14056 40500 14068
rect 40455 14028 40500 14056
rect 40494 14016 40500 14028
rect 40552 14016 40558 14068
rect 25498 13948 25504 14000
rect 25556 13988 25562 14000
rect 34146 13988 34152 14000
rect 25556 13960 26464 13988
rect 34107 13960 34152 13988
rect 25556 13948 25562 13960
rect 23569 13923 23627 13929
rect 23569 13889 23581 13923
rect 23615 13920 23627 13923
rect 23615 13892 25360 13920
rect 23615 13889 23627 13892
rect 23569 13883 23627 13889
rect 20073 13855 20131 13861
rect 20073 13852 20085 13855
rect 19392 13824 20085 13852
rect 19392 13812 19398 13824
rect 20073 13821 20085 13824
rect 20119 13821 20131 13855
rect 23658 13852 23664 13864
rect 23619 13824 23664 13852
rect 20073 13815 20131 13821
rect 23658 13812 23664 13824
rect 23716 13812 23722 13864
rect 25332 13852 25360 13892
rect 25682 13880 25688 13932
rect 25740 13920 25746 13932
rect 25961 13923 26019 13929
rect 25961 13920 25973 13923
rect 25740 13892 25973 13920
rect 25740 13880 25746 13892
rect 25961 13889 25973 13892
rect 26007 13889 26019 13923
rect 26234 13920 26240 13932
rect 26195 13892 26240 13920
rect 25961 13883 26019 13889
rect 26234 13880 26240 13892
rect 26292 13880 26298 13932
rect 26436 13929 26464 13960
rect 34146 13948 34152 13960
rect 34204 13948 34210 14000
rect 35897 13991 35955 13997
rect 35897 13957 35909 13991
rect 35943 13988 35955 13991
rect 36170 13988 36176 14000
rect 35943 13960 36176 13988
rect 35943 13957 35955 13960
rect 35897 13951 35955 13957
rect 36170 13948 36176 13960
rect 36228 13948 36234 14000
rect 40862 13988 40868 14000
rect 40823 13960 40868 13988
rect 40862 13948 40868 13960
rect 40920 13948 40926 14000
rect 26421 13923 26479 13929
rect 26421 13889 26433 13923
rect 26467 13889 26479 13923
rect 30006 13920 30012 13932
rect 29967 13892 30012 13920
rect 26421 13883 26479 13889
rect 30006 13880 30012 13892
rect 30064 13880 30070 13932
rect 30190 13920 30196 13932
rect 30151 13892 30196 13920
rect 30190 13880 30196 13892
rect 30248 13880 30254 13932
rect 33042 13920 33048 13932
rect 33003 13892 33048 13920
rect 33042 13880 33048 13892
rect 33100 13880 33106 13932
rect 33229 13923 33287 13929
rect 33229 13889 33241 13923
rect 33275 13920 33287 13923
rect 33410 13920 33416 13932
rect 33275 13892 33416 13920
rect 33275 13889 33287 13892
rect 33229 13883 33287 13889
rect 33410 13880 33416 13892
rect 33468 13880 33474 13932
rect 33778 13920 33784 13932
rect 33739 13892 33784 13920
rect 33778 13880 33784 13892
rect 33836 13880 33842 13932
rect 40678 13920 40684 13932
rect 40639 13892 40684 13920
rect 40678 13880 40684 13892
rect 40736 13880 40742 13932
rect 40773 13923 40831 13929
rect 40773 13889 40785 13923
rect 40819 13920 40831 13923
rect 40954 13920 40960 13932
rect 40819 13892 40960 13920
rect 40819 13889 40831 13892
rect 40773 13883 40831 13889
rect 40954 13880 40960 13892
rect 41012 13880 41018 13932
rect 41049 13923 41107 13929
rect 41049 13889 41061 13923
rect 41095 13920 41107 13923
rect 42978 13920 42984 13932
rect 41095 13892 42984 13920
rect 41095 13889 41107 13892
rect 41049 13883 41107 13889
rect 42978 13880 42984 13892
rect 43036 13880 43042 13932
rect 26694 13852 26700 13864
rect 25332 13824 26700 13852
rect 26694 13812 26700 13824
rect 26752 13812 26758 13864
rect 29917 13855 29975 13861
rect 29917 13821 29929 13855
rect 29963 13852 29975 13855
rect 30558 13852 30564 13864
rect 29963 13824 30564 13852
rect 29963 13821 29975 13824
rect 29917 13815 29975 13821
rect 30558 13812 30564 13824
rect 30616 13812 30622 13864
rect 47949 13855 48007 13861
rect 47949 13821 47961 13855
rect 47995 13852 48007 13855
rect 48314 13852 48320 13864
rect 47995 13824 48320 13852
rect 47995 13821 48007 13824
rect 47949 13815 48007 13821
rect 48314 13812 48320 13824
rect 48372 13812 48378 13864
rect 34974 13744 34980 13796
rect 35032 13784 35038 13796
rect 35802 13784 35808 13796
rect 35032 13756 35808 13784
rect 35032 13744 35038 13756
rect 35802 13744 35808 13756
rect 35860 13784 35866 13796
rect 36173 13787 36231 13793
rect 36173 13784 36185 13787
rect 35860 13756 36185 13784
rect 35860 13744 35866 13756
rect 36173 13753 36185 13756
rect 36219 13753 36231 13787
rect 36173 13747 36231 13753
rect 21453 13719 21511 13725
rect 21453 13685 21465 13719
rect 21499 13716 21511 13719
rect 21634 13716 21640 13728
rect 21499 13688 21640 13716
rect 21499 13685 21511 13688
rect 21453 13679 21511 13685
rect 21634 13676 21640 13688
rect 21692 13676 21698 13728
rect 23198 13716 23204 13728
rect 23159 13688 23204 13716
rect 23198 13676 23204 13688
rect 23256 13676 23262 13728
rect 30374 13716 30380 13728
rect 30335 13688 30380 13716
rect 30374 13676 30380 13688
rect 30432 13676 30438 13728
rect 36354 13716 36360 13728
rect 36315 13688 36360 13716
rect 36354 13676 36360 13688
rect 36412 13676 36418 13728
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 20993 13515 21051 13521
rect 20993 13481 21005 13515
rect 21039 13512 21051 13515
rect 21082 13512 21088 13524
rect 21039 13484 21088 13512
rect 21039 13481 21051 13484
rect 20993 13475 21051 13481
rect 21082 13472 21088 13484
rect 21140 13472 21146 13524
rect 26602 13472 26608 13524
rect 26660 13512 26666 13524
rect 27338 13512 27344 13524
rect 26660 13484 27344 13512
rect 26660 13472 26666 13484
rect 27338 13472 27344 13484
rect 27396 13472 27402 13524
rect 28537 13515 28595 13521
rect 28537 13481 28549 13515
rect 28583 13512 28595 13515
rect 30006 13512 30012 13524
rect 28583 13484 30012 13512
rect 28583 13481 28595 13484
rect 28537 13475 28595 13481
rect 30006 13472 30012 13484
rect 30064 13472 30070 13524
rect 32677 13515 32735 13521
rect 32677 13481 32689 13515
rect 32723 13512 32735 13515
rect 33410 13512 33416 13524
rect 32723 13484 33416 13512
rect 32723 13481 32735 13484
rect 32677 13475 32735 13481
rect 33410 13472 33416 13484
rect 33468 13472 33474 13524
rect 36265 13515 36323 13521
rect 36265 13481 36277 13515
rect 36311 13512 36323 13515
rect 36906 13512 36912 13524
rect 36311 13484 36912 13512
rect 36311 13481 36323 13484
rect 36265 13475 36323 13481
rect 36906 13472 36912 13484
rect 36964 13472 36970 13524
rect 19978 13404 19984 13456
rect 20036 13444 20042 13456
rect 20165 13447 20223 13453
rect 20165 13444 20177 13447
rect 20036 13416 20177 13444
rect 20036 13404 20042 13416
rect 20165 13413 20177 13416
rect 20211 13413 20223 13447
rect 20165 13407 20223 13413
rect 30466 13404 30472 13456
rect 30524 13444 30530 13456
rect 30742 13444 30748 13456
rect 30524 13416 30748 13444
rect 30524 13404 30530 13416
rect 30742 13404 30748 13416
rect 30800 13444 30806 13456
rect 31018 13444 31024 13456
rect 30800 13416 31024 13444
rect 30800 13404 30806 13416
rect 31018 13404 31024 13416
rect 31076 13404 31082 13456
rect 33318 13404 33324 13456
rect 33376 13444 33382 13456
rect 37182 13444 37188 13456
rect 33376 13416 37188 13444
rect 33376 13404 33382 13416
rect 37182 13404 37188 13416
rect 37240 13404 37246 13456
rect 18322 13336 18328 13388
rect 18380 13336 18386 13388
rect 22646 13376 22652 13388
rect 22607 13348 22652 13376
rect 22646 13336 22652 13348
rect 22704 13336 22710 13388
rect 27614 13376 27620 13388
rect 23768 13348 27620 13376
rect 16206 13308 16212 13320
rect 16167 13280 16212 13308
rect 16206 13268 16212 13280
rect 16264 13268 16270 13320
rect 18233 13311 18291 13317
rect 18233 13277 18245 13311
rect 18279 13308 18291 13311
rect 18340 13308 18368 13336
rect 18506 13308 18512 13320
rect 18279 13280 18368 13308
rect 18467 13280 18512 13308
rect 18279 13277 18291 13280
rect 18233 13271 18291 13277
rect 18506 13268 18512 13280
rect 18564 13268 18570 13320
rect 18693 13311 18751 13317
rect 18693 13277 18705 13311
rect 18739 13277 18751 13311
rect 19886 13308 19892 13320
rect 19847 13280 19892 13308
rect 18693 13271 18751 13277
rect 16476 13243 16534 13249
rect 16476 13209 16488 13243
rect 16522 13240 16534 13243
rect 17034 13240 17040 13252
rect 16522 13212 17040 13240
rect 16522 13209 16534 13212
rect 16476 13203 16534 13209
rect 17034 13200 17040 13212
rect 17092 13200 17098 13252
rect 18322 13240 18328 13252
rect 17604 13212 18328 13240
rect 17604 13181 17632 13212
rect 18322 13200 18328 13212
rect 18380 13240 18386 13252
rect 18708 13240 18736 13271
rect 19886 13268 19892 13280
rect 19944 13268 19950 13320
rect 19981 13311 20039 13317
rect 19981 13277 19993 13311
rect 20027 13308 20039 13311
rect 20070 13308 20076 13320
rect 20027 13280 20076 13308
rect 20027 13277 20039 13280
rect 19981 13271 20039 13277
rect 20070 13268 20076 13280
rect 20128 13268 20134 13320
rect 20165 13311 20223 13317
rect 20165 13277 20177 13311
rect 20211 13308 20223 13311
rect 20254 13308 20260 13320
rect 20211 13280 20260 13308
rect 20211 13277 20223 13280
rect 20165 13271 20223 13277
rect 20254 13268 20260 13280
rect 20312 13268 20318 13320
rect 21174 13308 21180 13320
rect 21135 13280 21180 13308
rect 21174 13268 21180 13280
rect 21232 13268 21238 13320
rect 21453 13311 21511 13317
rect 21453 13277 21465 13311
rect 21499 13277 21511 13311
rect 21634 13308 21640 13320
rect 21595 13280 21640 13308
rect 21453 13271 21511 13277
rect 18380 13212 18736 13240
rect 21468 13240 21496 13271
rect 21634 13268 21640 13280
rect 21692 13268 21698 13320
rect 22916 13311 22974 13317
rect 22916 13277 22928 13311
rect 22962 13308 22974 13311
rect 23198 13308 23204 13320
rect 22962 13280 23204 13308
rect 22962 13277 22974 13280
rect 22916 13271 22974 13277
rect 23198 13268 23204 13280
rect 23256 13268 23262 13320
rect 23768 13252 23796 13348
rect 26050 13308 26056 13320
rect 26011 13280 26056 13308
rect 26050 13268 26056 13280
rect 26108 13268 26114 13320
rect 26252 13317 26280 13348
rect 27614 13336 27620 13348
rect 27672 13336 27678 13388
rect 28718 13336 28724 13388
rect 28776 13376 28782 13388
rect 30006 13376 30012 13388
rect 28776 13348 30012 13376
rect 28776 13336 28782 13348
rect 30006 13336 30012 13348
rect 30064 13376 30070 13388
rect 31297 13379 31355 13385
rect 31297 13376 31309 13379
rect 30064 13348 31309 13376
rect 30064 13336 30070 13348
rect 31297 13345 31309 13348
rect 31343 13345 31355 13379
rect 31297 13339 31355 13345
rect 33134 13336 33140 13388
rect 33192 13376 33198 13388
rect 33505 13379 33563 13385
rect 33505 13376 33517 13379
rect 33192 13348 33517 13376
rect 33192 13336 33198 13348
rect 33505 13345 33517 13348
rect 33551 13345 33563 13379
rect 33505 13339 33563 13345
rect 36357 13379 36415 13385
rect 36357 13345 36369 13379
rect 36403 13376 36415 13379
rect 36446 13376 36452 13388
rect 36403 13348 36452 13376
rect 36403 13345 36415 13348
rect 36357 13339 36415 13345
rect 36446 13336 36452 13348
rect 36504 13336 36510 13388
rect 37642 13376 37648 13388
rect 37603 13348 37648 13376
rect 37642 13336 37648 13348
rect 37700 13336 37706 13388
rect 37737 13379 37795 13385
rect 37737 13345 37749 13379
rect 37783 13376 37795 13379
rect 38470 13376 38476 13388
rect 37783 13348 38476 13376
rect 37783 13345 37795 13348
rect 37737 13339 37795 13345
rect 38470 13336 38476 13348
rect 38528 13336 38534 13388
rect 46842 13376 46848 13388
rect 46803 13348 46848 13376
rect 46842 13336 46848 13348
rect 46900 13336 46906 13388
rect 48314 13376 48320 13388
rect 48275 13348 48320 13376
rect 48314 13336 48320 13348
rect 48372 13336 48378 13388
rect 26237 13311 26295 13317
rect 26237 13277 26249 13311
rect 26283 13277 26295 13311
rect 26237 13271 26295 13277
rect 26513 13311 26571 13317
rect 26513 13277 26525 13311
rect 26559 13308 26571 13311
rect 26602 13308 26608 13320
rect 26559 13280 26608 13308
rect 26559 13277 26571 13280
rect 26513 13271 26571 13277
rect 26602 13268 26608 13280
rect 26660 13268 26666 13320
rect 27157 13311 27215 13317
rect 27157 13277 27169 13311
rect 27203 13277 27215 13311
rect 28350 13308 28356 13320
rect 28311 13280 28356 13308
rect 27157 13271 27215 13277
rect 22094 13240 22100 13252
rect 21468 13212 22100 13240
rect 18380 13200 18386 13212
rect 22094 13200 22100 13212
rect 22152 13240 22158 13252
rect 23750 13240 23756 13252
rect 22152 13212 23756 13240
rect 22152 13200 22158 13212
rect 23750 13200 23756 13212
rect 23808 13200 23814 13252
rect 25866 13200 25872 13252
rect 25924 13240 25930 13252
rect 27172 13240 27200 13271
rect 28350 13268 28356 13280
rect 28408 13268 28414 13320
rect 28626 13268 28632 13320
rect 28684 13308 28690 13320
rect 29914 13308 29920 13320
rect 28684 13280 28729 13308
rect 29875 13280 29920 13308
rect 28684 13268 28690 13280
rect 29914 13268 29920 13280
rect 29972 13268 29978 13320
rect 30101 13311 30159 13317
rect 30101 13277 30113 13311
rect 30147 13277 30159 13311
rect 30101 13271 30159 13277
rect 30377 13311 30435 13317
rect 30377 13277 30389 13311
rect 30423 13308 30435 13311
rect 30466 13308 30472 13320
rect 30423 13280 30472 13308
rect 30423 13277 30435 13280
rect 30377 13271 30435 13277
rect 28534 13240 28540 13252
rect 25924 13212 28540 13240
rect 25924 13200 25930 13212
rect 28534 13200 28540 13212
rect 28592 13200 28598 13252
rect 29638 13200 29644 13252
rect 29696 13240 29702 13252
rect 30116 13240 30144 13271
rect 30466 13268 30472 13280
rect 30524 13268 30530 13320
rect 30561 13311 30619 13317
rect 30561 13277 30573 13311
rect 30607 13308 30619 13311
rect 33321 13311 33379 13317
rect 33321 13308 33333 13311
rect 30607 13280 33333 13308
rect 30607 13277 30619 13280
rect 30561 13271 30619 13277
rect 33321 13277 33333 13280
rect 33367 13277 33379 13311
rect 33321 13271 33379 13277
rect 33410 13268 33416 13320
rect 33468 13308 33474 13320
rect 33597 13311 33655 13317
rect 33597 13308 33609 13311
rect 33468 13280 33609 13308
rect 33468 13268 33474 13280
rect 33597 13277 33609 13280
rect 33643 13277 33655 13311
rect 33597 13271 33655 13277
rect 35802 13268 35808 13320
rect 35860 13308 35866 13320
rect 35989 13311 36047 13317
rect 35989 13308 36001 13311
rect 35860 13280 36001 13308
rect 35860 13268 35866 13280
rect 35989 13277 36001 13280
rect 36035 13277 36047 13311
rect 35989 13271 36047 13277
rect 36722 13268 36728 13320
rect 36780 13308 36786 13320
rect 37553 13311 37611 13317
rect 37553 13308 37565 13311
rect 36780 13280 37565 13308
rect 36780 13268 36786 13280
rect 37553 13277 37565 13280
rect 37599 13277 37611 13311
rect 37553 13271 37611 13277
rect 37826 13268 37832 13320
rect 37884 13308 37890 13320
rect 37884 13280 37929 13308
rect 37884 13268 37890 13280
rect 30650 13240 30656 13252
rect 29696 13212 30656 13240
rect 29696 13200 29702 13212
rect 30650 13200 30656 13212
rect 30708 13200 30714 13252
rect 31564 13243 31622 13249
rect 31564 13209 31576 13243
rect 31610 13240 31622 13243
rect 33137 13243 33195 13249
rect 33137 13240 33149 13243
rect 31610 13212 33149 13240
rect 31610 13209 31622 13212
rect 31564 13203 31622 13209
rect 33137 13209 33149 13212
rect 33183 13209 33195 13243
rect 33137 13203 33195 13209
rect 36170 13200 36176 13252
rect 36228 13240 36234 13252
rect 36449 13243 36507 13249
rect 36449 13240 36461 13243
rect 36228 13212 36461 13240
rect 36228 13200 36234 13212
rect 36449 13209 36461 13212
rect 36495 13209 36507 13243
rect 36449 13203 36507 13209
rect 47854 13200 47860 13252
rect 47912 13240 47918 13252
rect 48133 13243 48191 13249
rect 48133 13240 48145 13243
rect 47912 13212 48145 13240
rect 47912 13200 47918 13212
rect 48133 13209 48145 13212
rect 48179 13209 48191 13243
rect 48133 13203 48191 13209
rect 17589 13175 17647 13181
rect 17589 13141 17601 13175
rect 17635 13141 17647 13175
rect 18046 13172 18052 13184
rect 18007 13144 18052 13172
rect 17589 13135 17647 13141
rect 18046 13132 18052 13144
rect 18104 13132 18110 13184
rect 24026 13172 24032 13184
rect 23987 13144 24032 13172
rect 24026 13132 24032 13144
rect 24084 13132 24090 13184
rect 26418 13132 26424 13184
rect 26476 13172 26482 13184
rect 26697 13175 26755 13181
rect 26697 13172 26709 13175
rect 26476 13144 26709 13172
rect 26476 13132 26482 13144
rect 26697 13141 26709 13144
rect 26743 13141 26755 13175
rect 26697 13135 26755 13141
rect 27982 13132 27988 13184
rect 28040 13172 28046 13184
rect 28169 13175 28227 13181
rect 28169 13172 28181 13175
rect 28040 13144 28181 13172
rect 28040 13132 28046 13144
rect 28169 13141 28181 13144
rect 28215 13141 28227 13175
rect 28169 13135 28227 13141
rect 36081 13175 36139 13181
rect 36081 13141 36093 13175
rect 36127 13172 36139 13175
rect 36814 13172 36820 13184
rect 36127 13144 36820 13172
rect 36127 13141 36139 13144
rect 36081 13135 36139 13141
rect 36814 13132 36820 13144
rect 36872 13132 36878 13184
rect 37366 13172 37372 13184
rect 37327 13144 37372 13172
rect 37366 13132 37372 13144
rect 37424 13132 37430 13184
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 17034 12968 17040 12980
rect 16995 12940 17040 12968
rect 17034 12928 17040 12940
rect 17092 12928 17098 12980
rect 20441 12971 20499 12977
rect 20441 12937 20453 12971
rect 20487 12968 20499 12971
rect 21634 12968 21640 12980
rect 20487 12940 21640 12968
rect 20487 12937 20499 12940
rect 20441 12931 20499 12937
rect 21634 12928 21640 12940
rect 21692 12928 21698 12980
rect 23293 12971 23351 12977
rect 23293 12937 23305 12971
rect 23339 12968 23351 12971
rect 23382 12968 23388 12980
rect 23339 12940 23388 12968
rect 23339 12937 23351 12940
rect 23293 12931 23351 12937
rect 23382 12928 23388 12940
rect 23440 12928 23446 12980
rect 25225 12971 25283 12977
rect 25225 12937 25237 12971
rect 25271 12968 25283 12971
rect 25314 12968 25320 12980
rect 25271 12940 25320 12968
rect 25271 12937 25283 12940
rect 25225 12931 25283 12937
rect 25314 12928 25320 12940
rect 25372 12968 25378 12980
rect 26050 12968 26056 12980
rect 25372 12940 26056 12968
rect 25372 12928 25378 12940
rect 26050 12928 26056 12940
rect 26108 12928 26114 12980
rect 26602 12928 26608 12980
rect 26660 12928 26666 12980
rect 33597 12971 33655 12977
rect 33597 12937 33609 12971
rect 33643 12968 33655 12971
rect 33778 12968 33784 12980
rect 33643 12940 33784 12968
rect 33643 12937 33655 12940
rect 33597 12931 33655 12937
rect 33778 12928 33784 12940
rect 33836 12928 33842 12980
rect 35529 12971 35587 12977
rect 35529 12937 35541 12971
rect 35575 12937 35587 12971
rect 36722 12968 36728 12980
rect 36683 12940 36728 12968
rect 35529 12931 35587 12937
rect 21358 12900 21364 12912
rect 20180 12872 21364 12900
rect 17221 12835 17279 12841
rect 17221 12801 17233 12835
rect 17267 12832 17279 12835
rect 18046 12832 18052 12844
rect 17267 12804 18052 12832
rect 17267 12801 17279 12804
rect 17221 12795 17279 12801
rect 18046 12792 18052 12804
rect 18104 12792 18110 12844
rect 4706 12724 4712 12776
rect 4764 12764 4770 12776
rect 17497 12767 17555 12773
rect 17497 12764 17509 12767
rect 4764 12736 17509 12764
rect 4764 12724 4770 12736
rect 17497 12733 17509 12736
rect 17543 12764 17555 12767
rect 20180 12764 20208 12872
rect 21358 12860 21364 12872
rect 21416 12860 21422 12912
rect 26620 12900 26648 12928
rect 28718 12900 28724 12912
rect 23492 12872 26648 12900
rect 27724 12872 28724 12900
rect 20438 12792 20444 12844
rect 20496 12832 20502 12844
rect 20496 12804 20668 12832
rect 20496 12792 20502 12804
rect 17543 12736 20208 12764
rect 17543 12733 17555 12736
rect 17497 12727 17555 12733
rect 20254 12724 20260 12776
rect 20312 12764 20318 12776
rect 20640 12773 20668 12804
rect 21174 12792 21180 12844
rect 21232 12832 21238 12844
rect 23492 12841 23520 12872
rect 23477 12835 23535 12841
rect 23477 12832 23489 12835
rect 21232 12804 23489 12832
rect 21232 12792 21238 12804
rect 23477 12801 23489 12804
rect 23523 12801 23535 12835
rect 23750 12832 23756 12844
rect 23711 12804 23756 12832
rect 23477 12795 23535 12801
rect 23750 12792 23756 12804
rect 23808 12792 23814 12844
rect 23937 12835 23995 12841
rect 23937 12801 23949 12835
rect 23983 12832 23995 12835
rect 24026 12832 24032 12844
rect 23983 12804 24032 12832
rect 23983 12801 23995 12804
rect 23937 12795 23995 12801
rect 24026 12792 24032 12804
rect 24084 12792 24090 12844
rect 26326 12832 26332 12844
rect 26384 12841 26390 12844
rect 27724 12841 27752 12872
rect 28718 12860 28724 12872
rect 28776 12860 28782 12912
rect 30276 12903 30334 12909
rect 30276 12869 30288 12903
rect 30322 12900 30334 12903
rect 30374 12900 30380 12912
rect 30322 12872 30380 12900
rect 30322 12869 30334 12872
rect 30276 12863 30334 12869
rect 30374 12860 30380 12872
rect 30432 12860 30438 12912
rect 33318 12860 33324 12912
rect 33376 12900 33382 12912
rect 33413 12903 33471 12909
rect 33413 12900 33425 12903
rect 33376 12872 33425 12900
rect 33376 12860 33382 12872
rect 33413 12869 33425 12872
rect 33459 12869 33471 12903
rect 35544 12900 35572 12931
rect 36722 12928 36728 12940
rect 36780 12968 36786 12980
rect 36998 12968 37004 12980
rect 36780 12940 37004 12968
rect 36780 12928 36786 12940
rect 36998 12928 37004 12940
rect 37056 12928 37062 12980
rect 42334 12968 42340 12980
rect 37292 12940 42340 12968
rect 37292 12900 37320 12940
rect 42334 12928 42340 12940
rect 42392 12928 42398 12980
rect 47854 12968 47860 12980
rect 47815 12940 47860 12968
rect 47854 12928 47860 12940
rect 47912 12928 47918 12980
rect 35544 12872 37320 12900
rect 33413 12863 33471 12869
rect 37366 12860 37372 12912
rect 37424 12900 37430 12912
rect 38758 12903 38816 12909
rect 38758 12900 38770 12903
rect 37424 12872 38770 12900
rect 37424 12860 37430 12872
rect 38758 12869 38770 12872
rect 38804 12869 38816 12903
rect 38758 12863 38816 12869
rect 27982 12841 27988 12844
rect 26296 12804 26332 12832
rect 26326 12792 26332 12804
rect 26384 12795 26396 12841
rect 26605 12835 26663 12841
rect 26605 12801 26617 12835
rect 26651 12832 26663 12835
rect 27709 12835 27767 12841
rect 27709 12832 27721 12835
rect 26651 12804 27721 12832
rect 26651 12801 26663 12804
rect 26605 12795 26663 12801
rect 27709 12801 27721 12804
rect 27755 12801 27767 12835
rect 27976 12832 27988 12841
rect 27943 12804 27988 12832
rect 27709 12795 27767 12801
rect 27976 12795 27988 12804
rect 26384 12792 26390 12795
rect 27982 12792 27988 12795
rect 28040 12792 28046 12844
rect 29822 12792 29828 12844
rect 29880 12832 29886 12844
rect 30006 12832 30012 12844
rect 29880 12804 30012 12832
rect 29880 12792 29886 12804
rect 30006 12792 30012 12804
rect 30064 12792 30070 12844
rect 33226 12832 33232 12844
rect 33139 12804 33232 12832
rect 33226 12792 33232 12804
rect 33284 12832 33290 12844
rect 33284 12804 33456 12832
rect 33284 12792 33290 12804
rect 20533 12767 20591 12773
rect 20533 12764 20545 12767
rect 20312 12736 20545 12764
rect 20312 12724 20318 12736
rect 20533 12733 20545 12736
rect 20579 12733 20591 12767
rect 20533 12727 20591 12733
rect 20625 12767 20683 12773
rect 20625 12733 20637 12767
rect 20671 12764 20683 12767
rect 23290 12764 23296 12776
rect 20671 12736 23296 12764
rect 20671 12733 20683 12736
rect 20625 12727 20683 12733
rect 23290 12724 23296 12736
rect 23348 12724 23354 12776
rect 17405 12699 17463 12705
rect 17405 12665 17417 12699
rect 17451 12696 17463 12699
rect 18230 12696 18236 12708
rect 17451 12668 18236 12696
rect 17451 12665 17463 12668
rect 17405 12659 17463 12665
rect 18230 12656 18236 12668
rect 18288 12656 18294 12708
rect 33428 12696 33456 12804
rect 34606 12792 34612 12844
rect 34664 12832 34670 12844
rect 34885 12835 34943 12841
rect 34885 12832 34897 12835
rect 34664 12804 34897 12832
rect 34664 12792 34670 12804
rect 34885 12801 34897 12804
rect 34931 12801 34943 12835
rect 34885 12795 34943 12801
rect 35069 12835 35127 12841
rect 35069 12801 35081 12835
rect 35115 12832 35127 12835
rect 35713 12835 35771 12841
rect 35713 12832 35725 12835
rect 35115 12804 35725 12832
rect 35115 12801 35127 12804
rect 35069 12795 35127 12801
rect 35713 12801 35725 12804
rect 35759 12801 35771 12835
rect 35713 12795 35771 12801
rect 35897 12835 35955 12841
rect 35897 12801 35909 12835
rect 35943 12801 35955 12835
rect 35897 12795 35955 12801
rect 36357 12835 36415 12841
rect 36357 12801 36369 12835
rect 36403 12832 36415 12835
rect 36630 12832 36636 12844
rect 36403 12804 36636 12832
rect 36403 12801 36415 12804
rect 36357 12795 36415 12801
rect 34790 12724 34796 12776
rect 34848 12764 34854 12776
rect 35084 12764 35112 12795
rect 34848 12736 35112 12764
rect 34848 12724 34854 12736
rect 35802 12696 35808 12708
rect 33428 12668 35808 12696
rect 35802 12656 35808 12668
rect 35860 12656 35866 12708
rect 35912 12696 35940 12795
rect 36630 12792 36636 12804
rect 36688 12792 36694 12844
rect 39025 12835 39083 12841
rect 39025 12801 39037 12835
rect 39071 12832 39083 12835
rect 40218 12832 40224 12844
rect 39071 12804 40224 12832
rect 39071 12801 39083 12804
rect 39025 12795 39083 12801
rect 40218 12792 40224 12804
rect 40276 12792 40282 12844
rect 46385 12835 46443 12841
rect 46385 12801 46397 12835
rect 46431 12832 46443 12835
rect 46750 12832 46756 12844
rect 46431 12804 46756 12832
rect 46431 12801 46443 12804
rect 46385 12795 46443 12801
rect 46750 12792 46756 12804
rect 46808 12792 46814 12844
rect 47486 12792 47492 12844
rect 47544 12832 47550 12844
rect 47670 12832 47676 12844
rect 47544 12804 47676 12832
rect 47544 12792 47550 12804
rect 47670 12792 47676 12804
rect 47728 12832 47734 12844
rect 47765 12835 47823 12841
rect 47765 12832 47777 12835
rect 47728 12804 47777 12832
rect 47728 12792 47734 12804
rect 47765 12801 47777 12804
rect 47811 12801 47823 12835
rect 47765 12795 47823 12801
rect 36446 12764 36452 12776
rect 36407 12736 36452 12764
rect 36446 12724 36452 12736
rect 36504 12724 36510 12776
rect 37550 12696 37556 12708
rect 35912 12668 37556 12696
rect 37550 12656 37556 12668
rect 37608 12656 37614 12708
rect 17954 12588 17960 12640
rect 18012 12628 18018 12640
rect 20073 12631 20131 12637
rect 20073 12628 20085 12631
rect 18012 12600 20085 12628
rect 18012 12588 18018 12600
rect 20073 12597 20085 12600
rect 20119 12597 20131 12631
rect 29086 12628 29092 12640
rect 29047 12600 29092 12628
rect 20073 12591 20131 12597
rect 29086 12588 29092 12600
rect 29144 12588 29150 12640
rect 31386 12628 31392 12640
rect 31347 12600 31392 12628
rect 31386 12588 31392 12600
rect 31444 12588 31450 12640
rect 35069 12631 35127 12637
rect 35069 12597 35081 12631
rect 35115 12628 35127 12631
rect 35434 12628 35440 12640
rect 35115 12600 35440 12628
rect 35115 12597 35127 12600
rect 35069 12591 35127 12597
rect 35434 12588 35440 12600
rect 35492 12588 35498 12640
rect 35897 12631 35955 12637
rect 35897 12597 35909 12631
rect 35943 12628 35955 12631
rect 36170 12628 36176 12640
rect 35943 12600 36176 12628
rect 35943 12597 35955 12600
rect 35897 12591 35955 12597
rect 36170 12588 36176 12600
rect 36228 12588 36234 12640
rect 36354 12628 36360 12640
rect 36315 12600 36360 12628
rect 36354 12588 36360 12600
rect 36412 12588 36418 12640
rect 37458 12588 37464 12640
rect 37516 12628 37522 12640
rect 37645 12631 37703 12637
rect 37645 12628 37657 12631
rect 37516 12600 37657 12628
rect 37516 12588 37522 12600
rect 37645 12597 37657 12600
rect 37691 12597 37703 12631
rect 37645 12591 37703 12597
rect 46477 12631 46535 12637
rect 46477 12597 46489 12631
rect 46523 12628 46535 12631
rect 46658 12628 46664 12640
rect 46523 12600 46664 12628
rect 46523 12597 46535 12600
rect 46477 12591 46535 12597
rect 46658 12588 46664 12600
rect 46716 12588 46722 12640
rect 47026 12628 47032 12640
rect 46987 12600 47032 12628
rect 47026 12588 47032 12600
rect 47084 12588 47090 12640
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 17494 12424 17500 12436
rect 17407 12396 17500 12424
rect 17420 12297 17448 12396
rect 17494 12384 17500 12396
rect 17552 12424 17558 12436
rect 20530 12424 20536 12436
rect 17552 12396 20536 12424
rect 17552 12384 17558 12396
rect 20530 12384 20536 12396
rect 20588 12384 20594 12436
rect 26145 12427 26203 12433
rect 26145 12393 26157 12427
rect 26191 12424 26203 12427
rect 26326 12424 26332 12436
rect 26191 12396 26332 12424
rect 26191 12393 26203 12396
rect 26145 12387 26203 12393
rect 26326 12384 26332 12396
rect 26384 12384 26390 12436
rect 26513 12427 26571 12433
rect 26513 12393 26525 12427
rect 26559 12424 26571 12427
rect 26602 12424 26608 12436
rect 26559 12396 26608 12424
rect 26559 12393 26571 12396
rect 26513 12387 26571 12393
rect 26602 12384 26608 12396
rect 26660 12384 26666 12436
rect 28350 12384 28356 12436
rect 28408 12424 28414 12436
rect 28445 12427 28503 12433
rect 28445 12424 28457 12427
rect 28408 12396 28457 12424
rect 28408 12384 28414 12396
rect 28445 12393 28457 12396
rect 28491 12393 28503 12427
rect 30190 12424 30196 12436
rect 30151 12396 30196 12424
rect 28445 12387 28503 12393
rect 30190 12384 30196 12396
rect 30248 12384 30254 12436
rect 34698 12384 34704 12436
rect 34756 12424 34762 12436
rect 34977 12427 35035 12433
rect 34977 12424 34989 12427
rect 34756 12396 34989 12424
rect 34756 12384 34762 12396
rect 34977 12393 34989 12396
rect 35023 12393 35035 12427
rect 34977 12387 35035 12393
rect 35894 12384 35900 12436
rect 35952 12424 35958 12436
rect 36354 12424 36360 12436
rect 35952 12396 36360 12424
rect 35952 12384 35958 12396
rect 36354 12384 36360 12396
rect 36412 12384 36418 12436
rect 37826 12384 37832 12436
rect 37884 12424 37890 12436
rect 38013 12427 38071 12433
rect 38013 12424 38025 12427
rect 37884 12396 38025 12424
rect 37884 12384 37890 12396
rect 38013 12393 38025 12396
rect 38059 12393 38071 12427
rect 38013 12387 38071 12393
rect 20254 12356 20260 12368
rect 20215 12328 20260 12356
rect 20254 12316 20260 12328
rect 20312 12316 20318 12368
rect 29086 12316 29092 12368
rect 29144 12356 29150 12368
rect 47026 12356 47032 12368
rect 29144 12328 37136 12356
rect 29144 12316 29150 12328
rect 17405 12291 17463 12297
rect 17405 12257 17417 12291
rect 17451 12257 17463 12291
rect 19978 12288 19984 12300
rect 19939 12260 19984 12288
rect 17405 12251 17463 12257
rect 19978 12248 19984 12260
rect 20036 12248 20042 12300
rect 23290 12248 23296 12300
rect 23348 12288 23354 12300
rect 23569 12291 23627 12297
rect 23569 12288 23581 12291
rect 23348 12260 23581 12288
rect 23348 12248 23354 12260
rect 23569 12257 23581 12260
rect 23615 12288 23627 12291
rect 23842 12288 23848 12300
rect 23615 12260 23848 12288
rect 23615 12257 23627 12260
rect 23569 12251 23627 12257
rect 23842 12248 23848 12260
rect 23900 12248 23906 12300
rect 26602 12288 26608 12300
rect 26515 12260 26608 12288
rect 26602 12248 26608 12260
rect 26660 12288 26666 12300
rect 30558 12288 30564 12300
rect 26660 12260 30564 12288
rect 26660 12248 26666 12260
rect 30558 12248 30564 12260
rect 30616 12248 30622 12300
rect 33778 12248 33784 12300
rect 33836 12288 33842 12300
rect 33965 12291 34023 12297
rect 33965 12288 33977 12291
rect 33836 12260 33977 12288
rect 33836 12248 33842 12260
rect 33965 12257 33977 12260
rect 34011 12257 34023 12291
rect 35897 12291 35955 12297
rect 35897 12288 35909 12291
rect 33965 12251 34023 12257
rect 35176 12260 35909 12288
rect 2409 12223 2467 12229
rect 2409 12189 2421 12223
rect 2455 12220 2467 12223
rect 2590 12220 2596 12232
rect 2455 12192 2596 12220
rect 2455 12189 2467 12192
rect 2409 12183 2467 12189
rect 2590 12180 2596 12192
rect 2648 12180 2654 12232
rect 17221 12223 17279 12229
rect 17221 12189 17233 12223
rect 17267 12220 17279 12223
rect 17954 12220 17960 12232
rect 17267 12192 17960 12220
rect 17267 12189 17279 12192
rect 17221 12183 17279 12189
rect 17954 12180 17960 12192
rect 18012 12180 18018 12232
rect 18049 12223 18107 12229
rect 18049 12189 18061 12223
rect 18095 12189 18107 12223
rect 18049 12183 18107 12189
rect 18233 12223 18291 12229
rect 18233 12189 18245 12223
rect 18279 12220 18291 12223
rect 18322 12220 18328 12232
rect 18279 12192 18328 12220
rect 18279 12189 18291 12192
rect 18233 12183 18291 12189
rect 18064 12152 18092 12183
rect 18322 12180 18328 12192
rect 18380 12220 18386 12232
rect 18693 12223 18751 12229
rect 18693 12220 18705 12223
rect 18380 12192 18705 12220
rect 18380 12180 18386 12192
rect 18693 12189 18705 12192
rect 18739 12189 18751 12223
rect 18693 12183 18751 12189
rect 18877 12223 18935 12229
rect 18877 12189 18889 12223
rect 18923 12189 18935 12223
rect 18877 12183 18935 12189
rect 19889 12223 19947 12229
rect 19889 12189 19901 12223
rect 19935 12220 19947 12223
rect 23385 12223 23443 12229
rect 19935 12192 20024 12220
rect 19935 12189 19947 12192
rect 19889 12183 19947 12189
rect 18892 12152 18920 12183
rect 19996 12164 20024 12192
rect 23385 12189 23397 12223
rect 23431 12220 23443 12223
rect 24026 12220 24032 12232
rect 23431 12192 24032 12220
rect 23431 12189 23443 12192
rect 23385 12183 23443 12189
rect 24026 12180 24032 12192
rect 24084 12180 24090 12232
rect 25409 12223 25467 12229
rect 25409 12189 25421 12223
rect 25455 12220 25467 12223
rect 25866 12220 25872 12232
rect 25455 12192 25872 12220
rect 25455 12189 25467 12192
rect 25409 12183 25467 12189
rect 25866 12180 25872 12192
rect 25924 12180 25930 12232
rect 26329 12223 26387 12229
rect 26329 12189 26341 12223
rect 26375 12220 26387 12223
rect 26418 12220 26424 12232
rect 26375 12192 26424 12220
rect 26375 12189 26387 12192
rect 26329 12183 26387 12189
rect 26418 12180 26424 12192
rect 26476 12180 26482 12232
rect 28629 12223 28687 12229
rect 28629 12189 28641 12223
rect 28675 12189 28687 12223
rect 28629 12183 28687 12189
rect 28905 12223 28963 12229
rect 28905 12189 28917 12223
rect 28951 12189 28963 12223
rect 29086 12220 29092 12232
rect 29047 12192 29092 12220
rect 28905 12183 28963 12189
rect 17328 12124 18920 12152
rect 17328 12096 17356 12124
rect 19978 12112 19984 12164
rect 20036 12112 20042 12164
rect 22922 12112 22928 12164
rect 22980 12152 22986 12164
rect 23477 12155 23535 12161
rect 23477 12152 23489 12155
rect 22980 12124 23489 12152
rect 22980 12112 22986 12124
rect 23477 12121 23489 12124
rect 23523 12121 23535 12155
rect 23477 12115 23535 12121
rect 2222 12044 2228 12096
rect 2280 12084 2286 12096
rect 2317 12087 2375 12093
rect 2317 12084 2329 12087
rect 2280 12056 2329 12084
rect 2280 12044 2286 12056
rect 2317 12053 2329 12056
rect 2363 12053 2375 12087
rect 2317 12047 2375 12053
rect 16853 12087 16911 12093
rect 16853 12053 16865 12087
rect 16899 12084 16911 12087
rect 17034 12084 17040 12096
rect 16899 12056 17040 12084
rect 16899 12053 16911 12056
rect 16853 12047 16911 12053
rect 17034 12044 17040 12056
rect 17092 12044 17098 12096
rect 17310 12084 17316 12096
rect 17271 12056 17316 12084
rect 17310 12044 17316 12056
rect 17368 12044 17374 12096
rect 18230 12084 18236 12096
rect 18191 12056 18236 12084
rect 18230 12044 18236 12056
rect 18288 12044 18294 12096
rect 18785 12087 18843 12093
rect 18785 12053 18797 12087
rect 18831 12084 18843 12087
rect 18966 12084 18972 12096
rect 18831 12056 18972 12084
rect 18831 12053 18843 12056
rect 18785 12047 18843 12053
rect 18966 12044 18972 12056
rect 19024 12044 19030 12096
rect 20806 12044 20812 12096
rect 20864 12084 20870 12096
rect 23017 12087 23075 12093
rect 23017 12084 23029 12087
rect 20864 12056 23029 12084
rect 20864 12044 20870 12056
rect 23017 12053 23029 12056
rect 23063 12053 23075 12087
rect 25590 12084 25596 12096
rect 25551 12056 25596 12084
rect 23017 12047 23075 12053
rect 25590 12044 25596 12056
rect 25648 12044 25654 12096
rect 28644 12084 28672 12183
rect 28920 12152 28948 12183
rect 29086 12180 29092 12192
rect 29144 12180 29150 12232
rect 30282 12180 30288 12232
rect 30340 12220 30346 12232
rect 30377 12223 30435 12229
rect 30377 12220 30389 12223
rect 30340 12192 30389 12220
rect 30340 12180 30346 12192
rect 30377 12189 30389 12192
rect 30423 12189 30435 12223
rect 30377 12183 30435 12189
rect 30653 12223 30711 12229
rect 30653 12189 30665 12223
rect 30699 12189 30711 12223
rect 30653 12183 30711 12189
rect 30837 12223 30895 12229
rect 30837 12189 30849 12223
rect 30883 12220 30895 12223
rect 31386 12220 31392 12232
rect 30883 12192 31392 12220
rect 30883 12189 30895 12192
rect 30837 12183 30895 12189
rect 30098 12152 30104 12164
rect 28920 12124 30104 12152
rect 30098 12112 30104 12124
rect 30156 12152 30162 12164
rect 30668 12152 30696 12183
rect 31386 12180 31392 12192
rect 31444 12220 31450 12232
rect 35176 12229 35204 12260
rect 35897 12257 35909 12260
rect 35943 12257 35955 12291
rect 35897 12251 35955 12257
rect 35986 12248 35992 12300
rect 36044 12288 36050 12300
rect 36173 12291 36231 12297
rect 36173 12288 36185 12291
rect 36044 12260 36185 12288
rect 36044 12248 36050 12260
rect 36173 12257 36185 12260
rect 36219 12288 36231 12291
rect 36998 12288 37004 12300
rect 36219 12260 37004 12288
rect 36219 12257 36231 12260
rect 36173 12251 36231 12257
rect 36998 12248 37004 12260
rect 37056 12248 37062 12300
rect 34885 12223 34943 12229
rect 34885 12220 34897 12223
rect 31444 12192 34897 12220
rect 31444 12180 31450 12192
rect 34885 12189 34897 12192
rect 34931 12189 34943 12223
rect 34885 12183 34943 12189
rect 35161 12223 35219 12229
rect 35161 12189 35173 12223
rect 35207 12189 35219 12223
rect 35161 12183 35219 12189
rect 35253 12223 35311 12229
rect 35253 12189 35265 12223
rect 35299 12220 35311 12223
rect 35342 12220 35348 12232
rect 35299 12192 35348 12220
rect 35299 12189 35311 12192
rect 35253 12183 35311 12189
rect 35342 12180 35348 12192
rect 35400 12180 35406 12232
rect 35434 12180 35440 12232
rect 35492 12220 35498 12232
rect 36081 12223 36139 12229
rect 36081 12220 36093 12223
rect 35492 12192 36093 12220
rect 35492 12180 35498 12192
rect 36081 12189 36093 12192
rect 36127 12189 36139 12223
rect 36081 12183 36139 12189
rect 36265 12223 36323 12229
rect 36265 12189 36277 12223
rect 36311 12189 36323 12223
rect 36265 12183 36323 12189
rect 30156 12124 30696 12152
rect 33781 12155 33839 12161
rect 30156 12112 30162 12124
rect 33781 12121 33793 12155
rect 33827 12152 33839 12155
rect 34698 12152 34704 12164
rect 33827 12124 34704 12152
rect 33827 12121 33839 12124
rect 33781 12115 33839 12121
rect 34698 12112 34704 12124
rect 34756 12112 34762 12164
rect 30282 12084 30288 12096
rect 28644 12056 30288 12084
rect 30282 12044 30288 12056
rect 30340 12044 30346 12096
rect 33413 12087 33471 12093
rect 33413 12053 33425 12087
rect 33459 12084 33471 12087
rect 33502 12084 33508 12096
rect 33459 12056 33508 12084
rect 33459 12053 33471 12056
rect 33413 12047 33471 12053
rect 33502 12044 33508 12056
rect 33560 12044 33566 12096
rect 33873 12087 33931 12093
rect 33873 12053 33885 12087
rect 33919 12084 33931 12087
rect 35437 12087 35495 12093
rect 35437 12084 35449 12087
rect 33919 12056 35449 12084
rect 33919 12053 33931 12056
rect 33873 12047 33931 12053
rect 35437 12053 35449 12056
rect 35483 12053 35495 12087
rect 35437 12047 35495 12053
rect 35526 12044 35532 12096
rect 35584 12084 35590 12096
rect 36280 12084 36308 12183
rect 36354 12180 36360 12232
rect 36412 12220 36418 12232
rect 36412 12192 36505 12220
rect 36412 12180 36418 12192
rect 35584 12056 36308 12084
rect 36372 12084 36400 12180
rect 37108 12152 37136 12328
rect 46492 12328 47032 12356
rect 39298 12288 39304 12300
rect 37660 12260 39304 12288
rect 37458 12220 37464 12232
rect 37419 12192 37464 12220
rect 37458 12180 37464 12192
rect 37516 12180 37522 12232
rect 37660 12229 37688 12260
rect 39298 12248 39304 12260
rect 39356 12248 39362 12300
rect 46492 12297 46520 12328
rect 47026 12316 47032 12328
rect 47084 12316 47090 12368
rect 46477 12291 46535 12297
rect 46477 12257 46489 12291
rect 46523 12257 46535 12291
rect 46658 12288 46664 12300
rect 46619 12260 46664 12288
rect 46477 12251 46535 12257
rect 46658 12248 46664 12260
rect 46716 12248 46722 12300
rect 48222 12288 48228 12300
rect 48183 12260 48228 12288
rect 48222 12248 48228 12260
rect 48280 12248 48286 12300
rect 37645 12223 37703 12229
rect 37645 12189 37657 12223
rect 37691 12189 37703 12223
rect 37645 12183 37703 12189
rect 37829 12223 37887 12229
rect 37829 12189 37841 12223
rect 37875 12189 37887 12223
rect 37829 12183 37887 12189
rect 37737 12155 37795 12161
rect 37737 12152 37749 12155
rect 37108 12124 37749 12152
rect 37737 12121 37749 12124
rect 37783 12121 37795 12155
rect 37737 12115 37795 12121
rect 37844 12084 37872 12183
rect 36372 12056 37872 12084
rect 35584 12044 35590 12056
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 19426 11840 19432 11892
rect 19484 11880 19490 11892
rect 19981 11883 20039 11889
rect 19981 11880 19993 11883
rect 19484 11852 19993 11880
rect 19484 11840 19490 11852
rect 19981 11849 19993 11852
rect 20027 11849 20039 11883
rect 19981 11843 20039 11849
rect 20346 11840 20352 11892
rect 20404 11880 20410 11892
rect 21269 11883 21327 11889
rect 21269 11880 21281 11883
rect 20404 11852 21281 11880
rect 20404 11840 20410 11852
rect 21269 11849 21281 11852
rect 21315 11880 21327 11883
rect 22278 11880 22284 11892
rect 21315 11852 22140 11880
rect 22239 11852 22284 11880
rect 21315 11849 21327 11852
rect 21269 11843 21327 11849
rect 2222 11812 2228 11824
rect 2183 11784 2228 11812
rect 2222 11772 2228 11784
rect 2280 11772 2286 11824
rect 18966 11812 18972 11824
rect 18927 11784 18972 11812
rect 18966 11772 18972 11784
rect 19024 11812 19030 11824
rect 20165 11815 20223 11821
rect 20165 11812 20177 11815
rect 19024 11784 20177 11812
rect 19024 11772 19030 11784
rect 20165 11781 20177 11784
rect 20211 11781 20223 11815
rect 20165 11775 20223 11781
rect 21192 11784 21588 11812
rect 17034 11744 17040 11756
rect 16995 11716 17040 11744
rect 17034 11704 17040 11716
rect 17092 11704 17098 11756
rect 19889 11747 19947 11753
rect 19889 11744 19901 11747
rect 19260 11716 19901 11744
rect 2038 11676 2044 11688
rect 1999 11648 2044 11676
rect 2038 11636 2044 11648
rect 2096 11636 2102 11688
rect 2774 11676 2780 11688
rect 2735 11648 2780 11676
rect 2774 11636 2780 11648
rect 2832 11636 2838 11688
rect 18230 11568 18236 11620
rect 18288 11608 18294 11620
rect 19260 11617 19288 11716
rect 19889 11713 19901 11716
rect 19935 11713 19947 11747
rect 19889 11707 19947 11713
rect 19978 11704 19984 11756
rect 20036 11744 20042 11756
rect 21192 11753 21220 11784
rect 21177 11747 21235 11753
rect 21177 11744 21189 11747
rect 20036 11716 21189 11744
rect 20036 11704 20042 11716
rect 21177 11713 21189 11716
rect 21223 11713 21235 11747
rect 21177 11707 21235 11713
rect 21453 11747 21511 11753
rect 21453 11713 21465 11747
rect 21499 11713 21511 11747
rect 21560 11744 21588 11784
rect 21910 11772 21916 11824
rect 21968 11812 21974 11824
rect 22005 11815 22063 11821
rect 22005 11812 22017 11815
rect 21968 11784 22017 11812
rect 21968 11772 21974 11784
rect 22005 11781 22017 11784
rect 22051 11781 22063 11815
rect 22112 11812 22140 11852
rect 22278 11840 22284 11852
rect 22336 11840 22342 11892
rect 22373 11883 22431 11889
rect 22373 11849 22385 11883
rect 22419 11849 22431 11883
rect 25314 11880 25320 11892
rect 25275 11852 25320 11880
rect 22373 11843 22431 11849
rect 22388 11812 22416 11843
rect 25314 11840 25320 11852
rect 25372 11840 25378 11892
rect 28721 11883 28779 11889
rect 28721 11849 28733 11883
rect 28767 11880 28779 11883
rect 28994 11880 29000 11892
rect 28767 11852 29000 11880
rect 28767 11849 28779 11852
rect 28721 11843 28779 11849
rect 28994 11840 29000 11852
rect 29052 11880 29058 11892
rect 31018 11880 31024 11892
rect 29052 11852 31024 11880
rect 29052 11840 29058 11852
rect 31018 11840 31024 11852
rect 31076 11840 31082 11892
rect 34790 11840 34796 11892
rect 34848 11880 34854 11892
rect 34885 11883 34943 11889
rect 34885 11880 34897 11883
rect 34848 11852 34897 11880
rect 34848 11840 34854 11852
rect 34885 11849 34897 11852
rect 34931 11880 34943 11883
rect 36449 11883 36507 11889
rect 34931 11852 36124 11880
rect 34931 11849 34943 11852
rect 34885 11843 34943 11849
rect 22112 11784 22416 11812
rect 35345 11815 35403 11821
rect 22005 11775 22063 11781
rect 35345 11781 35357 11815
rect 35391 11812 35403 11815
rect 35434 11812 35440 11824
rect 35391 11784 35440 11812
rect 35391 11781 35403 11784
rect 35345 11775 35403 11781
rect 35434 11772 35440 11784
rect 35492 11772 35498 11824
rect 22189 11747 22247 11753
rect 22189 11744 22201 11747
rect 21560 11716 22201 11744
rect 21453 11707 21511 11713
rect 22189 11713 22201 11716
rect 22235 11713 22247 11747
rect 22554 11744 22560 11756
rect 22515 11716 22560 11744
rect 22189 11707 22247 11713
rect 19429 11679 19487 11685
rect 19429 11645 19441 11679
rect 19475 11676 19487 11679
rect 19996 11676 20024 11704
rect 21468 11676 21496 11707
rect 22554 11704 22560 11716
rect 22612 11704 22618 11756
rect 23842 11704 23848 11756
rect 23900 11744 23906 11756
rect 28534 11744 28540 11756
rect 23900 11716 25544 11744
rect 28495 11716 28540 11744
rect 23900 11704 23906 11716
rect 21542 11676 21548 11688
rect 19475 11648 20024 11676
rect 20180 11648 21548 11676
rect 19475 11645 19487 11648
rect 19429 11639 19487 11645
rect 20180 11617 20208 11648
rect 21542 11636 21548 11648
rect 21600 11636 21606 11688
rect 25222 11636 25228 11688
rect 25280 11676 25286 11688
rect 25516 11685 25544 11716
rect 28534 11704 28540 11716
rect 28592 11704 28598 11756
rect 30650 11744 30656 11756
rect 30611 11716 30656 11744
rect 30650 11704 30656 11716
rect 30708 11704 30714 11756
rect 30837 11747 30895 11753
rect 30837 11713 30849 11747
rect 30883 11713 30895 11747
rect 30837 11707 30895 11713
rect 25409 11679 25467 11685
rect 25409 11676 25421 11679
rect 25280 11648 25421 11676
rect 25280 11636 25286 11648
rect 25409 11645 25421 11648
rect 25455 11645 25467 11679
rect 25409 11639 25467 11645
rect 25501 11679 25559 11685
rect 25501 11645 25513 11679
rect 25547 11645 25559 11679
rect 25501 11639 25559 11645
rect 29638 11636 29644 11688
rect 29696 11676 29702 11688
rect 30852 11676 30880 11707
rect 31018 11704 31024 11756
rect 31076 11744 31082 11756
rect 31113 11747 31171 11753
rect 31113 11744 31125 11747
rect 31076 11716 31125 11744
rect 31076 11704 31082 11716
rect 31113 11713 31125 11716
rect 31159 11713 31171 11747
rect 31113 11707 31171 11713
rect 31297 11747 31355 11753
rect 31297 11713 31309 11747
rect 31343 11744 31355 11747
rect 32493 11747 32551 11753
rect 32493 11744 32505 11747
rect 31343 11716 32505 11744
rect 31343 11713 31355 11716
rect 31297 11707 31355 11713
rect 32493 11713 32505 11716
rect 32539 11713 32551 11747
rect 32493 11707 32551 11713
rect 32677 11747 32735 11753
rect 32677 11713 32689 11747
rect 32723 11744 32735 11747
rect 33134 11744 33140 11756
rect 32723 11716 33140 11744
rect 32723 11713 32735 11716
rect 32677 11707 32735 11713
rect 29696 11648 30880 11676
rect 29696 11636 29702 11648
rect 19245 11611 19303 11617
rect 19245 11608 19257 11611
rect 18288 11580 19257 11608
rect 18288 11568 18294 11580
rect 19245 11577 19257 11580
rect 19291 11577 19303 11611
rect 19245 11571 19303 11577
rect 20165 11611 20223 11617
rect 20165 11577 20177 11611
rect 20211 11577 20223 11611
rect 20165 11571 20223 11577
rect 31570 11568 31576 11620
rect 31628 11608 31634 11620
rect 32692 11608 32720 11707
rect 33134 11704 33140 11716
rect 33192 11704 33198 11756
rect 33502 11744 33508 11756
rect 33463 11716 33508 11744
rect 33502 11704 33508 11716
rect 33560 11704 33566 11756
rect 34698 11744 34704 11756
rect 34659 11716 34704 11744
rect 34698 11704 34704 11716
rect 34756 11704 34762 11756
rect 35526 11744 35532 11756
rect 35487 11716 35532 11744
rect 35526 11704 35532 11716
rect 35584 11704 35590 11756
rect 35621 11747 35679 11753
rect 35621 11713 35633 11747
rect 35667 11744 35679 11747
rect 35986 11744 35992 11756
rect 35667 11716 35992 11744
rect 35667 11713 35679 11716
rect 35621 11707 35679 11713
rect 35986 11704 35992 11716
rect 36044 11704 36050 11756
rect 36096 11753 36124 11852
rect 36449 11849 36461 11883
rect 36495 11880 36507 11883
rect 36906 11880 36912 11892
rect 36495 11852 36912 11880
rect 36495 11849 36507 11852
rect 36449 11843 36507 11849
rect 36906 11840 36912 11852
rect 36964 11840 36970 11892
rect 37550 11880 37556 11892
rect 37511 11852 37556 11880
rect 37550 11840 37556 11852
rect 37608 11840 37614 11892
rect 36081 11747 36139 11753
rect 36081 11713 36093 11747
rect 36127 11713 36139 11747
rect 36262 11744 36268 11756
rect 36223 11716 36268 11744
rect 36081 11707 36139 11713
rect 36262 11704 36268 11716
rect 36320 11744 36326 11756
rect 36630 11744 36636 11756
rect 36320 11716 36636 11744
rect 36320 11704 36326 11716
rect 36630 11704 36636 11716
rect 36688 11704 36694 11756
rect 37461 11747 37519 11753
rect 37461 11713 37473 11747
rect 37507 11713 37519 11747
rect 37642 11744 37648 11756
rect 37603 11716 37648 11744
rect 37461 11707 37519 11713
rect 32769 11679 32827 11685
rect 32769 11645 32781 11679
rect 32815 11676 32827 11679
rect 33042 11676 33048 11688
rect 32815 11648 33048 11676
rect 32815 11645 32827 11648
rect 32769 11639 32827 11645
rect 33042 11636 33048 11648
rect 33100 11676 33106 11688
rect 34517 11679 34575 11685
rect 34517 11676 34529 11679
rect 33100 11648 34529 11676
rect 33100 11636 33106 11648
rect 34517 11645 34529 11648
rect 34563 11645 34575 11679
rect 37476 11676 37504 11707
rect 37642 11704 37648 11716
rect 37700 11704 37706 11756
rect 34517 11639 34575 11645
rect 36096 11648 37504 11676
rect 35342 11608 35348 11620
rect 31628 11580 32720 11608
rect 35303 11580 35348 11608
rect 31628 11568 31634 11580
rect 35342 11568 35348 11580
rect 35400 11568 35406 11620
rect 16206 11500 16212 11552
rect 16264 11540 16270 11552
rect 16853 11543 16911 11549
rect 16853 11540 16865 11543
rect 16264 11512 16865 11540
rect 16264 11500 16270 11512
rect 16853 11509 16865 11512
rect 16899 11509 16911 11543
rect 16853 11503 16911 11509
rect 21453 11543 21511 11549
rect 21453 11509 21465 11543
rect 21499 11540 21511 11543
rect 22462 11540 22468 11552
rect 21499 11512 22468 11540
rect 21499 11509 21511 11512
rect 21453 11503 21511 11509
rect 22462 11500 22468 11512
rect 22520 11500 22526 11552
rect 24946 11540 24952 11552
rect 24907 11512 24952 11540
rect 24946 11500 24952 11512
rect 25004 11500 25010 11552
rect 32306 11540 32312 11552
rect 32267 11512 32312 11540
rect 32306 11500 32312 11512
rect 32364 11500 32370 11552
rect 33321 11543 33379 11549
rect 33321 11509 33333 11543
rect 33367 11540 33379 11543
rect 33410 11540 33416 11552
rect 33367 11512 33416 11540
rect 33367 11509 33379 11512
rect 33321 11503 33379 11509
rect 33410 11500 33416 11512
rect 33468 11500 33474 11552
rect 34606 11500 34612 11552
rect 34664 11540 34670 11552
rect 36096 11549 36124 11648
rect 36081 11543 36139 11549
rect 36081 11540 36093 11543
rect 34664 11512 36093 11540
rect 34664 11500 34670 11512
rect 36081 11509 36093 11512
rect 36127 11509 36139 11543
rect 36081 11503 36139 11509
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 2038 11336 2044 11348
rect 1999 11308 2044 11336
rect 2038 11296 2044 11308
rect 2096 11296 2102 11348
rect 17310 11336 17316 11348
rect 17271 11308 17316 11336
rect 17310 11296 17316 11308
rect 17368 11296 17374 11348
rect 22922 11336 22928 11348
rect 22883 11308 22928 11336
rect 22922 11296 22928 11308
rect 22980 11296 22986 11348
rect 26510 11336 26516 11348
rect 26206 11308 26516 11336
rect 18138 11268 18144 11280
rect 18051 11240 18144 11268
rect 18138 11228 18144 11240
rect 18196 11268 18202 11280
rect 26206 11268 26234 11308
rect 26510 11296 26516 11308
rect 26568 11296 26574 11348
rect 33042 11336 33048 11348
rect 33003 11308 33048 11336
rect 33042 11296 33048 11308
rect 33100 11296 33106 11348
rect 34606 11296 34612 11348
rect 34664 11336 34670 11348
rect 35069 11339 35127 11345
rect 35069 11336 35081 11339
rect 34664 11308 35081 11336
rect 34664 11296 34670 11308
rect 35069 11305 35081 11308
rect 35115 11305 35127 11339
rect 35069 11299 35127 11305
rect 35526 11296 35532 11348
rect 35584 11336 35590 11348
rect 35621 11339 35679 11345
rect 35621 11336 35633 11339
rect 35584 11308 35633 11336
rect 35584 11296 35590 11308
rect 35621 11305 35633 11308
rect 35667 11305 35679 11339
rect 35621 11299 35679 11305
rect 18196 11240 26234 11268
rect 18196 11228 18202 11240
rect 22462 11200 22468 11212
rect 22423 11172 22468 11200
rect 22462 11160 22468 11172
rect 22520 11160 22526 11212
rect 25130 11200 25136 11212
rect 25091 11172 25136 11200
rect 25130 11160 25136 11172
rect 25188 11160 25194 11212
rect 26421 11203 26479 11209
rect 26421 11169 26433 11203
rect 26467 11200 26479 11203
rect 26602 11200 26608 11212
rect 26467 11172 26608 11200
rect 26467 11169 26479 11172
rect 26421 11163 26479 11169
rect 26602 11160 26608 11172
rect 26660 11160 26666 11212
rect 29638 11200 29644 11212
rect 28736 11172 29644 11200
rect 15933 11135 15991 11141
rect 15933 11101 15945 11135
rect 15979 11132 15991 11135
rect 17310 11132 17316 11144
rect 15979 11104 17316 11132
rect 15979 11101 15991 11104
rect 15933 11095 15991 11101
rect 16316 11076 16344 11104
rect 17310 11092 17316 11104
rect 17368 11092 17374 11144
rect 17954 11132 17960 11144
rect 17915 11104 17960 11132
rect 17954 11092 17960 11104
rect 18012 11092 18018 11144
rect 18230 11132 18236 11144
rect 18191 11104 18236 11132
rect 18230 11092 18236 11104
rect 18288 11092 18294 11144
rect 19705 11135 19763 11141
rect 19705 11101 19717 11135
rect 19751 11132 19763 11135
rect 19978 11132 19984 11144
rect 19751 11104 19984 11132
rect 19751 11101 19763 11104
rect 19705 11095 19763 11101
rect 19978 11092 19984 11104
rect 20036 11092 20042 11144
rect 22370 11092 22376 11144
rect 22428 11132 22434 11144
rect 22557 11135 22615 11141
rect 22557 11132 22569 11135
rect 22428 11104 22569 11132
rect 22428 11092 22434 11104
rect 22557 11101 22569 11104
rect 22603 11132 22615 11135
rect 23382 11132 23388 11144
rect 22603 11104 23388 11132
rect 22603 11101 22615 11104
rect 22557 11095 22615 11101
rect 23382 11092 23388 11104
rect 23440 11092 23446 11144
rect 24946 11132 24952 11144
rect 24907 11104 24952 11132
rect 24946 11092 24952 11104
rect 25004 11092 25010 11144
rect 26694 11132 26700 11144
rect 26655 11104 26700 11132
rect 26694 11092 26700 11104
rect 26752 11092 26758 11144
rect 28537 11135 28595 11141
rect 28537 11132 28549 11135
rect 26804 11104 28549 11132
rect 16206 11073 16212 11076
rect 16200 11064 16212 11073
rect 16167 11036 16212 11064
rect 16200 11027 16212 11036
rect 16206 11024 16212 11027
rect 16264 11024 16270 11076
rect 16298 11024 16304 11076
rect 16356 11024 16362 11076
rect 18248 11064 18276 11092
rect 23658 11064 23664 11076
rect 18248 11036 23664 11064
rect 23658 11024 23664 11036
rect 23716 11064 23722 11076
rect 26804 11064 26832 11104
rect 28537 11101 28549 11104
rect 28583 11132 28595 11135
rect 28626 11132 28632 11144
rect 28583 11104 28632 11132
rect 28583 11101 28595 11104
rect 28537 11095 28595 11101
rect 28626 11092 28632 11104
rect 28684 11092 28690 11144
rect 28736 11141 28764 11172
rect 29638 11160 29644 11172
rect 29696 11160 29702 11212
rect 28721 11135 28779 11141
rect 28721 11101 28733 11135
rect 28767 11101 28779 11135
rect 28994 11132 29000 11144
rect 28955 11104 29000 11132
rect 28721 11095 28779 11101
rect 28994 11092 29000 11104
rect 29052 11092 29058 11144
rect 29086 11092 29092 11144
rect 29144 11132 29150 11144
rect 29733 11135 29791 11141
rect 29733 11132 29745 11135
rect 29144 11104 29745 11132
rect 29144 11092 29150 11104
rect 29733 11101 29745 11104
rect 29779 11132 29791 11135
rect 29822 11132 29828 11144
rect 29779 11104 29828 11132
rect 29779 11101 29791 11104
rect 29733 11095 29791 11101
rect 29822 11092 29828 11104
rect 29880 11132 29886 11144
rect 31662 11132 31668 11144
rect 29880 11104 31668 11132
rect 29880 11092 29886 11104
rect 31662 11092 31668 11104
rect 31720 11092 31726 11144
rect 31932 11135 31990 11141
rect 31932 11101 31944 11135
rect 31978 11132 31990 11135
rect 32306 11132 32312 11144
rect 31978 11104 32312 11132
rect 31978 11101 31990 11104
rect 31932 11095 31990 11101
rect 32306 11092 32312 11104
rect 32364 11092 32370 11144
rect 33060 11132 33088 11296
rect 35636 11268 35664 11299
rect 36262 11296 36268 11348
rect 36320 11336 36326 11348
rect 37093 11339 37151 11345
rect 37093 11336 37105 11339
rect 36320 11308 37105 11336
rect 36320 11296 36326 11308
rect 37093 11305 37105 11308
rect 37139 11305 37151 11339
rect 37093 11299 37151 11305
rect 37642 11268 37648 11280
rect 35636 11240 37648 11268
rect 34698 11160 34704 11212
rect 34756 11200 34762 11212
rect 34756 11172 35112 11200
rect 34756 11160 34762 11172
rect 35084 11141 35112 11172
rect 35728 11172 36492 11200
rect 35728 11141 35756 11172
rect 34885 11135 34943 11141
rect 34885 11132 34897 11135
rect 33060 11104 34897 11132
rect 34885 11101 34897 11104
rect 34931 11101 34943 11135
rect 34885 11095 34943 11101
rect 35069 11135 35127 11141
rect 35069 11101 35081 11135
rect 35115 11101 35127 11135
rect 35069 11095 35127 11101
rect 35529 11135 35587 11141
rect 35529 11101 35541 11135
rect 35575 11101 35587 11135
rect 35529 11095 35587 11101
rect 35713 11135 35771 11141
rect 35713 11101 35725 11135
rect 35759 11101 35771 11135
rect 36357 11135 36415 11141
rect 36357 11132 36369 11135
rect 35713 11095 35771 11101
rect 35820 11104 36369 11132
rect 23716 11036 26832 11064
rect 26881 11067 26939 11073
rect 23716 11024 23722 11036
rect 26881 11033 26893 11067
rect 26927 11064 26939 11067
rect 28258 11064 28264 11076
rect 26927 11036 28264 11064
rect 26927 11033 26939 11036
rect 26881 11027 26939 11033
rect 28258 11024 28264 11036
rect 28316 11024 28322 11076
rect 29546 11024 29552 11076
rect 29604 11064 29610 11076
rect 29978 11067 30036 11073
rect 29978 11064 29990 11067
rect 29604 11036 29990 11064
rect 29604 11024 29610 11036
rect 29978 11033 29990 11036
rect 30024 11033 30036 11067
rect 35544 11064 35572 11095
rect 35820 11064 35848 11104
rect 36357 11101 36369 11104
rect 36403 11101 36415 11135
rect 36357 11095 36415 11101
rect 29978 11027 30036 11033
rect 31128 11036 35848 11064
rect 36173 11067 36231 11073
rect 31128 11008 31156 11036
rect 36173 11033 36185 11067
rect 36219 11064 36231 11067
rect 36464 11064 36492 11172
rect 37200 11141 37228 11240
rect 37642 11228 37648 11240
rect 37700 11228 37706 11280
rect 36541 11135 36599 11141
rect 36541 11101 36553 11135
rect 36587 11132 36599 11135
rect 37001 11135 37059 11141
rect 37001 11132 37013 11135
rect 36587 11104 37013 11132
rect 36587 11101 36599 11104
rect 36541 11095 36599 11101
rect 37001 11101 37013 11104
rect 37047 11101 37059 11135
rect 37001 11095 37059 11101
rect 37185 11135 37243 11141
rect 37185 11101 37197 11135
rect 37231 11101 37243 11135
rect 37185 11095 37243 11101
rect 37458 11064 37464 11076
rect 36219 11036 37464 11064
rect 36219 11033 36231 11036
rect 36173 11027 36231 11033
rect 37458 11024 37464 11036
rect 37516 11024 37522 11076
rect 17770 10996 17776 11008
rect 17731 10968 17776 10996
rect 17770 10956 17776 10968
rect 17828 10956 17834 11008
rect 19426 10956 19432 11008
rect 19484 10996 19490 11008
rect 19521 10999 19579 11005
rect 19521 10996 19533 10999
rect 19484 10968 19533 10996
rect 19484 10956 19490 10968
rect 19521 10965 19533 10968
rect 19567 10965 19579 10999
rect 19521 10959 19579 10965
rect 24581 10999 24639 11005
rect 24581 10965 24593 10999
rect 24627 10996 24639 10999
rect 24670 10996 24676 11008
rect 24627 10968 24676 10996
rect 24627 10965 24639 10968
rect 24581 10959 24639 10965
rect 24670 10956 24676 10968
rect 24728 10956 24734 11008
rect 25038 10996 25044 11008
rect 24999 10968 25044 10996
rect 25038 10956 25044 10968
rect 25096 10956 25102 11008
rect 29181 10999 29239 11005
rect 29181 10965 29193 10999
rect 29227 10996 29239 10999
rect 29730 10996 29736 11008
rect 29227 10968 29736 10996
rect 29227 10965 29239 10968
rect 29181 10959 29239 10965
rect 29730 10956 29736 10968
rect 29788 10956 29794 11008
rect 31110 10996 31116 11008
rect 31071 10968 31116 10996
rect 31110 10956 31116 10968
rect 31168 10956 31174 11008
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 19334 10792 19340 10804
rect 19168 10764 19340 10792
rect 17580 10727 17638 10733
rect 17580 10693 17592 10727
rect 17626 10724 17638 10727
rect 17770 10724 17776 10736
rect 17626 10696 17776 10724
rect 17626 10693 17638 10696
rect 17580 10687 17638 10693
rect 17770 10684 17776 10696
rect 17828 10684 17834 10736
rect 2961 10659 3019 10665
rect 2961 10625 2973 10659
rect 3007 10656 3019 10659
rect 4614 10656 4620 10668
rect 3007 10628 4620 10656
rect 3007 10625 3019 10628
rect 2961 10619 3019 10625
rect 4614 10616 4620 10628
rect 4672 10616 4678 10668
rect 17310 10656 17316 10668
rect 17271 10628 17316 10656
rect 17310 10616 17316 10628
rect 17368 10616 17374 10668
rect 19168 10665 19196 10764
rect 19334 10752 19340 10764
rect 19392 10752 19398 10804
rect 22554 10752 22560 10804
rect 22612 10792 22618 10804
rect 22649 10795 22707 10801
rect 22649 10792 22661 10795
rect 22612 10764 22661 10792
rect 22612 10752 22618 10764
rect 22649 10761 22661 10764
rect 22695 10761 22707 10795
rect 22649 10755 22707 10761
rect 24581 10795 24639 10801
rect 24581 10761 24593 10795
rect 24627 10792 24639 10795
rect 25038 10792 25044 10804
rect 24627 10764 25044 10792
rect 24627 10761 24639 10764
rect 24581 10755 24639 10761
rect 19426 10733 19432 10736
rect 19420 10724 19432 10733
rect 19387 10696 19432 10724
rect 19420 10687 19432 10696
rect 19426 10684 19432 10687
rect 19484 10684 19490 10736
rect 21542 10684 21548 10736
rect 21600 10724 21606 10736
rect 22278 10724 22284 10736
rect 21600 10696 22140 10724
rect 22191 10696 22284 10724
rect 21600 10684 21606 10696
rect 19153 10659 19211 10665
rect 19153 10625 19165 10659
rect 19199 10625 19211 10659
rect 19153 10619 19211 10625
rect 20714 10616 20720 10668
rect 20772 10656 20778 10668
rect 21269 10659 21327 10665
rect 21269 10656 21281 10659
rect 20772 10628 21281 10656
rect 20772 10616 20778 10628
rect 21269 10625 21281 10628
rect 21315 10625 21327 10659
rect 21450 10656 21456 10668
rect 21411 10628 21456 10656
rect 21269 10619 21327 10625
rect 21450 10616 21456 10628
rect 21508 10616 21514 10668
rect 21818 10616 21824 10668
rect 21876 10656 21882 10668
rect 22112 10665 22140 10696
rect 22278 10684 22284 10696
rect 22336 10724 22342 10736
rect 23937 10727 23995 10733
rect 23937 10724 23949 10727
rect 22336 10696 23949 10724
rect 22336 10684 22342 10696
rect 23937 10693 23949 10696
rect 23983 10693 23995 10727
rect 23937 10687 23995 10693
rect 22005 10659 22063 10665
rect 22005 10656 22017 10659
rect 21876 10628 22017 10656
rect 21876 10616 21882 10628
rect 22005 10625 22017 10628
rect 22051 10625 22063 10659
rect 22005 10619 22063 10625
rect 22098 10659 22156 10665
rect 22098 10625 22110 10659
rect 22144 10625 22156 10659
rect 22098 10619 22156 10625
rect 22186 10616 22192 10668
rect 22244 10656 22250 10668
rect 22373 10659 22431 10665
rect 22373 10656 22385 10659
rect 22244 10628 22385 10656
rect 22244 10616 22250 10628
rect 22373 10625 22385 10628
rect 22419 10625 22431 10659
rect 22373 10619 22431 10625
rect 22511 10659 22569 10665
rect 22511 10625 22523 10659
rect 22557 10656 22569 10659
rect 22738 10656 22744 10668
rect 22557 10628 22744 10656
rect 22557 10625 22569 10628
rect 22511 10619 22569 10625
rect 22738 10616 22744 10628
rect 22796 10656 22802 10668
rect 22796 10628 23336 10656
rect 22796 10616 22802 10628
rect 23109 10591 23167 10597
rect 23109 10588 23121 10591
rect 22204 10560 23121 10588
rect 22204 10464 22232 10560
rect 23109 10557 23121 10560
rect 23155 10557 23167 10591
rect 23308 10588 23336 10628
rect 23382 10616 23388 10668
rect 23440 10656 23446 10668
rect 23845 10659 23903 10665
rect 23845 10656 23857 10659
rect 23440 10628 23857 10656
rect 23440 10616 23446 10628
rect 23845 10625 23857 10628
rect 23891 10625 23903 10659
rect 24026 10656 24032 10668
rect 23987 10628 24032 10656
rect 23845 10619 23903 10625
rect 24026 10616 24032 10628
rect 24084 10616 24090 10668
rect 24596 10588 24624 10755
rect 25038 10752 25044 10764
rect 25096 10752 25102 10804
rect 29546 10792 29552 10804
rect 29507 10764 29552 10792
rect 29546 10752 29552 10764
rect 29604 10752 29610 10804
rect 34517 10795 34575 10801
rect 34517 10761 34529 10795
rect 34563 10792 34575 10795
rect 34698 10792 34704 10804
rect 34563 10764 34704 10792
rect 34563 10761 34575 10764
rect 34517 10755 34575 10761
rect 34698 10752 34704 10764
rect 34756 10752 34762 10804
rect 26206 10696 28580 10724
rect 24854 10616 24860 10668
rect 24912 10656 24918 10668
rect 25694 10659 25752 10665
rect 25694 10656 25706 10659
rect 24912 10628 25706 10656
rect 24912 10616 24918 10628
rect 25694 10625 25706 10628
rect 25740 10625 25752 10659
rect 25694 10619 25752 10625
rect 25961 10659 26019 10665
rect 25961 10625 25973 10659
rect 26007 10656 26019 10659
rect 26206 10656 26234 10696
rect 26007 10628 26234 10656
rect 26007 10625 26019 10628
rect 25961 10619 26019 10625
rect 28258 10616 28264 10668
rect 28316 10665 28322 10668
rect 28552 10665 28580 10696
rect 28316 10656 28328 10665
rect 28537 10659 28595 10665
rect 28316 10628 28361 10656
rect 28316 10619 28328 10628
rect 28537 10625 28549 10659
rect 28583 10656 28595 10659
rect 29086 10656 29092 10668
rect 28583 10628 29092 10656
rect 28583 10625 28595 10628
rect 28537 10619 28595 10625
rect 28316 10616 28322 10619
rect 29086 10616 29092 10628
rect 29144 10616 29150 10668
rect 29730 10656 29736 10668
rect 29691 10628 29736 10656
rect 29730 10616 29736 10628
rect 29788 10616 29794 10668
rect 30009 10659 30067 10665
rect 30009 10625 30021 10659
rect 30055 10656 30067 10659
rect 31110 10656 31116 10668
rect 30055 10628 31116 10656
rect 30055 10625 30067 10628
rect 30009 10619 30067 10625
rect 31110 10616 31116 10628
rect 31168 10616 31174 10668
rect 31662 10616 31668 10668
rect 31720 10656 31726 10668
rect 33410 10665 33416 10668
rect 33137 10659 33195 10665
rect 33137 10656 33149 10659
rect 31720 10628 33149 10656
rect 31720 10616 31726 10628
rect 33137 10625 33149 10628
rect 33183 10625 33195 10659
rect 33404 10656 33416 10665
rect 33371 10628 33416 10656
rect 33137 10619 33195 10625
rect 33404 10619 33416 10628
rect 33410 10616 33416 10619
rect 33468 10616 33474 10668
rect 23308 10560 24624 10588
rect 29917 10591 29975 10597
rect 23109 10551 23167 10557
rect 29917 10557 29929 10591
rect 29963 10588 29975 10591
rect 31570 10588 31576 10600
rect 29963 10560 31576 10588
rect 29963 10557 29975 10560
rect 29917 10551 29975 10557
rect 31570 10548 31576 10560
rect 31628 10548 31634 10600
rect 22462 10480 22468 10532
rect 22520 10520 22526 10532
rect 23293 10523 23351 10529
rect 23293 10520 23305 10523
rect 22520 10492 23305 10520
rect 22520 10480 22526 10492
rect 23293 10489 23305 10492
rect 23339 10489 23351 10523
rect 23293 10483 23351 10489
rect 2314 10452 2320 10464
rect 2275 10424 2320 10452
rect 2314 10412 2320 10424
rect 2372 10412 2378 10464
rect 2869 10455 2927 10461
rect 2869 10421 2881 10455
rect 2915 10452 2927 10455
rect 3234 10452 3240 10464
rect 2915 10424 3240 10452
rect 2915 10421 2927 10424
rect 2869 10415 2927 10421
rect 3234 10412 3240 10424
rect 3292 10412 3298 10464
rect 18693 10455 18751 10461
rect 18693 10421 18705 10455
rect 18739 10452 18751 10455
rect 18874 10452 18880 10464
rect 18739 10424 18880 10452
rect 18739 10421 18751 10424
rect 18693 10415 18751 10421
rect 18874 10412 18880 10424
rect 18932 10412 18938 10464
rect 20533 10455 20591 10461
rect 20533 10421 20545 10455
rect 20579 10452 20591 10455
rect 20714 10452 20720 10464
rect 20579 10424 20720 10452
rect 20579 10421 20591 10424
rect 20533 10415 20591 10421
rect 20714 10412 20720 10424
rect 20772 10412 20778 10464
rect 21361 10455 21419 10461
rect 21361 10421 21373 10455
rect 21407 10452 21419 10455
rect 22186 10452 22192 10464
rect 21407 10424 22192 10452
rect 21407 10421 21419 10424
rect 21361 10415 21419 10421
rect 22186 10412 22192 10424
rect 22244 10412 22250 10464
rect 23198 10452 23204 10464
rect 23159 10424 23204 10452
rect 23198 10412 23204 10424
rect 23256 10412 23262 10464
rect 23842 10412 23848 10464
rect 23900 10452 23906 10464
rect 25222 10452 25228 10464
rect 23900 10424 25228 10452
rect 23900 10412 23906 10424
rect 25222 10412 25228 10424
rect 25280 10412 25286 10464
rect 26878 10412 26884 10464
rect 26936 10452 26942 10464
rect 27157 10455 27215 10461
rect 27157 10452 27169 10455
rect 26936 10424 27169 10452
rect 26936 10412 26942 10424
rect 27157 10421 27169 10424
rect 27203 10421 27215 10455
rect 27157 10415 27215 10421
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 17954 10208 17960 10260
rect 18012 10248 18018 10260
rect 18233 10251 18291 10257
rect 18233 10248 18245 10251
rect 18012 10220 18245 10248
rect 18012 10208 18018 10220
rect 18233 10217 18245 10220
rect 18279 10217 18291 10251
rect 18233 10211 18291 10217
rect 19889 10251 19947 10257
rect 19889 10217 19901 10251
rect 19935 10248 19947 10251
rect 19978 10248 19984 10260
rect 19935 10220 19984 10248
rect 19935 10217 19947 10220
rect 19889 10211 19947 10217
rect 19978 10208 19984 10220
rect 20036 10208 20042 10260
rect 20714 10208 20720 10260
rect 20772 10248 20778 10260
rect 21637 10251 21695 10257
rect 21637 10248 21649 10251
rect 20772 10220 21649 10248
rect 20772 10208 20778 10220
rect 21637 10217 21649 10220
rect 21683 10217 21695 10251
rect 21818 10248 21824 10260
rect 21779 10220 21824 10248
rect 21637 10211 21695 10217
rect 21818 10208 21824 10220
rect 21876 10208 21882 10260
rect 26237 10251 26295 10257
rect 21928 10220 25544 10248
rect 2314 10140 2320 10192
rect 2372 10180 2378 10192
rect 21928 10180 21956 10220
rect 23842 10180 23848 10192
rect 2372 10152 3464 10180
rect 2372 10140 2378 10152
rect 1578 10112 1584 10124
rect 1539 10084 1584 10112
rect 1578 10072 1584 10084
rect 1636 10072 1642 10124
rect 3234 10112 3240 10124
rect 3195 10084 3240 10112
rect 3234 10072 3240 10084
rect 3292 10072 3298 10124
rect 3436 10121 3464 10152
rect 18708 10152 21956 10180
rect 22066 10152 23520 10180
rect 23803 10152 23848 10180
rect 3421 10115 3479 10121
rect 3421 10081 3433 10115
rect 3467 10081 3479 10115
rect 3421 10075 3479 10081
rect 18414 10044 18420 10056
rect 18375 10016 18420 10044
rect 18414 10004 18420 10016
rect 18472 10004 18478 10056
rect 18506 10004 18512 10056
rect 18564 10044 18570 10056
rect 18708 10053 18736 10152
rect 20530 10112 20536 10124
rect 20443 10084 20536 10112
rect 20530 10072 20536 10084
rect 20588 10112 20594 10124
rect 22066 10112 22094 10152
rect 20588 10084 22094 10112
rect 20588 10072 20594 10084
rect 23198 10072 23204 10124
rect 23256 10112 23262 10124
rect 23385 10115 23443 10121
rect 23385 10112 23397 10115
rect 23256 10084 23397 10112
rect 23256 10072 23262 10084
rect 23385 10081 23397 10084
rect 23431 10081 23443 10115
rect 23492 10112 23520 10152
rect 23842 10140 23848 10152
rect 23900 10140 23906 10192
rect 24854 10180 24860 10192
rect 24815 10152 24860 10180
rect 24854 10140 24860 10152
rect 24912 10140 24918 10192
rect 25130 10112 25136 10124
rect 23492 10084 25136 10112
rect 23385 10075 23443 10081
rect 25130 10072 25136 10084
rect 25188 10072 25194 10124
rect 25516 10112 25544 10220
rect 26237 10217 26249 10251
rect 26283 10248 26295 10251
rect 26694 10248 26700 10260
rect 26283 10220 26700 10248
rect 26283 10217 26295 10220
rect 26237 10211 26295 10217
rect 26694 10208 26700 10220
rect 26752 10208 26758 10260
rect 26234 10112 26240 10124
rect 25516 10084 26240 10112
rect 26234 10072 26240 10084
rect 26292 10112 26298 10124
rect 26292 10084 26740 10112
rect 26292 10072 26298 10084
rect 18693 10047 18751 10053
rect 18693 10044 18705 10047
rect 18564 10016 18705 10044
rect 18564 10004 18570 10016
rect 18693 10013 18705 10016
rect 18739 10013 18751 10047
rect 18874 10044 18880 10056
rect 18835 10016 18880 10044
rect 18693 10007 18751 10013
rect 18874 10004 18880 10016
rect 18932 10004 18938 10056
rect 20349 10047 20407 10053
rect 20349 10013 20361 10047
rect 20395 10044 20407 10047
rect 20714 10044 20720 10056
rect 20395 10016 20720 10044
rect 20395 10013 20407 10016
rect 20349 10007 20407 10013
rect 20714 10004 20720 10016
rect 20772 10004 20778 10056
rect 22738 10004 22744 10056
rect 22796 10044 22802 10056
rect 22833 10047 22891 10053
rect 22833 10044 22845 10047
rect 22796 10016 22845 10044
rect 22796 10004 22802 10016
rect 22833 10013 22845 10016
rect 22879 10013 22891 10047
rect 22833 10007 22891 10013
rect 23477 10047 23535 10053
rect 23477 10013 23489 10047
rect 23523 10044 23535 10047
rect 24026 10044 24032 10056
rect 23523 10016 24032 10044
rect 23523 10013 23535 10016
rect 23477 10007 23535 10013
rect 24026 10004 24032 10016
rect 24084 10004 24090 10056
rect 24670 10044 24676 10056
rect 24631 10016 24676 10044
rect 24670 10004 24676 10016
rect 24728 10004 24734 10056
rect 25314 10004 25320 10056
rect 25372 10044 25378 10056
rect 25590 10044 25596 10056
rect 25372 10016 25596 10044
rect 25372 10004 25378 10016
rect 25590 10004 25596 10016
rect 25648 10044 25654 10056
rect 26712 10053 26740 10084
rect 26421 10047 26479 10053
rect 26421 10044 26433 10047
rect 25648 10016 26433 10044
rect 25648 10004 25654 10016
rect 26421 10013 26433 10016
rect 26467 10013 26479 10047
rect 26421 10007 26479 10013
rect 26697 10047 26755 10053
rect 26697 10013 26709 10047
rect 26743 10013 26755 10047
rect 26878 10044 26884 10056
rect 26839 10016 26884 10044
rect 26697 10007 26755 10013
rect 26878 10004 26884 10016
rect 26936 10004 26942 10056
rect 18892 9908 18920 10004
rect 20257 9979 20315 9985
rect 20257 9945 20269 9979
rect 20303 9976 20315 9979
rect 20806 9976 20812 9988
rect 20303 9948 20812 9976
rect 20303 9945 20315 9948
rect 20257 9939 20315 9945
rect 20806 9936 20812 9948
rect 20864 9936 20870 9988
rect 21450 9976 21456 9988
rect 21363 9948 21456 9976
rect 21450 9936 21456 9948
rect 21508 9936 21514 9988
rect 22278 9936 22284 9988
rect 22336 9976 22342 9988
rect 22649 9979 22707 9985
rect 22649 9976 22661 9979
rect 22336 9948 22661 9976
rect 22336 9936 22342 9948
rect 22649 9945 22661 9948
rect 22695 9976 22707 9979
rect 23198 9976 23204 9988
rect 22695 9948 23204 9976
rect 22695 9945 22707 9948
rect 22649 9939 22707 9945
rect 23198 9936 23204 9948
rect 23256 9976 23262 9988
rect 23256 9948 24716 9976
rect 23256 9936 23262 9948
rect 21266 9908 21272 9920
rect 18892 9880 21272 9908
rect 21266 9868 21272 9880
rect 21324 9908 21330 9920
rect 21468 9908 21496 9936
rect 21324 9880 21496 9908
rect 21663 9911 21721 9917
rect 21324 9868 21330 9880
rect 21663 9877 21675 9911
rect 21709 9908 21721 9911
rect 22465 9911 22523 9917
rect 22465 9908 22477 9911
rect 21709 9880 22477 9908
rect 21709 9877 21721 9880
rect 21663 9871 21721 9877
rect 22465 9877 22477 9880
rect 22511 9908 22523 9911
rect 23290 9908 23296 9920
rect 22511 9880 23296 9908
rect 22511 9877 22523 9880
rect 22465 9871 22523 9877
rect 23290 9868 23296 9880
rect 23348 9868 23354 9920
rect 24688 9908 24716 9948
rect 26896 9908 26924 10004
rect 24688 9880 26924 9908
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 18414 9664 18420 9716
rect 18472 9704 18478 9716
rect 22189 9707 22247 9713
rect 18472 9676 22140 9704
rect 18472 9664 18478 9676
rect 20714 9596 20720 9648
rect 20772 9636 20778 9648
rect 21085 9639 21143 9645
rect 21085 9636 21097 9639
rect 20772 9608 21097 9636
rect 20772 9596 20778 9608
rect 21085 9605 21097 9608
rect 21131 9605 21143 9639
rect 21266 9636 21272 9648
rect 21227 9608 21272 9636
rect 21085 9599 21143 9605
rect 21266 9596 21272 9608
rect 21324 9596 21330 9648
rect 22112 9636 22140 9676
rect 22189 9673 22201 9707
rect 22235 9704 22247 9707
rect 22370 9704 22376 9716
rect 22235 9676 22376 9704
rect 22235 9673 22247 9676
rect 22189 9667 22247 9673
rect 22370 9664 22376 9676
rect 22428 9664 22434 9716
rect 23845 9707 23903 9713
rect 22480 9676 23796 9704
rect 22480 9636 22508 9676
rect 22112 9608 22508 9636
rect 23768 9636 23796 9676
rect 23845 9673 23857 9707
rect 23891 9704 23903 9707
rect 24026 9704 24032 9716
rect 23891 9676 24032 9704
rect 23891 9673 23903 9676
rect 23845 9667 23903 9673
rect 24026 9664 24032 9676
rect 24084 9664 24090 9716
rect 25314 9704 25320 9716
rect 24136 9676 25320 9704
rect 24136 9636 24164 9676
rect 25314 9664 25320 9676
rect 25372 9664 25378 9716
rect 23768 9608 24164 9636
rect 21453 9571 21511 9577
rect 21453 9537 21465 9571
rect 21499 9568 21511 9571
rect 22005 9571 22063 9577
rect 22005 9568 22017 9571
rect 21499 9540 22017 9568
rect 21499 9537 21511 9540
rect 21453 9531 21511 9537
rect 22005 9537 22017 9540
rect 22051 9537 22063 9571
rect 22186 9568 22192 9580
rect 22147 9540 22192 9568
rect 22005 9531 22063 9537
rect 22186 9528 22192 9540
rect 22244 9528 22250 9580
rect 22738 9528 22744 9580
rect 22796 9568 22802 9580
rect 23017 9571 23075 9577
rect 23017 9568 23029 9571
rect 22796 9540 23029 9568
rect 22796 9528 22802 9540
rect 23017 9537 23029 9540
rect 23063 9537 23075 9571
rect 23198 9568 23204 9580
rect 23159 9540 23204 9568
rect 23017 9531 23075 9537
rect 23198 9528 23204 9540
rect 23256 9528 23262 9580
rect 23290 9528 23296 9580
rect 23348 9568 23354 9580
rect 23661 9571 23719 9577
rect 23661 9568 23673 9571
rect 23348 9540 23673 9568
rect 23348 9528 23354 9540
rect 23661 9537 23673 9540
rect 23707 9537 23719 9571
rect 23661 9531 23719 9537
rect 23845 9571 23903 9577
rect 23845 9537 23857 9571
rect 23891 9537 23903 9571
rect 23845 9531 23903 9537
rect 2038 9500 2044 9512
rect 1999 9472 2044 9500
rect 2038 9460 2044 9472
rect 2096 9460 2102 9512
rect 2225 9503 2283 9509
rect 2225 9469 2237 9503
rect 2271 9500 2283 9503
rect 2866 9500 2872 9512
rect 2271 9472 2872 9500
rect 2271 9469 2283 9472
rect 2225 9463 2283 9469
rect 2866 9460 2872 9472
rect 2924 9460 2930 9512
rect 2958 9460 2964 9512
rect 3016 9500 3022 9512
rect 23109 9503 23167 9509
rect 3016 9472 3061 9500
rect 3016 9460 3022 9472
rect 23109 9469 23121 9503
rect 23155 9500 23167 9503
rect 23860 9500 23888 9531
rect 23155 9472 23888 9500
rect 23155 9469 23167 9472
rect 23109 9463 23167 9469
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 2038 9120 2044 9172
rect 2096 9160 2102 9172
rect 2133 9163 2191 9169
rect 2133 9160 2145 9163
rect 2096 9132 2145 9160
rect 2096 9120 2102 9132
rect 2133 9129 2145 9132
rect 2179 9129 2191 9163
rect 2866 9160 2872 9172
rect 2827 9132 2872 9160
rect 2133 9123 2191 9129
rect 2866 9120 2872 9132
rect 2924 9120 2930 9172
rect 39574 9120 39580 9172
rect 39632 9160 39638 9172
rect 47949 9163 48007 9169
rect 47949 9160 47961 9163
rect 39632 9132 47961 9160
rect 39632 9120 39638 9132
rect 47949 9129 47961 9132
rect 47995 9129 48007 9163
rect 47949 9123 48007 9129
rect 2774 8916 2780 8968
rect 2832 8956 2838 8968
rect 2961 8959 3019 8965
rect 2961 8956 2973 8959
rect 2832 8928 2973 8956
rect 2832 8916 2838 8928
rect 2961 8925 2973 8928
rect 3007 8956 3019 8959
rect 4982 8956 4988 8968
rect 3007 8928 4988 8956
rect 3007 8925 3019 8928
rect 2961 8919 3019 8925
rect 4982 8916 4988 8928
rect 5040 8916 5046 8968
rect 48222 8888 48228 8900
rect 48183 8860 48228 8888
rect 48222 8848 48228 8860
rect 48280 8848 48286 8900
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 48222 8440 48228 8492
rect 48280 8480 48286 8492
rect 48317 8483 48375 8489
rect 48317 8480 48329 8483
rect 48280 8452 48329 8480
rect 48280 8440 48286 8452
rect 48317 8449 48329 8452
rect 48363 8449 48375 8483
rect 48317 8443 48375 8449
rect 28534 8372 28540 8424
rect 28592 8412 28598 8424
rect 48041 8415 48099 8421
rect 48041 8412 48053 8415
rect 28592 8384 48053 8412
rect 28592 8372 28598 8384
rect 48041 8381 48053 8384
rect 48087 8381 48099 8415
rect 48041 8375 48099 8381
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 3418 7828 3424 7880
rect 3476 7868 3482 7880
rect 3476 7840 3521 7868
rect 3476 7828 3482 7840
rect 1578 7800 1584 7812
rect 1539 7772 1584 7800
rect 1578 7760 1584 7772
rect 1636 7760 1642 7812
rect 2866 7760 2872 7812
rect 2924 7800 2930 7812
rect 3237 7803 3295 7809
rect 3237 7800 3249 7803
rect 2924 7772 3249 7800
rect 2924 7760 2930 7772
rect 3237 7769 3249 7772
rect 3283 7769 3295 7803
rect 3237 7763 3295 7769
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 2866 7528 2872 7540
rect 2827 7500 2872 7528
rect 2866 7488 2872 7500
rect 2924 7488 2930 7540
rect 3418 7460 3424 7472
rect 2332 7432 3424 7460
rect 2332 7401 2360 7432
rect 3418 7420 3424 7432
rect 3476 7420 3482 7472
rect 2317 7395 2375 7401
rect 2317 7361 2329 7395
rect 2363 7361 2375 7395
rect 2317 7355 2375 7361
rect 2777 7395 2835 7401
rect 2777 7361 2789 7395
rect 2823 7392 2835 7395
rect 3142 7392 3148 7404
rect 2823 7364 3148 7392
rect 2823 7361 2835 7364
rect 2777 7355 2835 7361
rect 3142 7352 3148 7364
rect 3200 7392 3206 7404
rect 5442 7392 5448 7404
rect 3200 7364 5448 7392
rect 3200 7352 3206 7364
rect 5442 7352 5448 7364
rect 5500 7352 5506 7404
rect 3418 7188 3424 7200
rect 3379 7160 3424 7188
rect 3418 7148 3424 7160
rect 3476 7148 3482 7200
rect 43254 7188 43260 7200
rect 43215 7160 43260 7188
rect 43254 7148 43260 7160
rect 43312 7148 43318 7200
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 1578 6848 1584 6860
rect 1539 6820 1584 6848
rect 1578 6808 1584 6820
rect 1636 6808 1642 6860
rect 3418 6848 3424 6860
rect 3379 6820 3424 6848
rect 3418 6808 3424 6820
rect 3476 6808 3482 6860
rect 32214 6808 32220 6860
rect 32272 6848 32278 6860
rect 32309 6851 32367 6857
rect 32309 6848 32321 6851
rect 32272 6820 32321 6848
rect 32272 6808 32278 6820
rect 32309 6817 32321 6820
rect 32355 6817 32367 6851
rect 32309 6811 32367 6817
rect 42797 6851 42855 6857
rect 42797 6817 42809 6851
rect 42843 6848 42855 6851
rect 43254 6848 43260 6860
rect 42843 6820 43260 6848
rect 42843 6817 42855 6820
rect 42797 6811 42855 6817
rect 43254 6808 43260 6820
rect 43312 6808 43318 6860
rect 44637 6851 44695 6857
rect 44637 6817 44649 6851
rect 44683 6848 44695 6851
rect 46842 6848 46848 6860
rect 44683 6820 46848 6848
rect 44683 6817 44695 6820
rect 44637 6811 44695 6817
rect 46842 6808 46848 6820
rect 46900 6808 46906 6860
rect 31389 6783 31447 6789
rect 31389 6749 31401 6783
rect 31435 6780 31447 6783
rect 31849 6783 31907 6789
rect 31849 6780 31861 6783
rect 31435 6752 31861 6780
rect 31435 6749 31447 6752
rect 31389 6743 31447 6749
rect 31849 6749 31861 6752
rect 31895 6749 31907 6783
rect 31849 6743 31907 6749
rect 46106 6740 46112 6792
rect 46164 6780 46170 6792
rect 46201 6783 46259 6789
rect 46201 6780 46213 6783
rect 46164 6752 46213 6780
rect 46164 6740 46170 6752
rect 46201 6749 46213 6752
rect 46247 6749 46259 6783
rect 46201 6743 46259 6749
rect 47029 6783 47087 6789
rect 47029 6749 47041 6783
rect 47075 6780 47087 6783
rect 47302 6780 47308 6792
rect 47075 6752 47308 6780
rect 47075 6749 47087 6752
rect 47029 6743 47087 6749
rect 47302 6740 47308 6752
rect 47360 6740 47366 6792
rect 47670 6780 47676 6792
rect 47631 6752 47676 6780
rect 47670 6740 47676 6752
rect 47728 6740 47734 6792
rect 47946 6740 47952 6792
rect 48004 6780 48010 6792
rect 48133 6783 48191 6789
rect 48133 6780 48145 6783
rect 48004 6752 48145 6780
rect 48004 6740 48010 6752
rect 48133 6749 48145 6752
rect 48179 6749 48191 6783
rect 48133 6743 48191 6749
rect 2406 6672 2412 6724
rect 2464 6712 2470 6724
rect 3237 6715 3295 6721
rect 3237 6712 3249 6715
rect 2464 6684 3249 6712
rect 2464 6672 2470 6684
rect 3237 6681 3249 6684
rect 3283 6681 3295 6715
rect 3237 6675 3295 6681
rect 32033 6715 32091 6721
rect 32033 6681 32045 6715
rect 32079 6712 32091 6715
rect 32398 6712 32404 6724
rect 32079 6684 32404 6712
rect 32079 6681 32091 6684
rect 32033 6675 32091 6681
rect 32398 6672 32404 6684
rect 32456 6672 32462 6724
rect 42981 6715 43039 6721
rect 42981 6681 42993 6715
rect 43027 6712 43039 6715
rect 43070 6712 43076 6724
rect 43027 6684 43076 6712
rect 43027 6681 43039 6684
rect 42981 6675 43039 6681
rect 43070 6672 43076 6684
rect 43128 6672 43134 6724
rect 46290 6604 46296 6656
rect 46348 6644 46354 6656
rect 46937 6647 46995 6653
rect 46937 6644 46949 6647
rect 46348 6616 46949 6644
rect 46348 6604 46354 6616
rect 46937 6613 46949 6616
rect 46983 6613 46995 6647
rect 47578 6644 47584 6656
rect 47539 6616 47584 6644
rect 46937 6607 46995 6613
rect 47578 6604 47584 6616
rect 47636 6604 47642 6656
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 2406 6440 2412 6452
rect 2367 6412 2412 6440
rect 2406 6400 2412 6412
rect 2464 6400 2470 6452
rect 32398 6440 32404 6452
rect 32359 6412 32404 6440
rect 32398 6400 32404 6412
rect 32456 6400 32462 6452
rect 43070 6440 43076 6452
rect 43031 6412 43076 6440
rect 43070 6400 43076 6412
rect 43128 6400 43134 6452
rect 47302 6372 47308 6384
rect 41386 6344 47308 6372
rect 2498 6304 2504 6316
rect 2459 6276 2504 6304
rect 2498 6264 2504 6276
rect 2556 6264 2562 6316
rect 32493 6307 32551 6313
rect 32493 6273 32505 6307
rect 32539 6304 32551 6307
rect 41386 6304 41414 6344
rect 47302 6332 47308 6344
rect 47360 6332 47366 6384
rect 32539 6276 41414 6304
rect 42981 6307 43039 6313
rect 32539 6273 32551 6276
rect 32493 6267 32551 6273
rect 42981 6273 42993 6307
rect 43027 6304 43039 6307
rect 43070 6304 43076 6316
rect 43027 6276 43076 6304
rect 43027 6273 43039 6276
rect 42981 6267 43039 6273
rect 43070 6264 43076 6276
rect 43128 6264 43134 6316
rect 46382 6304 46388 6316
rect 46343 6276 46388 6304
rect 46382 6264 46388 6276
rect 46440 6264 46446 6316
rect 47210 6304 47216 6316
rect 47123 6276 47216 6304
rect 47210 6264 47216 6276
rect 47268 6304 47274 6316
rect 47762 6304 47768 6316
rect 47268 6276 47348 6304
rect 47723 6276 47768 6304
rect 47268 6264 47274 6276
rect 47320 6248 47348 6276
rect 47762 6264 47768 6276
rect 47820 6264 47826 6316
rect 47302 6196 47308 6248
rect 47360 6196 47366 6248
rect 1857 6103 1915 6109
rect 1857 6069 1869 6103
rect 1903 6100 1915 6103
rect 2958 6100 2964 6112
rect 1903 6072 2964 6100
rect 1903 6069 1915 6072
rect 1857 6063 1915 6069
rect 2958 6060 2964 6072
rect 3016 6060 3022 6112
rect 3145 6103 3203 6109
rect 3145 6069 3157 6103
rect 3191 6100 3203 6103
rect 3418 6100 3424 6112
rect 3191 6072 3424 6100
rect 3191 6069 3203 6072
rect 3145 6063 3203 6069
rect 3418 6060 3424 6072
rect 3476 6060 3482 6112
rect 46477 6103 46535 6109
rect 46477 6069 46489 6103
rect 46523 6100 46535 6103
rect 46934 6100 46940 6112
rect 46523 6072 46940 6100
rect 46523 6069 46535 6072
rect 46477 6063 46535 6069
rect 46934 6060 46940 6072
rect 46992 6060 46998 6112
rect 47026 6060 47032 6112
rect 47084 6100 47090 6112
rect 47121 6103 47179 6109
rect 47121 6100 47133 6103
rect 47084 6072 47133 6100
rect 47084 6060 47090 6072
rect 47121 6069 47133 6072
rect 47167 6069 47179 6103
rect 47121 6063 47179 6069
rect 47857 6103 47915 6109
rect 47857 6069 47869 6103
rect 47903 6100 47915 6103
rect 48130 6100 48136 6112
rect 47903 6072 48136 6100
rect 47903 6069 47915 6072
rect 47857 6063 47915 6069
rect 48130 6060 48136 6072
rect 48188 6060 48194 6112
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 2498 5788 2504 5840
rect 2556 5828 2562 5840
rect 46842 5828 46848 5840
rect 2556 5800 4200 5828
rect 2556 5788 2562 5800
rect 3418 5760 3424 5772
rect 3379 5732 3424 5760
rect 3418 5720 3424 5732
rect 3476 5720 3482 5772
rect 4172 5701 4200 5800
rect 45664 5800 46848 5828
rect 45664 5704 45692 5800
rect 46842 5788 46848 5800
rect 46900 5788 46906 5840
rect 46106 5760 46112 5772
rect 46067 5732 46112 5760
rect 46106 5720 46112 5732
rect 46164 5720 46170 5772
rect 46290 5760 46296 5772
rect 46251 5732 46296 5760
rect 46290 5720 46296 5732
rect 46348 5720 46354 5772
rect 47118 5760 47124 5772
rect 47079 5732 47124 5760
rect 47118 5720 47124 5732
rect 47176 5720 47182 5772
rect 4157 5695 4215 5701
rect 4157 5661 4169 5695
rect 4203 5692 4215 5695
rect 17586 5692 17592 5704
rect 4203 5664 17592 5692
rect 4203 5661 4215 5664
rect 4157 5655 4215 5661
rect 17586 5652 17592 5664
rect 17644 5652 17650 5704
rect 45646 5692 45652 5704
rect 45559 5664 45652 5692
rect 45646 5652 45652 5664
rect 45704 5652 45710 5704
rect 1578 5624 1584 5636
rect 1539 5596 1584 5624
rect 1578 5584 1584 5596
rect 1636 5584 1642 5636
rect 3237 5627 3295 5633
rect 3237 5593 3249 5627
rect 3283 5624 3295 5627
rect 4065 5627 4123 5633
rect 4065 5624 4077 5627
rect 3283 5596 4077 5624
rect 3283 5593 3295 5596
rect 3237 5587 3295 5593
rect 4065 5593 4077 5596
rect 4111 5593 4123 5627
rect 4065 5587 4123 5593
rect 45554 5556 45560 5568
rect 45515 5528 45560 5556
rect 45554 5516 45560 5528
rect 45612 5516 45618 5568
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 47026 5284 47032 5296
rect 46987 5256 47032 5284
rect 47026 5244 47032 5256
rect 47084 5244 47090 5296
rect 4614 5216 4620 5228
rect 4575 5188 4620 5216
rect 4614 5176 4620 5188
rect 4672 5216 4678 5228
rect 12526 5216 12532 5228
rect 4672 5188 12532 5216
rect 4672 5176 4678 5188
rect 12526 5176 12532 5188
rect 12584 5176 12590 5228
rect 2774 5148 2780 5160
rect 2735 5120 2780 5148
rect 2774 5108 2780 5120
rect 2832 5108 2838 5160
rect 3050 5108 3056 5160
rect 3108 5148 3114 5160
rect 3789 5151 3847 5157
rect 3789 5148 3801 5151
rect 3108 5120 3801 5148
rect 3108 5108 3114 5120
rect 3789 5117 3801 5120
rect 3835 5117 3847 5151
rect 3789 5111 3847 5117
rect 3973 5151 4031 5157
rect 3973 5117 3985 5151
rect 4019 5117 4031 5151
rect 3973 5111 4031 5117
rect 46753 5151 46811 5157
rect 46753 5117 46765 5151
rect 46799 5117 46811 5151
rect 47210 5148 47216 5160
rect 47171 5120 47216 5148
rect 46753 5111 46811 5117
rect 2498 5040 2504 5092
rect 2556 5080 2562 5092
rect 3988 5080 4016 5111
rect 2556 5052 4016 5080
rect 46768 5080 46796 5111
rect 47210 5108 47216 5120
rect 47268 5108 47274 5160
rect 48406 5080 48412 5092
rect 46768 5052 48412 5080
rect 2556 5040 2562 5052
rect 48406 5040 48412 5052
rect 48464 5040 48470 5092
rect 4525 5015 4583 5021
rect 4525 4981 4537 5015
rect 4571 5012 4583 5015
rect 4798 5012 4804 5024
rect 4571 4984 4804 5012
rect 4571 4981 4583 4984
rect 4525 4975 4583 4981
rect 4798 4972 4804 4984
rect 4856 4972 4862 5024
rect 44726 5012 44732 5024
rect 44687 4984 44732 5012
rect 44726 4972 44732 4984
rect 44784 4972 44790 5024
rect 47949 5015 48007 5021
rect 47949 4981 47961 5015
rect 47995 5012 48007 5015
rect 48314 5012 48320 5024
rect 47995 4984 48320 5012
rect 47995 4981 48007 4984
rect 47949 4975 48007 4981
rect 48314 4972 48320 4984
rect 48372 4972 48378 5024
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 2498 4808 2504 4820
rect 2459 4780 2504 4808
rect 2498 4768 2504 4780
rect 2556 4768 2562 4820
rect 3050 4808 3056 4820
rect 3011 4780 3056 4808
rect 3050 4768 3056 4780
rect 3108 4768 3114 4820
rect 1765 4743 1823 4749
rect 1765 4709 1777 4743
rect 1811 4740 1823 4743
rect 47762 4740 47768 4752
rect 1811 4712 6914 4740
rect 1811 4709 1823 4712
rect 1765 4703 1823 4709
rect 6886 4672 6914 4712
rect 45204 4712 47768 4740
rect 18230 4672 18236 4684
rect 6886 4644 18236 4672
rect 18230 4632 18236 4644
rect 18288 4632 18294 4684
rect 1302 4564 1308 4616
rect 1360 4604 1366 4616
rect 1581 4607 1639 4613
rect 1581 4604 1593 4607
rect 1360 4576 1593 4604
rect 1360 4564 1366 4576
rect 1581 4573 1593 4576
rect 1627 4573 1639 4607
rect 1581 4567 1639 4573
rect 2961 4607 3019 4613
rect 2961 4573 2973 4607
rect 3007 4604 3019 4607
rect 3234 4604 3240 4616
rect 3007 4576 3240 4604
rect 3007 4573 3019 4576
rect 2961 4567 3019 4573
rect 3234 4564 3240 4576
rect 3292 4604 3298 4616
rect 4062 4604 4068 4616
rect 3292 4576 4068 4604
rect 3292 4564 3298 4576
rect 4062 4564 4068 4576
rect 4120 4564 4126 4616
rect 4157 4607 4215 4613
rect 4157 4573 4169 4607
rect 4203 4573 4215 4607
rect 4157 4567 4215 4573
rect 4617 4607 4675 4613
rect 4617 4573 4629 4607
rect 4663 4604 4675 4607
rect 4706 4604 4712 4616
rect 4663 4576 4712 4604
rect 4663 4573 4675 4576
rect 4617 4567 4675 4573
rect 4172 4536 4200 4567
rect 4706 4564 4712 4576
rect 4764 4564 4770 4616
rect 5442 4604 5448 4616
rect 5403 4576 5448 4604
rect 5442 4564 5448 4576
rect 5500 4604 5506 4616
rect 24854 4604 24860 4616
rect 5500 4576 24860 4604
rect 5500 4564 5506 4576
rect 24854 4564 24860 4576
rect 24912 4564 24918 4616
rect 39022 4604 39028 4616
rect 38983 4576 39028 4604
rect 39022 4564 39028 4576
rect 39080 4564 39086 4616
rect 43070 4604 43076 4616
rect 43031 4576 43076 4604
rect 43070 4564 43076 4576
rect 43128 4564 43134 4616
rect 43901 4607 43959 4613
rect 43901 4573 43913 4607
rect 43947 4604 43959 4607
rect 44358 4604 44364 4616
rect 43947 4576 44364 4604
rect 43947 4573 43959 4576
rect 43901 4567 43959 4573
rect 44358 4564 44364 4576
rect 44416 4564 44422 4616
rect 44542 4604 44548 4616
rect 44503 4576 44548 4604
rect 44542 4564 44548 4576
rect 44600 4564 44606 4616
rect 45204 4613 45232 4712
rect 47762 4700 47768 4712
rect 47820 4700 47826 4752
rect 46842 4672 46848 4684
rect 46803 4644 46848 4672
rect 46842 4632 46848 4644
rect 46900 4632 46906 4684
rect 48130 4672 48136 4684
rect 48091 4644 48136 4672
rect 48130 4632 48136 4644
rect 48188 4632 48194 4684
rect 48314 4672 48320 4684
rect 48275 4644 48320 4672
rect 48314 4632 48320 4644
rect 48372 4632 48378 4684
rect 45189 4607 45247 4613
rect 45189 4573 45201 4607
rect 45235 4573 45247 4607
rect 45189 4567 45247 4573
rect 46017 4607 46075 4613
rect 46017 4573 46029 4607
rect 46063 4604 46075 4607
rect 46750 4604 46756 4616
rect 46063 4576 46756 4604
rect 46063 4573 46075 4576
rect 46017 4567 46075 4573
rect 46750 4564 46756 4576
rect 46808 4564 46814 4616
rect 4982 4536 4988 4548
rect 4172 4508 4988 4536
rect 4982 4496 4988 4508
rect 5040 4536 5046 4548
rect 19426 4536 19432 4548
rect 5040 4508 19432 4536
rect 5040 4496 5046 4508
rect 19426 4496 19432 4508
rect 19484 4496 19490 4548
rect 3510 4428 3516 4480
rect 3568 4468 3574 4480
rect 4065 4471 4123 4477
rect 4065 4468 4077 4471
rect 3568 4440 4077 4468
rect 3568 4428 3574 4440
rect 4065 4437 4077 4440
rect 4111 4437 4123 4471
rect 5350 4468 5356 4480
rect 5311 4440 5356 4468
rect 4065 4431 4123 4437
rect 5350 4428 5356 4440
rect 5408 4428 5414 4480
rect 43165 4471 43223 4477
rect 43165 4437 43177 4471
rect 43211 4468 43223 4471
rect 45094 4468 45100 4480
rect 43211 4440 45100 4468
rect 43211 4437 43223 4440
rect 43165 4431 43223 4437
rect 45094 4428 45100 4440
rect 45152 4428 45158 4480
rect 45281 4471 45339 4477
rect 45281 4437 45293 4471
rect 45327 4468 45339 4471
rect 45370 4468 45376 4480
rect 45327 4440 45376 4468
rect 45327 4437 45339 4440
rect 45281 4431 45339 4437
rect 45370 4428 45376 4440
rect 45428 4428 45434 4480
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 1673 4199 1731 4205
rect 1673 4165 1685 4199
rect 1719 4196 1731 4199
rect 2774 4196 2780 4208
rect 1719 4168 2780 4196
rect 1719 4165 1731 4168
rect 1673 4159 1731 4165
rect 2774 4156 2780 4168
rect 2832 4156 2838 4208
rect 44269 4199 44327 4205
rect 5644 4168 6776 4196
rect 4062 4128 4068 4140
rect 3975 4100 4068 4128
rect 4062 4088 4068 4100
rect 4120 4128 4126 4140
rect 5644 4128 5672 4168
rect 5810 4128 5816 4140
rect 4120 4100 5672 4128
rect 5771 4100 5816 4128
rect 4120 4088 4126 4100
rect 5810 4088 5816 4100
rect 5868 4128 5874 4140
rect 6641 4131 6699 4137
rect 6641 4128 6653 4131
rect 5868 4100 6653 4128
rect 5868 4088 5874 4100
rect 6641 4097 6653 4100
rect 6687 4097 6699 4131
rect 6748 4128 6776 4168
rect 44269 4165 44281 4199
rect 44315 4196 44327 4199
rect 44315 4168 44496 4196
rect 44315 4165 44327 4168
rect 44269 4159 44327 4165
rect 7558 4128 7564 4140
rect 6748 4100 7420 4128
rect 7519 4100 7564 4128
rect 6641 4091 6699 4097
rect 6656 4060 6684 4091
rect 7392 4060 7420 4100
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 10505 4131 10563 4137
rect 10505 4097 10517 4131
rect 10551 4097 10563 4131
rect 12526 4128 12532 4140
rect 12487 4100 12532 4128
rect 10505 4091 10563 4097
rect 10520 4060 10548 4091
rect 12526 4088 12532 4100
rect 12584 4088 12590 4140
rect 13170 4128 13176 4140
rect 13131 4100 13176 4128
rect 13170 4088 13176 4100
rect 13228 4088 13234 4140
rect 18601 4131 18659 4137
rect 18601 4097 18613 4131
rect 18647 4097 18659 4131
rect 18601 4091 18659 4097
rect 26145 4131 26203 4137
rect 26145 4097 26157 4131
rect 26191 4128 26203 4131
rect 27154 4128 27160 4140
rect 26191 4100 26225 4128
rect 27115 4100 27160 4128
rect 26191 4097 26203 4100
rect 26145 4091 26203 4097
rect 6656 4032 7328 4060
rect 7392 4032 10548 4060
rect 1949 3995 2007 4001
rect 1949 3961 1961 3995
rect 1995 3992 2007 3995
rect 7190 3992 7196 4004
rect 1995 3964 7196 3992
rect 1995 3961 2007 3964
rect 1949 3955 2007 3961
rect 7190 3952 7196 3964
rect 7248 3952 7254 4004
rect 7300 3992 7328 4032
rect 18616 3992 18644 4091
rect 24854 4020 24860 4072
rect 24912 4060 24918 4072
rect 26160 4060 26188 4091
rect 27154 4088 27160 4100
rect 27212 4088 27218 4140
rect 38378 4128 38384 4140
rect 38339 4100 38384 4128
rect 38378 4088 38384 4100
rect 38436 4088 38442 4140
rect 39022 4128 39028 4140
rect 38983 4100 39028 4128
rect 39022 4088 39028 4100
rect 39080 4088 39086 4140
rect 41509 4131 41567 4137
rect 41509 4097 41521 4131
rect 41555 4128 41567 4131
rect 41966 4128 41972 4140
rect 41555 4100 41972 4128
rect 41555 4097 41567 4100
rect 41509 4091 41567 4097
rect 41966 4088 41972 4100
rect 42024 4088 42030 4140
rect 44468 4128 44496 4168
rect 44468 4100 44588 4128
rect 24912 4032 26234 4060
rect 24912 4020 24918 4032
rect 7300 3964 18644 3992
rect 18693 3995 18751 4001
rect 18693 3961 18705 3995
rect 18739 3992 18751 3995
rect 20162 3992 20168 4004
rect 18739 3964 20168 3992
rect 18739 3961 18751 3964
rect 18693 3955 18751 3961
rect 20162 3952 20168 3964
rect 20220 3952 20226 4004
rect 26206 3992 26234 4032
rect 38194 4020 38200 4072
rect 38252 4060 38258 4072
rect 39209 4063 39267 4069
rect 39209 4060 39221 4063
rect 38252 4032 39221 4060
rect 38252 4020 38258 4032
rect 39209 4029 39221 4032
rect 39255 4029 39267 4063
rect 40494 4060 40500 4072
rect 40455 4032 40500 4060
rect 39209 4023 39267 4029
rect 40494 4020 40500 4032
rect 40552 4020 40558 4072
rect 43993 4063 44051 4069
rect 43993 4029 44005 4063
rect 44039 4060 44051 4063
rect 44174 4060 44180 4072
rect 44039 4032 44180 4060
rect 44039 4029 44051 4032
rect 43993 4023 44051 4029
rect 44174 4020 44180 4032
rect 44232 4020 44238 4072
rect 44453 4063 44511 4069
rect 44453 4029 44465 4063
rect 44499 4029 44511 4063
rect 44453 4023 44511 4029
rect 38102 3992 38108 4004
rect 26206 3964 38108 3992
rect 38102 3952 38108 3964
rect 38160 3952 38166 4004
rect 38378 3952 38384 4004
rect 38436 3992 38442 4004
rect 44082 3992 44088 4004
rect 38436 3964 44088 3992
rect 38436 3952 38442 3964
rect 44082 3952 44088 3964
rect 44140 3952 44146 4004
rect 3053 3927 3111 3933
rect 3053 3893 3065 3927
rect 3099 3924 3111 3927
rect 3694 3924 3700 3936
rect 3099 3896 3700 3924
rect 3099 3893 3111 3896
rect 3053 3887 3111 3893
rect 3694 3884 3700 3896
rect 3752 3884 3758 3936
rect 4157 3927 4215 3933
rect 4157 3893 4169 3927
rect 4203 3924 4215 3927
rect 4614 3924 4620 3936
rect 4203 3896 4620 3924
rect 4203 3893 4215 3896
rect 4157 3887 4215 3893
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 4982 3924 4988 3936
rect 4943 3896 4988 3924
rect 4982 3884 4988 3896
rect 5040 3884 5046 3936
rect 5905 3927 5963 3933
rect 5905 3893 5917 3927
rect 5951 3924 5963 3927
rect 6086 3924 6092 3936
rect 5951 3896 6092 3924
rect 5951 3893 5963 3896
rect 5905 3887 5963 3893
rect 6086 3884 6092 3896
rect 6144 3884 6150 3936
rect 6733 3927 6791 3933
rect 6733 3893 6745 3927
rect 6779 3924 6791 3927
rect 6822 3924 6828 3936
rect 6779 3896 6828 3924
rect 6779 3893 6791 3896
rect 6733 3887 6791 3893
rect 6822 3884 6828 3896
rect 6880 3884 6886 3936
rect 7650 3924 7656 3936
rect 7611 3896 7656 3924
rect 7650 3884 7656 3896
rect 7708 3884 7714 3936
rect 10597 3927 10655 3933
rect 10597 3893 10609 3927
rect 10643 3924 10655 3927
rect 10686 3924 10692 3936
rect 10643 3896 10692 3924
rect 10643 3893 10655 3896
rect 10597 3887 10655 3893
rect 10686 3884 10692 3896
rect 10744 3884 10750 3936
rect 12437 3927 12495 3933
rect 12437 3893 12449 3927
rect 12483 3924 12495 3927
rect 12526 3924 12532 3936
rect 12483 3896 12532 3924
rect 12483 3893 12495 3896
rect 12437 3887 12495 3893
rect 12526 3884 12532 3896
rect 12584 3884 12590 3936
rect 13265 3927 13323 3933
rect 13265 3893 13277 3927
rect 13311 3924 13323 3927
rect 13354 3924 13360 3936
rect 13311 3896 13360 3924
rect 13311 3893 13323 3896
rect 13265 3887 13323 3893
rect 13354 3884 13360 3896
rect 13412 3884 13418 3936
rect 20070 3924 20076 3936
rect 20031 3896 20076 3924
rect 20070 3884 20076 3896
rect 20128 3884 20134 3936
rect 24762 3884 24768 3936
rect 24820 3924 24826 3936
rect 25317 3927 25375 3933
rect 25317 3924 25329 3927
rect 24820 3896 25329 3924
rect 24820 3884 24826 3896
rect 25317 3893 25329 3896
rect 25363 3893 25375 3927
rect 25317 3887 25375 3893
rect 25958 3884 25964 3936
rect 26016 3924 26022 3936
rect 26053 3927 26111 3933
rect 26053 3924 26065 3927
rect 26016 3896 26065 3924
rect 26016 3884 26022 3896
rect 26053 3893 26065 3896
rect 26099 3893 26111 3927
rect 26053 3887 26111 3893
rect 27249 3927 27307 3933
rect 27249 3893 27261 3927
rect 27295 3924 27307 3927
rect 27338 3924 27344 3936
rect 27295 3896 27344 3924
rect 27295 3893 27307 3896
rect 27249 3887 27307 3893
rect 27338 3884 27344 3896
rect 27396 3884 27402 3936
rect 38473 3927 38531 3933
rect 38473 3893 38485 3927
rect 38519 3924 38531 3927
rect 38930 3924 38936 3936
rect 38519 3896 38936 3924
rect 38519 3893 38531 3896
rect 38473 3887 38531 3893
rect 38930 3884 38936 3896
rect 38988 3884 38994 3936
rect 40770 3884 40776 3936
rect 40828 3924 40834 3936
rect 41417 3927 41475 3933
rect 41417 3924 41429 3927
rect 40828 3896 41429 3924
rect 40828 3884 40834 3896
rect 41417 3893 41429 3896
rect 41463 3893 41475 3927
rect 44468 3924 44496 4023
rect 44560 3992 44588 4100
rect 46750 4088 46756 4140
rect 46808 4128 46814 4140
rect 46808 4100 46853 4128
rect 46808 4088 46814 4100
rect 47210 4088 47216 4140
rect 47268 4128 47274 4140
rect 47765 4131 47823 4137
rect 47765 4128 47777 4131
rect 47268 4100 47777 4128
rect 47268 4088 47274 4100
rect 47765 4097 47777 4100
rect 47811 4097 47823 4131
rect 47765 4091 47823 4097
rect 45738 4060 45744 4072
rect 45699 4032 45744 4060
rect 45738 4020 45744 4032
rect 45796 4020 45802 4072
rect 46569 4063 46627 4069
rect 46569 4029 46581 4063
rect 46615 4060 46627 4063
rect 47854 4060 47860 4072
rect 46615 4032 47860 4060
rect 46615 4029 46627 4032
rect 46569 4023 46627 4029
rect 47854 4020 47860 4032
rect 47912 4020 47918 4072
rect 47578 3992 47584 4004
rect 44560 3964 47584 3992
rect 47578 3952 47584 3964
rect 47636 3952 47642 4004
rect 47946 3924 47952 3936
rect 44468 3896 47952 3924
rect 41417 3887 41475 3893
rect 47946 3884 47952 3896
rect 48004 3884 48010 3936
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 7190 3680 7196 3732
rect 7248 3720 7254 3732
rect 12802 3720 12808 3732
rect 7248 3692 12808 3720
rect 7248 3680 7254 3692
rect 12802 3680 12808 3692
rect 12860 3680 12866 3732
rect 27154 3720 27160 3732
rect 26206 3692 27160 3720
rect 4798 3652 4804 3664
rect 3252 3624 4804 3652
rect 3252 3593 3280 3624
rect 4798 3612 4804 3624
rect 4856 3612 4862 3664
rect 4890 3612 4896 3664
rect 4948 3652 4954 3664
rect 13170 3652 13176 3664
rect 4948 3624 13176 3652
rect 4948 3612 4954 3624
rect 13170 3612 13176 3624
rect 13228 3612 13234 3664
rect 17586 3612 17592 3664
rect 17644 3652 17650 3664
rect 26206 3652 26234 3692
rect 27154 3680 27160 3692
rect 27212 3720 27218 3732
rect 43070 3720 43076 3732
rect 27212 3692 43076 3720
rect 27212 3680 27218 3692
rect 43070 3680 43076 3692
rect 43128 3680 43134 3732
rect 44082 3680 44088 3732
rect 44140 3720 44146 3732
rect 47302 3720 47308 3732
rect 44140 3692 47308 3720
rect 44140 3680 44146 3692
rect 47302 3680 47308 3692
rect 47360 3680 47366 3732
rect 17644 3624 26234 3652
rect 17644 3612 17650 3624
rect 30282 3612 30288 3664
rect 30340 3652 30346 3664
rect 38194 3652 38200 3664
rect 30340 3624 33548 3652
rect 38155 3624 38200 3652
rect 30340 3612 30346 3624
rect 3237 3587 3295 3593
rect 3237 3553 3249 3587
rect 3283 3553 3295 3587
rect 3237 3547 3295 3553
rect 3421 3587 3479 3593
rect 3421 3553 3433 3587
rect 3467 3584 3479 3587
rect 4706 3584 4712 3596
rect 3467 3556 4712 3584
rect 3467 3553 3479 3556
rect 3421 3547 3479 3553
rect 4706 3544 4712 3556
rect 4764 3544 4770 3596
rect 6086 3584 6092 3596
rect 6047 3556 6092 3584
rect 6086 3544 6092 3556
rect 6144 3544 6150 3596
rect 6454 3584 6460 3596
rect 6415 3556 6460 3584
rect 6454 3544 6460 3556
rect 6512 3544 6518 3596
rect 10686 3584 10692 3596
rect 10647 3556 10692 3584
rect 10686 3544 10692 3556
rect 10744 3544 10750 3596
rect 10962 3584 10968 3596
rect 10923 3556 10968 3584
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 25958 3584 25964 3596
rect 25919 3556 25964 3584
rect 25958 3544 25964 3556
rect 26016 3544 26022 3596
rect 26418 3584 26424 3596
rect 26379 3556 26424 3584
rect 26418 3544 26424 3556
rect 26476 3544 26482 3596
rect 1578 3516 1584 3528
rect 1539 3488 1584 3516
rect 1578 3476 1584 3488
rect 1636 3476 1642 3528
rect 4154 3516 4160 3528
rect 4115 3488 4160 3516
rect 4154 3476 4160 3488
rect 4212 3476 4218 3528
rect 4801 3519 4859 3525
rect 4801 3485 4813 3519
rect 4847 3516 4859 3519
rect 4890 3516 4896 3528
rect 4847 3488 4896 3516
rect 4847 3485 4859 3488
rect 4801 3479 4859 3485
rect 4890 3476 4896 3488
rect 4948 3476 4954 3528
rect 5445 3519 5503 3525
rect 5445 3485 5457 3519
rect 5491 3516 5503 3519
rect 5905 3519 5963 3525
rect 5905 3516 5917 3519
rect 5491 3488 5917 3516
rect 5491 3485 5503 3488
rect 5445 3479 5503 3485
rect 5905 3485 5917 3488
rect 5951 3485 5963 3519
rect 5905 3479 5963 3485
rect 7466 3476 7472 3528
rect 7524 3516 7530 3528
rect 8205 3519 8263 3525
rect 8205 3516 8217 3519
rect 7524 3488 8217 3516
rect 7524 3476 7530 3488
rect 8205 3485 8217 3488
rect 8251 3485 8263 3519
rect 10502 3516 10508 3528
rect 10463 3488 10508 3516
rect 8205 3479 8263 3485
rect 10502 3476 10508 3488
rect 10560 3476 10566 3528
rect 13170 3516 13176 3528
rect 13131 3488 13176 3516
rect 13170 3476 13176 3488
rect 13228 3476 13234 3528
rect 16850 3476 16856 3528
rect 16908 3516 16914 3528
rect 16945 3519 17003 3525
rect 16945 3516 16957 3519
rect 16908 3488 16957 3516
rect 16908 3476 16914 3488
rect 16945 3485 16957 3488
rect 16991 3485 17003 3519
rect 17586 3516 17592 3528
rect 17547 3488 17592 3516
rect 16945 3479 17003 3485
rect 17586 3476 17592 3488
rect 17644 3476 17650 3528
rect 18877 3519 18935 3525
rect 18877 3485 18889 3519
rect 18923 3516 18935 3519
rect 19334 3516 19340 3528
rect 18923 3488 19340 3516
rect 18923 3485 18935 3488
rect 18877 3479 18935 3485
rect 19334 3476 19340 3488
rect 19392 3476 19398 3528
rect 19426 3476 19432 3528
rect 19484 3516 19490 3528
rect 19484 3488 19529 3516
rect 19484 3476 19490 3488
rect 19978 3476 19984 3528
rect 20036 3516 20042 3528
rect 20073 3519 20131 3525
rect 20073 3516 20085 3519
rect 20036 3488 20085 3516
rect 20036 3476 20042 3488
rect 20073 3485 20085 3488
rect 20119 3485 20131 3519
rect 20073 3479 20131 3485
rect 25317 3519 25375 3525
rect 25317 3485 25329 3519
rect 25363 3516 25375 3519
rect 25777 3519 25835 3525
rect 25777 3516 25789 3519
rect 25363 3488 25789 3516
rect 25363 3485 25375 3488
rect 25317 3479 25375 3485
rect 25777 3485 25789 3488
rect 25823 3485 25835 3519
rect 25777 3479 25835 3485
rect 27154 3476 27160 3528
rect 27212 3516 27218 3528
rect 28077 3519 28135 3525
rect 28077 3516 28089 3519
rect 27212 3488 28089 3516
rect 27212 3476 27218 3488
rect 28077 3485 28089 3488
rect 28123 3485 28135 3519
rect 28077 3479 28135 3485
rect 20349 3451 20407 3457
rect 20349 3417 20361 3451
rect 20395 3448 20407 3451
rect 33318 3448 33324 3460
rect 20395 3420 33324 3448
rect 20395 3417 20407 3420
rect 20349 3411 20407 3417
rect 33318 3408 33324 3420
rect 33376 3408 33382 3460
rect 33520 3448 33548 3624
rect 38194 3612 38200 3624
rect 38252 3612 38258 3664
rect 44177 3655 44235 3661
rect 44177 3652 44189 3655
rect 38304 3624 44189 3652
rect 34054 3544 34060 3596
rect 34112 3584 34118 3596
rect 38304 3584 38332 3624
rect 44177 3621 44189 3624
rect 44223 3621 44235 3655
rect 44177 3615 44235 3621
rect 45278 3612 45284 3664
rect 45336 3652 45342 3664
rect 45336 3624 45692 3652
rect 45336 3612 45342 3624
rect 40770 3584 40776 3596
rect 34112 3556 38332 3584
rect 40731 3556 40776 3584
rect 34112 3544 34118 3556
rect 40770 3544 40776 3556
rect 40828 3544 40834 3596
rect 41230 3584 41236 3596
rect 41191 3556 41236 3584
rect 41230 3544 41236 3556
rect 41288 3544 41294 3596
rect 44542 3544 44548 3596
rect 44600 3584 44606 3596
rect 45189 3587 45247 3593
rect 45189 3584 45201 3587
rect 44600 3556 45201 3584
rect 44600 3544 44606 3556
rect 45189 3553 45201 3556
rect 45235 3553 45247 3587
rect 45370 3584 45376 3596
rect 45331 3556 45376 3584
rect 45189 3547 45247 3553
rect 45370 3544 45376 3556
rect 45428 3544 45434 3596
rect 45664 3593 45692 3624
rect 45649 3587 45707 3593
rect 45649 3553 45661 3587
rect 45695 3553 45707 3587
rect 45649 3547 45707 3553
rect 38102 3516 38108 3528
rect 38063 3488 38108 3516
rect 38102 3476 38108 3488
rect 38160 3476 38166 3528
rect 38746 3516 38752 3528
rect 38707 3488 38752 3516
rect 38746 3476 38752 3488
rect 38804 3476 38810 3528
rect 40586 3516 40592 3528
rect 40547 3488 40592 3516
rect 40586 3476 40592 3488
rect 40644 3476 40650 3528
rect 41966 3476 41972 3528
rect 42024 3516 42030 3528
rect 43073 3519 43131 3525
rect 43073 3516 43085 3519
rect 42024 3488 43085 3516
rect 42024 3476 42030 3488
rect 43073 3485 43085 3488
rect 43119 3516 43131 3519
rect 48314 3516 48320 3528
rect 43119 3488 44312 3516
rect 48275 3488 48320 3516
rect 43119 3485 43131 3488
rect 43073 3479 43131 3485
rect 33520 3420 43760 3448
rect 4338 3340 4344 3392
rect 4396 3380 4402 3392
rect 4709 3383 4767 3389
rect 4709 3380 4721 3383
rect 4396 3352 4721 3380
rect 4396 3340 4402 3352
rect 4709 3349 4721 3352
rect 4755 3349 4767 3383
rect 4709 3343 4767 3349
rect 17034 3340 17040 3392
rect 17092 3380 17098 3392
rect 17497 3383 17555 3389
rect 17497 3380 17509 3383
rect 17092 3352 17509 3380
rect 17092 3340 17098 3352
rect 17497 3349 17509 3352
rect 17543 3349 17555 3383
rect 17497 3343 17555 3349
rect 19426 3340 19432 3392
rect 19484 3380 19490 3392
rect 19521 3383 19579 3389
rect 19521 3380 19533 3383
rect 19484 3352 19533 3380
rect 19484 3340 19490 3352
rect 19521 3349 19533 3352
rect 19567 3349 19579 3383
rect 19521 3343 19579 3349
rect 42794 3340 42800 3392
rect 42852 3380 42858 3392
rect 42981 3383 43039 3389
rect 42981 3380 42993 3383
rect 42852 3352 42993 3380
rect 42852 3340 42858 3352
rect 42981 3349 42993 3352
rect 43027 3349 43039 3383
rect 43732 3380 43760 3420
rect 43806 3408 43812 3460
rect 43864 3448 43870 3460
rect 43993 3451 44051 3457
rect 43993 3448 44005 3451
rect 43864 3420 44005 3448
rect 43864 3408 43870 3420
rect 43993 3417 44005 3420
rect 44039 3417 44051 3451
rect 44284 3448 44312 3488
rect 48314 3476 48320 3488
rect 48372 3476 48378 3528
rect 45646 3448 45652 3460
rect 44284 3420 45652 3448
rect 43993 3411 44051 3417
rect 45646 3408 45652 3420
rect 45704 3408 45710 3460
rect 48133 3383 48191 3389
rect 48133 3380 48145 3383
rect 43732 3352 48145 3380
rect 42981 3343 43039 3349
rect 48133 3349 48145 3352
rect 48179 3349 48191 3383
rect 48133 3343 48191 3349
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 47854 3176 47860 3188
rect 47815 3148 47860 3176
rect 47854 3136 47860 3148
rect 47912 3136 47918 3188
rect 3510 3108 3516 3120
rect 3471 3080 3516 3108
rect 3510 3068 3516 3080
rect 3568 3068 3574 3120
rect 4338 3108 4344 3120
rect 4299 3080 4344 3108
rect 4338 3068 4344 3080
rect 4396 3068 4402 3120
rect 7650 3108 7656 3120
rect 7611 3080 7656 3108
rect 7650 3068 7656 3080
rect 7708 3068 7714 3120
rect 13354 3108 13360 3120
rect 13315 3080 13360 3108
rect 13354 3068 13360 3080
rect 13412 3068 13418 3120
rect 17034 3108 17040 3120
rect 16995 3080 17040 3108
rect 17034 3068 17040 3080
rect 17092 3068 17098 3120
rect 19426 3068 19432 3120
rect 19484 3108 19490 3120
rect 19797 3111 19855 3117
rect 19797 3108 19809 3111
rect 19484 3080 19809 3108
rect 19484 3068 19490 3080
rect 19797 3077 19809 3080
rect 19843 3077 19855 3111
rect 27338 3108 27344 3120
rect 27299 3080 27344 3108
rect 19797 3071 19855 3077
rect 27338 3068 27344 3080
rect 27396 3068 27402 3120
rect 38930 3108 38936 3120
rect 38891 3080 38936 3108
rect 38930 3068 38936 3080
rect 38988 3068 38994 3120
rect 42794 3108 42800 3120
rect 42755 3080 42800 3108
rect 42794 3068 42800 3080
rect 42852 3068 42858 3120
rect 45094 3108 45100 3120
rect 45055 3080 45100 3108
rect 45094 3068 45100 3080
rect 45152 3068 45158 3120
rect 3694 3000 3700 3052
rect 3752 3040 3758 3052
rect 7466 3040 7472 3052
rect 3752 3012 3797 3040
rect 7427 3012 7472 3040
rect 3752 3000 3758 3012
rect 7466 3000 7472 3012
rect 7524 3000 7530 3052
rect 10502 3040 10508 3052
rect 10463 3012 10508 3040
rect 10502 3000 10508 3012
rect 10560 3000 10566 3052
rect 11606 3000 11612 3052
rect 11664 3040 11670 3052
rect 11701 3043 11759 3049
rect 11701 3040 11713 3043
rect 11664 3012 11713 3040
rect 11664 3000 11670 3012
rect 11701 3009 11713 3012
rect 11747 3009 11759 3043
rect 13170 3040 13176 3052
rect 13131 3012 13176 3040
rect 11701 3003 11759 3009
rect 13170 3000 13176 3012
rect 13228 3000 13234 3052
rect 16850 3040 16856 3052
rect 16811 3012 16856 3040
rect 16850 3000 16856 3012
rect 16908 3000 16914 3052
rect 24762 3040 24768 3052
rect 24723 3012 24768 3040
rect 24762 3000 24768 3012
rect 24820 3000 24826 3052
rect 27154 3040 27160 3052
rect 27115 3012 27160 3040
rect 27154 3000 27160 3012
rect 27212 3000 27218 3052
rect 38746 3040 38752 3052
rect 38707 3012 38752 3040
rect 38746 3000 38752 3012
rect 38804 3000 38810 3052
rect 40586 3000 40592 3052
rect 40644 3040 40650 3052
rect 41049 3043 41107 3049
rect 41049 3040 41061 3043
rect 40644 3012 41061 3040
rect 40644 3000 40650 3012
rect 41049 3009 41061 3012
rect 41095 3009 41107 3043
rect 41049 3003 41107 3009
rect 44358 3000 44364 3052
rect 44416 3040 44422 3052
rect 44913 3043 44971 3049
rect 44913 3040 44925 3043
rect 44416 3012 44925 3040
rect 44416 3000 44422 3012
rect 44913 3009 44925 3012
rect 44959 3009 44971 3043
rect 44913 3003 44971 3009
rect 46290 3000 46296 3052
rect 46348 3040 46354 3052
rect 47765 3043 47823 3049
rect 47765 3040 47777 3043
rect 46348 3012 47777 3040
rect 46348 3000 46354 3012
rect 47765 3009 47777 3012
rect 47811 3009 47823 3043
rect 47765 3003 47823 3009
rect 3234 2972 3240 2984
rect 3195 2944 3240 2972
rect 3234 2932 3240 2944
rect 3292 2932 3298 2984
rect 4157 2975 4215 2981
rect 4157 2941 4169 2975
rect 4203 2972 4215 2975
rect 4982 2972 4988 2984
rect 4203 2944 4988 2972
rect 4203 2941 4215 2944
rect 4157 2935 4215 2941
rect 4982 2932 4988 2944
rect 5040 2932 5046 2984
rect 5166 2972 5172 2984
rect 5127 2944 5172 2972
rect 5166 2932 5172 2944
rect 5224 2932 5230 2984
rect 7742 2932 7748 2984
rect 7800 2972 7806 2984
rect 7929 2975 7987 2981
rect 7929 2972 7941 2975
rect 7800 2944 7941 2972
rect 7800 2932 7806 2944
rect 7929 2941 7941 2944
rect 7975 2941 7987 2975
rect 7929 2935 7987 2941
rect 13538 2932 13544 2984
rect 13596 2972 13602 2984
rect 13633 2975 13691 2981
rect 13633 2972 13645 2975
rect 13596 2944 13645 2972
rect 13596 2932 13602 2944
rect 13633 2941 13645 2944
rect 13679 2941 13691 2975
rect 17402 2972 17408 2984
rect 17363 2944 17408 2972
rect 13633 2935 13691 2941
rect 17402 2932 17408 2944
rect 17460 2932 17466 2984
rect 19613 2975 19671 2981
rect 19613 2941 19625 2975
rect 19659 2972 19671 2975
rect 20070 2972 20076 2984
rect 19659 2944 20076 2972
rect 19659 2941 19671 2944
rect 19613 2935 19671 2941
rect 20070 2932 20076 2944
rect 20128 2932 20134 2984
rect 20622 2972 20628 2984
rect 20583 2944 20628 2972
rect 20622 2932 20628 2944
rect 20680 2932 20686 2984
rect 24946 2972 24952 2984
rect 24907 2944 24952 2972
rect 24946 2932 24952 2944
rect 25004 2932 25010 2984
rect 25774 2972 25780 2984
rect 25735 2944 25780 2972
rect 25774 2932 25780 2944
rect 25832 2932 25838 2984
rect 27706 2972 27712 2984
rect 27667 2944 27712 2972
rect 27706 2932 27712 2944
rect 27764 2932 27770 2984
rect 39298 2972 39304 2984
rect 39259 2944 39304 2972
rect 39298 2932 39304 2944
rect 39356 2932 39362 2984
rect 41877 2975 41935 2981
rect 41877 2941 41889 2975
rect 41923 2972 41935 2975
rect 42613 2975 42671 2981
rect 42613 2972 42625 2975
rect 41923 2944 42625 2972
rect 41923 2941 41935 2944
rect 41877 2935 41935 2941
rect 42613 2941 42625 2944
rect 42659 2941 42671 2975
rect 42613 2935 42671 2941
rect 43073 2975 43131 2981
rect 43073 2941 43085 2975
rect 43119 2941 43131 2975
rect 46750 2972 46756 2984
rect 46711 2944 46756 2972
rect 43073 2935 43131 2941
rect 11885 2907 11943 2913
rect 11885 2873 11897 2907
rect 11931 2904 11943 2907
rect 23566 2904 23572 2916
rect 11931 2876 23572 2904
rect 11931 2873 11943 2876
rect 11885 2867 11943 2873
rect 23566 2864 23572 2876
rect 23624 2864 23630 2916
rect 6638 2836 6644 2848
rect 6599 2808 6644 2836
rect 6638 2796 6644 2808
rect 6696 2796 6702 2848
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 12492 2808 12537 2836
rect 12492 2796 12498 2808
rect 41874 2796 41880 2848
rect 41932 2836 41938 2848
rect 43088 2836 43116 2935
rect 46750 2932 46756 2944
rect 46808 2932 46814 2984
rect 41932 2808 43116 2836
rect 41932 2796 41938 2808
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 12618 2592 12624 2644
rect 12676 2632 12682 2644
rect 14461 2635 14519 2641
rect 14461 2632 14473 2635
rect 12676 2604 14473 2632
rect 12676 2592 12682 2604
rect 14461 2601 14473 2604
rect 14507 2601 14519 2635
rect 14461 2595 14519 2601
rect 24946 2592 24952 2644
rect 25004 2632 25010 2644
rect 25409 2635 25467 2641
rect 25409 2632 25421 2635
rect 25004 2604 25421 2632
rect 25004 2592 25010 2604
rect 25409 2601 25421 2604
rect 25455 2601 25467 2635
rect 25409 2595 25467 2601
rect 29638 2592 29644 2644
rect 29696 2632 29702 2644
rect 29917 2635 29975 2641
rect 29917 2632 29929 2635
rect 29696 2604 29929 2632
rect 29696 2592 29702 2604
rect 29917 2601 29929 2604
rect 29963 2601 29975 2635
rect 29917 2595 29975 2601
rect 48958 2564 48964 2576
rect 44100 2536 48964 2564
rect 1578 2496 1584 2508
rect 1539 2468 1584 2496
rect 1578 2456 1584 2468
rect 1636 2456 1642 2508
rect 2958 2456 2964 2508
rect 3016 2496 3022 2508
rect 3421 2499 3479 2505
rect 3421 2496 3433 2499
rect 3016 2468 3433 2496
rect 3016 2456 3022 2468
rect 3421 2465 3433 2468
rect 3467 2465 3479 2499
rect 4062 2496 4068 2508
rect 4023 2468 4068 2496
rect 3421 2459 3479 2465
rect 4062 2456 4068 2468
rect 4120 2456 4126 2508
rect 4522 2496 4528 2508
rect 4483 2468 4528 2496
rect 4522 2456 4528 2468
rect 4580 2456 4586 2508
rect 6638 2496 6644 2508
rect 6599 2468 6644 2496
rect 6638 2456 6644 2468
rect 6696 2456 6702 2508
rect 6822 2496 6828 2508
rect 6783 2468 6828 2496
rect 6822 2456 6828 2468
rect 6880 2456 6886 2508
rect 7098 2496 7104 2508
rect 7059 2468 7104 2496
rect 7098 2456 7104 2468
rect 7156 2456 7162 2508
rect 11885 2499 11943 2505
rect 11885 2465 11897 2499
rect 11931 2496 11943 2499
rect 12434 2496 12440 2508
rect 11931 2468 12440 2496
rect 11931 2465 11943 2468
rect 11885 2459 11943 2465
rect 12434 2456 12440 2468
rect 12492 2456 12498 2508
rect 12894 2496 12900 2508
rect 12855 2468 12900 2496
rect 12894 2456 12900 2468
rect 12952 2456 12958 2508
rect 19334 2456 19340 2508
rect 19392 2496 19398 2508
rect 19429 2499 19487 2505
rect 19429 2496 19441 2499
rect 19392 2468 19441 2496
rect 19392 2456 19398 2468
rect 19429 2465 19441 2468
rect 19475 2465 19487 2499
rect 19429 2459 19487 2465
rect 19610 2456 19616 2508
rect 19668 2496 19674 2508
rect 44100 2505 44128 2536
rect 48958 2524 48964 2536
rect 49016 2524 49022 2576
rect 19889 2499 19947 2505
rect 19889 2496 19901 2499
rect 19668 2468 19901 2496
rect 19668 2456 19674 2468
rect 19889 2465 19901 2468
rect 19935 2465 19947 2499
rect 19889 2459 19947 2465
rect 44085 2499 44143 2505
rect 44085 2465 44097 2499
rect 44131 2465 44143 2499
rect 44085 2459 44143 2465
rect 44637 2499 44695 2505
rect 44637 2465 44649 2499
rect 44683 2496 44695 2499
rect 44726 2496 44732 2508
rect 44683 2468 44732 2496
rect 44683 2465 44695 2468
rect 44637 2459 44695 2465
rect 44726 2456 44732 2468
rect 44784 2456 44790 2508
rect 46753 2499 46811 2505
rect 46753 2465 46765 2499
rect 46799 2496 46811 2499
rect 47670 2496 47676 2508
rect 46799 2468 47676 2496
rect 46799 2465 46811 2468
rect 46753 2459 46811 2465
rect 47670 2456 47676 2468
rect 47728 2456 47734 2508
rect 14182 2388 14188 2440
rect 14240 2428 14246 2440
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 14240 2400 14289 2428
rect 14240 2388 14246 2400
rect 14277 2397 14289 2400
rect 14323 2397 14335 2431
rect 14277 2391 14335 2397
rect 25501 2431 25559 2437
rect 25501 2397 25513 2431
rect 25547 2428 25559 2431
rect 38378 2428 38384 2440
rect 25547 2400 38384 2428
rect 25547 2397 25559 2400
rect 25501 2391 25559 2397
rect 38378 2388 38384 2400
rect 38436 2388 38442 2440
rect 47213 2431 47271 2437
rect 47213 2397 47225 2431
rect 47259 2428 47271 2431
rect 47765 2431 47823 2437
rect 47765 2428 47777 2431
rect 47259 2400 47777 2428
rect 47259 2397 47271 2400
rect 47213 2391 47271 2397
rect 47765 2397 47777 2400
rect 47811 2397 47823 2431
rect 47765 2391 47823 2397
rect 3237 2363 3295 2369
rect 3237 2329 3249 2363
rect 3283 2329 3295 2363
rect 3237 2323 3295 2329
rect 4249 2363 4307 2369
rect 4249 2329 4261 2363
rect 4295 2360 4307 2363
rect 4614 2360 4620 2372
rect 4295 2332 4620 2360
rect 4295 2329 4307 2332
rect 4249 2323 4307 2329
rect 3252 2292 3280 2323
rect 4614 2320 4620 2332
rect 4672 2320 4678 2372
rect 12069 2363 12127 2369
rect 12069 2329 12081 2363
rect 12115 2360 12127 2363
rect 12526 2360 12532 2372
rect 12115 2332 12532 2360
rect 12115 2329 12127 2332
rect 12069 2323 12127 2329
rect 12526 2320 12532 2332
rect 12584 2320 12590 2372
rect 19613 2363 19671 2369
rect 19613 2329 19625 2363
rect 19659 2360 19671 2363
rect 20162 2360 20168 2372
rect 19659 2332 20168 2360
rect 19659 2329 19671 2332
rect 19613 2323 19671 2329
rect 20162 2320 20168 2332
rect 20220 2320 20226 2372
rect 28994 2320 29000 2372
rect 29052 2360 29058 2372
rect 29825 2363 29883 2369
rect 29825 2360 29837 2363
rect 29052 2332 29837 2360
rect 29052 2320 29058 2332
rect 29825 2329 29837 2332
rect 29871 2329 29883 2363
rect 29825 2323 29883 2329
rect 38654 2320 38660 2372
rect 38712 2360 38718 2372
rect 38933 2363 38991 2369
rect 38933 2360 38945 2363
rect 38712 2332 38945 2360
rect 38712 2320 38718 2332
rect 38933 2329 38945 2332
rect 38979 2329 38991 2363
rect 38933 2323 38991 2329
rect 44453 2363 44511 2369
rect 44453 2329 44465 2363
rect 44499 2360 44511 2363
rect 45554 2360 45560 2372
rect 44499 2332 45560 2360
rect 44499 2329 44511 2332
rect 44453 2323 44511 2329
rect 45554 2320 45560 2332
rect 45612 2320 45618 2372
rect 46934 2320 46940 2372
rect 46992 2360 46998 2372
rect 47029 2363 47087 2369
rect 47029 2360 47041 2363
rect 46992 2332 47041 2360
rect 46992 2320 46998 2332
rect 47029 2329 47041 2332
rect 47075 2329 47087 2363
rect 47029 2323 47087 2329
rect 5350 2292 5356 2304
rect 3252 2264 5356 2292
rect 5350 2252 5356 2264
rect 5408 2252 5414 2304
rect 30650 2252 30656 2304
rect 30708 2292 30714 2304
rect 38841 2295 38899 2301
rect 38841 2292 38853 2295
rect 30708 2264 38853 2292
rect 30708 2252 30714 2264
rect 38841 2261 38853 2264
rect 38887 2261 38899 2295
rect 38841 2255 38899 2261
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
rect 44174 2048 44180 2100
rect 44232 2088 44238 2100
rect 46842 2088 46848 2100
rect 44232 2060 46848 2088
rect 44232 2048 44238 2060
rect 46842 2048 46848 2060
rect 46900 2048 46906 2100
rect 2866 1640 2872 1692
rect 2924 1680 2930 1692
rect 5534 1680 5540 1692
rect 2924 1652 5540 1680
rect 2924 1640 2930 1652
rect 5534 1640 5540 1652
rect 5592 1640 5598 1692
<< via1 >>
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 7196 47200 7248 47252
rect 4804 47132 4856 47184
rect 8300 47132 8352 47184
rect 17408 47132 17460 47184
rect 20444 47132 20496 47184
rect 24676 47132 24728 47184
rect 43628 47132 43680 47184
rect 4988 47064 5040 47116
rect 6000 47064 6052 47116
rect 14188 47064 14240 47116
rect 39764 47064 39816 47116
rect 46756 47107 46808 47116
rect 46756 47073 46765 47107
rect 46765 47073 46799 47107
rect 46799 47073 46808 47107
rect 46756 47064 46808 47073
rect 4528 46996 4580 47048
rect 9036 46996 9088 47048
rect 12440 47039 12492 47048
rect 12440 47005 12449 47039
rect 12449 47005 12483 47039
rect 12483 47005 12492 47039
rect 12440 46996 12492 47005
rect 17500 47039 17552 47048
rect 17500 47005 17509 47039
rect 17509 47005 17543 47039
rect 17543 47005 17552 47039
rect 17500 46996 17552 47005
rect 19340 46996 19392 47048
rect 22468 46996 22520 47048
rect 23848 46996 23900 47048
rect 25320 47039 25372 47048
rect 25320 47005 25329 47039
rect 25329 47005 25363 47039
rect 25363 47005 25372 47039
rect 25320 46996 25372 47005
rect 29736 46996 29788 47048
rect 31760 46996 31812 47048
rect 33140 47039 33192 47048
rect 33140 47005 33149 47039
rect 33149 47005 33183 47039
rect 33183 47005 33192 47039
rect 33140 46996 33192 47005
rect 38936 47039 38988 47048
rect 38936 47005 38945 47039
rect 38945 47005 38979 47039
rect 38979 47005 38988 47039
rect 38936 46996 38988 47005
rect 40132 47039 40184 47048
rect 40132 47005 40141 47039
rect 40141 47005 40175 47039
rect 40175 47005 40184 47039
rect 40132 46996 40184 47005
rect 41512 47039 41564 47048
rect 41512 47005 41521 47039
rect 41521 47005 41555 47039
rect 41555 47005 41564 47039
rect 41512 46996 41564 47005
rect 42524 46996 42576 47048
rect 47216 47039 47268 47048
rect 47216 47005 47225 47039
rect 47225 47005 47259 47039
rect 47259 47005 47268 47039
rect 47216 46996 47268 47005
rect 48964 46996 49016 47048
rect 2320 46971 2372 46980
rect 2320 46937 2329 46971
rect 2329 46937 2363 46971
rect 2363 46937 2372 46971
rect 2320 46928 2372 46937
rect 1308 46860 1360 46912
rect 4712 46928 4764 46980
rect 13820 46928 13872 46980
rect 47032 46971 47084 46980
rect 47032 46937 47041 46971
rect 47041 46937 47075 46971
rect 47075 46937 47084 46971
rect 47032 46928 47084 46937
rect 47768 46928 47820 46980
rect 3516 46860 3568 46912
rect 32496 46903 32548 46912
rect 32496 46869 32505 46903
rect 32505 46869 32539 46903
rect 32539 46869 32548 46903
rect 32496 46860 32548 46869
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 1952 46656 2004 46708
rect 7196 46699 7248 46708
rect 3516 46631 3568 46640
rect 3516 46597 3525 46631
rect 3525 46597 3559 46631
rect 3559 46597 3568 46631
rect 3516 46588 3568 46597
rect 7196 46665 7205 46699
rect 7205 46665 7239 46699
rect 7239 46665 7248 46699
rect 7196 46656 7248 46665
rect 33140 46656 33192 46708
rect 4620 46588 4672 46640
rect 4528 46520 4580 46572
rect 6000 46563 6052 46572
rect 6000 46529 6009 46563
rect 6009 46529 6043 46563
rect 6043 46529 6052 46563
rect 6000 46520 6052 46529
rect 2596 46495 2648 46504
rect 2596 46461 2605 46495
rect 2605 46461 2639 46495
rect 2639 46461 2648 46495
rect 2596 46452 2648 46461
rect 5816 46495 5868 46504
rect 5816 46461 5825 46495
rect 5825 46461 5859 46495
rect 5859 46461 5868 46495
rect 5816 46452 5868 46461
rect 4068 46384 4120 46436
rect 12440 46588 12492 46640
rect 22468 46563 22520 46572
rect 22468 46529 22477 46563
rect 22477 46529 22511 46563
rect 22511 46529 22520 46563
rect 22468 46520 22520 46529
rect 25320 46588 25372 46640
rect 39764 46563 39816 46572
rect 39764 46529 39773 46563
rect 39773 46529 39807 46563
rect 39807 46529 39816 46563
rect 39764 46520 39816 46529
rect 41512 46520 41564 46572
rect 47400 46520 47452 46572
rect 12900 46452 12952 46504
rect 12992 46495 13044 46504
rect 12992 46461 13001 46495
rect 13001 46461 13035 46495
rect 13035 46461 13044 46495
rect 14372 46495 14424 46504
rect 12992 46452 13044 46461
rect 14372 46461 14381 46495
rect 14381 46461 14415 46495
rect 14415 46461 14424 46495
rect 14372 46452 14424 46461
rect 14556 46495 14608 46504
rect 14556 46461 14565 46495
rect 14565 46461 14599 46495
rect 14599 46461 14608 46495
rect 14556 46452 14608 46461
rect 14832 46495 14884 46504
rect 14832 46461 14841 46495
rect 14841 46461 14875 46495
rect 14875 46461 14884 46495
rect 14832 46452 14884 46461
rect 22652 46495 22704 46504
rect 22652 46461 22661 46495
rect 22661 46461 22695 46495
rect 22695 46461 22704 46495
rect 22652 46452 22704 46461
rect 23204 46495 23256 46504
rect 23204 46461 23213 46495
rect 23213 46461 23247 46495
rect 23247 46461 23256 46495
rect 23204 46452 23256 46461
rect 24952 46495 25004 46504
rect 24952 46461 24961 46495
rect 24961 46461 24995 46495
rect 24995 46461 25004 46495
rect 24952 46452 25004 46461
rect 25780 46495 25832 46504
rect 25780 46461 25789 46495
rect 25789 46461 25823 46495
rect 25823 46461 25832 46495
rect 25780 46452 25832 46461
rect 29368 46495 29420 46504
rect 29368 46461 29377 46495
rect 29377 46461 29411 46495
rect 29411 46461 29420 46495
rect 29368 46452 29420 46461
rect 29644 46495 29696 46504
rect 29644 46461 29653 46495
rect 29653 46461 29687 46495
rect 29687 46461 29696 46495
rect 29644 46452 29696 46461
rect 33232 46495 33284 46504
rect 33232 46461 33241 46495
rect 33241 46461 33275 46495
rect 33275 46461 33284 46495
rect 33232 46452 33284 46461
rect 33508 46495 33560 46504
rect 33508 46461 33517 46495
rect 33517 46461 33551 46495
rect 33551 46461 33560 46495
rect 33508 46452 33560 46461
rect 37648 46495 37700 46504
rect 37648 46461 37657 46495
rect 37657 46461 37691 46495
rect 37691 46461 37700 46495
rect 37648 46452 37700 46461
rect 39948 46495 40000 46504
rect 36728 46384 36780 46436
rect 39948 46461 39957 46495
rect 39957 46461 39991 46495
rect 39991 46461 40000 46495
rect 39948 46452 40000 46461
rect 42800 46495 42852 46504
rect 38660 46384 38712 46436
rect 42800 46461 42809 46495
rect 42809 46461 42843 46495
rect 42843 46461 42852 46495
rect 42800 46452 42852 46461
rect 41880 46384 41932 46436
rect 45928 46452 45980 46504
rect 46388 46495 46440 46504
rect 46388 46461 46397 46495
rect 46397 46461 46431 46495
rect 46431 46461 46440 46495
rect 46388 46452 46440 46461
rect 45836 46384 45888 46436
rect 4896 46316 4948 46368
rect 10508 46359 10560 46368
rect 10508 46325 10517 46359
rect 10517 46325 10551 46359
rect 10551 46325 10560 46359
rect 10508 46316 10560 46325
rect 12992 46316 13044 46368
rect 16856 46359 16908 46368
rect 16856 46325 16865 46359
rect 16865 46325 16899 46359
rect 16899 46325 16908 46359
rect 16856 46316 16908 46325
rect 19248 46316 19300 46368
rect 27068 46316 27120 46368
rect 35348 46316 35400 46368
rect 46664 46316 46716 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 5816 46112 5868 46164
rect 12900 46155 12952 46164
rect 12900 46121 12909 46155
rect 12909 46121 12943 46155
rect 12943 46121 12952 46155
rect 12900 46112 12952 46121
rect 13820 46112 13872 46164
rect 14556 46112 14608 46164
rect 22652 46155 22704 46164
rect 22652 46121 22661 46155
rect 22661 46121 22695 46155
rect 22695 46121 22704 46155
rect 22652 46112 22704 46121
rect 29368 46112 29420 46164
rect 33232 46155 33284 46164
rect 33232 46121 33241 46155
rect 33241 46121 33275 46155
rect 33275 46121 33284 46155
rect 33232 46112 33284 46121
rect 39948 46112 40000 46164
rect 45928 46155 45980 46164
rect 45928 46121 45937 46155
rect 45937 46121 45971 46155
rect 45971 46121 45980 46155
rect 45928 46112 45980 46121
rect 5080 46044 5132 46096
rect 2780 46019 2832 46028
rect 2780 45985 2789 46019
rect 2789 45985 2823 46019
rect 2823 45985 2832 46019
rect 2780 45976 2832 45985
rect 4620 45976 4672 46028
rect 10508 46019 10560 46028
rect 10508 45985 10517 46019
rect 10517 45985 10551 46019
rect 10551 45985 10560 46019
rect 10508 45976 10560 45985
rect 10968 45976 11020 46028
rect 15476 46019 15528 46028
rect 15476 45985 15485 46019
rect 15485 45985 15519 46019
rect 15519 45985 15528 46019
rect 15476 45976 15528 45985
rect 16856 46019 16908 46028
rect 16856 45985 16865 46019
rect 16865 45985 16899 46019
rect 16899 45985 16908 46019
rect 16856 45976 16908 45985
rect 25228 46044 25280 46096
rect 25136 46019 25188 46028
rect 4804 45908 4856 45960
rect 6368 45951 6420 45960
rect 6368 45917 6377 45951
rect 6377 45917 6411 45951
rect 6411 45917 6420 45951
rect 7012 45951 7064 45960
rect 6368 45908 6420 45917
rect 5540 45840 5592 45892
rect 7012 45917 7021 45951
rect 7021 45917 7055 45951
rect 7055 45917 7064 45951
rect 7012 45908 7064 45917
rect 13268 45908 13320 45960
rect 10692 45883 10744 45892
rect 6920 45815 6972 45824
rect 6920 45781 6929 45815
rect 6929 45781 6963 45815
rect 6963 45781 6972 45815
rect 6920 45772 6972 45781
rect 10692 45849 10701 45883
rect 10701 45849 10735 45883
rect 10735 45849 10744 45883
rect 10692 45840 10744 45849
rect 16672 45883 16724 45892
rect 16672 45849 16681 45883
rect 16681 45849 16715 45883
rect 16715 45849 16724 45883
rect 16672 45840 16724 45849
rect 25136 45985 25145 46019
rect 25145 45985 25179 46019
rect 25179 45985 25188 46019
rect 25136 45976 25188 45985
rect 29736 46019 29788 46028
rect 29736 45985 29745 46019
rect 29745 45985 29779 46019
rect 29779 45985 29788 46019
rect 29736 45976 29788 45985
rect 30288 45976 30340 46028
rect 35348 46019 35400 46028
rect 35348 45985 35357 46019
rect 35357 45985 35391 46019
rect 35391 45985 35400 46019
rect 35348 45976 35400 45985
rect 36084 46019 36136 46028
rect 36084 45985 36093 46019
rect 36093 45985 36127 46019
rect 36127 45985 36136 46019
rect 36084 45976 36136 45985
rect 24584 45951 24636 45960
rect 24584 45917 24593 45951
rect 24593 45917 24627 45951
rect 24627 45917 24636 45951
rect 24584 45908 24636 45917
rect 29000 45951 29052 45960
rect 29000 45917 29009 45951
rect 29009 45917 29043 45951
rect 29043 45917 29052 45951
rect 29000 45908 29052 45917
rect 33140 45951 33192 45960
rect 33140 45917 33149 45951
rect 33149 45917 33183 45951
rect 33183 45917 33192 45951
rect 33140 45908 33192 45917
rect 38292 45951 38344 45960
rect 38292 45917 38301 45951
rect 38301 45917 38335 45951
rect 38335 45917 38344 45951
rect 38292 45908 38344 45917
rect 38384 45908 38436 45960
rect 29920 45883 29972 45892
rect 29920 45849 29929 45883
rect 29929 45849 29963 45883
rect 29963 45849 29972 45883
rect 29920 45840 29972 45849
rect 35624 45840 35676 45892
rect 22560 45772 22612 45824
rect 25320 45772 25372 45824
rect 39120 45772 39172 45824
rect 40132 46019 40184 46028
rect 40132 45985 40141 46019
rect 40141 45985 40175 46019
rect 40175 45985 40184 46019
rect 40132 45976 40184 45985
rect 40592 46019 40644 46028
rect 40592 45985 40601 46019
rect 40601 45985 40635 46019
rect 40635 45985 40644 46019
rect 40592 45976 40644 45985
rect 46664 46019 46716 46028
rect 46664 45985 46673 46019
rect 46673 45985 46707 46019
rect 46707 45985 46716 46019
rect 46664 45976 46716 45985
rect 48320 46019 48372 46028
rect 48320 45985 48329 46019
rect 48329 45985 48363 46019
rect 48363 45985 48372 46019
rect 48320 45976 48372 45985
rect 46020 45951 46072 45960
rect 46020 45917 46029 45951
rect 46029 45917 46063 45951
rect 46063 45917 46072 45951
rect 46020 45908 46072 45917
rect 40316 45883 40368 45892
rect 40316 45849 40325 45883
rect 40325 45849 40359 45883
rect 40359 45849 40368 45883
rect 40316 45840 40368 45849
rect 47400 45772 47452 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 10692 45568 10744 45620
rect 24952 45568 25004 45620
rect 25320 45568 25372 45620
rect 38384 45568 38436 45620
rect 6920 45500 6972 45552
rect 7012 45500 7064 45552
rect 29920 45543 29972 45552
rect 5540 45432 5592 45484
rect 6736 45475 6788 45484
rect 6736 45441 6745 45475
rect 6745 45441 6779 45475
rect 6779 45441 6788 45475
rect 6736 45432 6788 45441
rect 2872 45407 2924 45416
rect 2872 45373 2881 45407
rect 2881 45373 2915 45407
rect 2915 45373 2924 45407
rect 2872 45364 2924 45373
rect 4896 45364 4948 45416
rect 5356 45364 5408 45416
rect 6368 45364 6420 45416
rect 7380 45407 7432 45416
rect 7380 45373 7389 45407
rect 7389 45373 7423 45407
rect 7423 45373 7432 45407
rect 7380 45364 7432 45373
rect 14372 45432 14424 45484
rect 15108 45475 15160 45484
rect 15108 45441 15117 45475
rect 15117 45441 15151 45475
rect 15151 45441 15160 45475
rect 15108 45432 15160 45441
rect 16672 45432 16724 45484
rect 24584 45432 24636 45484
rect 25228 45432 25280 45484
rect 29920 45509 29929 45543
rect 29929 45509 29963 45543
rect 29963 45509 29972 45543
rect 29920 45500 29972 45509
rect 35624 45543 35676 45552
rect 35624 45509 35633 45543
rect 35633 45509 35667 45543
rect 35667 45509 35676 45543
rect 35624 45500 35676 45509
rect 37648 45500 37700 45552
rect 39120 45543 39172 45552
rect 39120 45509 39129 45543
rect 39129 45509 39163 45543
rect 39163 45509 39172 45543
rect 39120 45500 39172 45509
rect 42800 45500 42852 45552
rect 29828 45475 29880 45484
rect 29828 45441 29837 45475
rect 29837 45441 29871 45475
rect 29871 45441 29880 45475
rect 29828 45432 29880 45441
rect 12532 45364 12584 45416
rect 22560 45364 22612 45416
rect 29000 45296 29052 45348
rect 37280 45432 37332 45484
rect 38292 45432 38344 45484
rect 38936 45475 38988 45484
rect 38936 45441 38945 45475
rect 38945 45441 38979 45475
rect 38979 45441 38988 45475
rect 38936 45432 38988 45441
rect 40132 45364 40184 45416
rect 46940 45500 46992 45552
rect 47032 45500 47084 45552
rect 45836 45432 45888 45484
rect 47400 45432 47452 45484
rect 46296 45364 46348 45416
rect 5448 45228 5500 45280
rect 6736 45228 6788 45280
rect 12532 45228 12584 45280
rect 25228 45228 25280 45280
rect 35716 45228 35768 45280
rect 48320 45228 48372 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 4988 45024 5040 45076
rect 5448 45024 5500 45076
rect 15108 45024 15160 45076
rect 40132 45024 40184 45076
rect 40316 45024 40368 45076
rect 7380 44956 7432 45008
rect 6828 44931 6880 44940
rect 6828 44897 6837 44931
rect 6837 44897 6871 44931
rect 6871 44897 6880 44931
rect 6828 44888 6880 44897
rect 2044 44820 2096 44872
rect 2320 44820 2372 44872
rect 5540 44820 5592 44872
rect 46848 44931 46900 44940
rect 46848 44897 46857 44931
rect 46857 44897 46891 44931
rect 46891 44897 46900 44931
rect 46848 44888 46900 44897
rect 48320 44931 48372 44940
rect 48320 44897 48329 44931
rect 48329 44897 48363 44931
rect 48363 44897 48372 44931
rect 48320 44888 48372 44897
rect 46020 44820 46072 44872
rect 46388 44820 46440 44872
rect 3240 44795 3292 44804
rect 3240 44761 3249 44795
rect 3249 44761 3283 44795
rect 3283 44761 3292 44795
rect 3240 44752 3292 44761
rect 47860 44752 47912 44804
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 4620 44480 4672 44532
rect 3240 44412 3292 44464
rect 5540 44412 5592 44464
rect 6828 44480 6880 44532
rect 15108 44480 15160 44532
rect 47860 44523 47912 44532
rect 47860 44489 47869 44523
rect 47869 44489 47903 44523
rect 47903 44489 47912 44523
rect 47860 44480 47912 44489
rect 13268 44412 13320 44464
rect 46940 44412 46992 44464
rect 2044 44387 2096 44396
rect 2044 44353 2053 44387
rect 2053 44353 2087 44387
rect 2087 44353 2096 44387
rect 2044 44344 2096 44353
rect 4988 44387 5040 44396
rect 3056 44276 3108 44328
rect 3148 44319 3200 44328
rect 3148 44285 3157 44319
rect 3157 44285 3191 44319
rect 3191 44285 3200 44319
rect 4988 44353 4997 44387
rect 4997 44353 5031 44387
rect 5031 44353 5040 44387
rect 4988 44344 5040 44353
rect 5172 44344 5224 44396
rect 37280 44344 37332 44396
rect 47216 44387 47268 44396
rect 47216 44353 47225 44387
rect 47225 44353 47259 44387
rect 47259 44353 47268 44387
rect 47216 44344 47268 44353
rect 5816 44319 5868 44328
rect 3148 44276 3200 44285
rect 5816 44285 5825 44319
rect 5825 44285 5859 44319
rect 5859 44285 5868 44319
rect 5816 44276 5868 44285
rect 33140 44276 33192 44328
rect 4620 44208 4672 44260
rect 5080 44208 5132 44260
rect 7288 44140 7340 44192
rect 29000 44140 29052 44192
rect 29644 44140 29696 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 3516 43800 3568 43852
rect 5264 43800 5316 43852
rect 5724 43843 5776 43852
rect 5724 43809 5733 43843
rect 5733 43809 5767 43843
rect 5767 43809 5776 43843
rect 5724 43800 5776 43809
rect 7288 43843 7340 43852
rect 7288 43809 7297 43843
rect 7297 43809 7331 43843
rect 7331 43809 7340 43843
rect 7288 43800 7340 43809
rect 2044 43732 2096 43784
rect 4988 43775 5040 43784
rect 4988 43741 4997 43775
rect 4997 43741 5031 43775
rect 5031 43741 5040 43775
rect 4988 43732 5040 43741
rect 5908 43664 5960 43716
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 5908 43435 5960 43444
rect 5908 43401 5917 43435
rect 5917 43401 5951 43435
rect 5951 43401 5960 43435
rect 5908 43392 5960 43401
rect 5172 43367 5224 43376
rect 5172 43333 5181 43367
rect 5181 43333 5215 43367
rect 5215 43333 5224 43367
rect 5172 43324 5224 43333
rect 2044 43299 2096 43308
rect 2044 43265 2053 43299
rect 2053 43265 2087 43299
rect 2087 43265 2096 43299
rect 2044 43256 2096 43265
rect 3516 43256 3568 43308
rect 6736 43324 6788 43376
rect 6000 43299 6052 43308
rect 6000 43265 6009 43299
rect 6009 43265 6043 43299
rect 6043 43265 6052 43299
rect 6000 43256 6052 43265
rect 29828 43256 29880 43308
rect 47676 43256 47728 43308
rect 2228 43231 2280 43240
rect 2228 43197 2237 43231
rect 2237 43197 2271 43231
rect 2271 43197 2280 43231
rect 2228 43188 2280 43197
rect 2780 43231 2832 43240
rect 2780 43197 2789 43231
rect 2789 43197 2823 43231
rect 2823 43197 2832 43231
rect 2780 43188 2832 43197
rect 47032 43095 47084 43104
rect 47032 43061 47041 43095
rect 47041 43061 47075 43095
rect 47075 43061 47084 43095
rect 47032 43052 47084 43061
rect 47860 43095 47912 43104
rect 47860 43061 47869 43095
rect 47869 43061 47903 43095
rect 47903 43061 47912 43095
rect 47860 43052 47912 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 2228 42848 2280 42900
rect 2504 42687 2556 42696
rect 2504 42653 2513 42687
rect 2513 42653 2547 42687
rect 2547 42653 2556 42687
rect 3516 42780 3568 42832
rect 3056 42755 3108 42764
rect 3056 42721 3065 42755
rect 3065 42721 3099 42755
rect 3099 42721 3108 42755
rect 3056 42712 3108 42721
rect 5264 42712 5316 42764
rect 47032 42712 47084 42764
rect 48228 42755 48280 42764
rect 48228 42721 48237 42755
rect 48237 42721 48271 42755
rect 48271 42721 48280 42755
rect 48228 42712 48280 42721
rect 2504 42644 2556 42653
rect 4988 42644 5040 42696
rect 5632 42576 5684 42628
rect 6000 42576 6052 42628
rect 13084 42576 13136 42628
rect 47860 42576 47912 42628
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 7288 41964 7340 42016
rect 46480 41964 46532 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 7288 41667 7340 41676
rect 7288 41633 7297 41667
rect 7297 41633 7331 41667
rect 7331 41633 7340 41667
rect 7288 41624 7340 41633
rect 46480 41667 46532 41676
rect 46480 41633 46489 41667
rect 46489 41633 46523 41667
rect 46523 41633 46532 41667
rect 46480 41624 46532 41633
rect 48228 41667 48280 41676
rect 48228 41633 48237 41667
rect 48237 41633 48271 41667
rect 48271 41633 48280 41667
rect 48228 41624 48280 41633
rect 3056 41488 3108 41540
rect 7104 41531 7156 41540
rect 7104 41497 7113 41531
rect 7113 41497 7147 41531
rect 7147 41497 7156 41531
rect 7104 41488 7156 41497
rect 47124 41488 47176 41540
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 7104 41216 7156 41268
rect 47124 41259 47176 41268
rect 47124 41225 47133 41259
rect 47133 41225 47167 41259
rect 47167 41225 47176 41259
rect 47124 41216 47176 41225
rect 6092 41080 6144 41132
rect 7380 41080 7432 41132
rect 46940 41080 46992 41132
rect 46480 40876 46532 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 46480 40579 46532 40588
rect 46480 40545 46489 40579
rect 46489 40545 46523 40579
rect 46523 40545 46532 40579
rect 46480 40536 46532 40545
rect 14740 40468 14792 40520
rect 19064 40468 19116 40520
rect 23664 40511 23716 40520
rect 23664 40477 23673 40511
rect 23673 40477 23707 40511
rect 23707 40477 23716 40511
rect 23664 40468 23716 40477
rect 23848 40511 23900 40520
rect 23848 40477 23857 40511
rect 23857 40477 23891 40511
rect 23891 40477 23900 40511
rect 23848 40468 23900 40477
rect 16028 40443 16080 40452
rect 16028 40409 16037 40443
rect 16037 40409 16071 40443
rect 16071 40409 16080 40443
rect 16028 40400 16080 40409
rect 45560 40400 45612 40452
rect 47124 40400 47176 40452
rect 48320 40443 48372 40452
rect 48320 40409 48329 40443
rect 48329 40409 48363 40443
rect 48363 40409 48372 40443
rect 48320 40400 48372 40409
rect 17776 40332 17828 40384
rect 22284 40332 22336 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 16028 40171 16080 40180
rect 16028 40137 16037 40171
rect 16037 40137 16071 40171
rect 16071 40137 16080 40171
rect 16028 40128 16080 40137
rect 24400 40128 24452 40180
rect 3240 40060 3292 40112
rect 8208 40060 8260 40112
rect 12992 40103 13044 40112
rect 12992 40069 13001 40103
rect 13001 40069 13035 40103
rect 13035 40069 13044 40103
rect 12992 40060 13044 40069
rect 17776 40103 17828 40112
rect 17776 40069 17785 40103
rect 17785 40069 17819 40103
rect 17819 40069 17828 40103
rect 17776 40060 17828 40069
rect 22192 40060 22244 40112
rect 14648 39967 14700 39976
rect 14648 39933 14657 39967
rect 14657 39933 14691 39967
rect 14691 39933 14700 39967
rect 14648 39924 14700 39933
rect 14924 39924 14976 39976
rect 13084 39856 13136 39908
rect 21732 39992 21784 40044
rect 24032 40060 24084 40112
rect 16948 39924 17000 39976
rect 19248 39967 19300 39976
rect 19248 39933 19257 39967
rect 19257 39933 19291 39967
rect 19291 39933 19300 39967
rect 19248 39924 19300 39933
rect 22284 39924 22336 39976
rect 19064 39856 19116 39908
rect 20904 39856 20956 39908
rect 24952 39992 25004 40044
rect 47124 40035 47176 40044
rect 47124 40001 47133 40035
rect 47133 40001 47167 40035
rect 47167 40001 47176 40035
rect 47124 39992 47176 40001
rect 23940 39967 23992 39976
rect 23940 39933 23949 39967
rect 23949 39933 23983 39967
rect 23983 39933 23992 39967
rect 23940 39924 23992 39933
rect 24492 39967 24544 39976
rect 24492 39933 24501 39967
rect 24501 39933 24535 39967
rect 24535 39933 24544 39967
rect 24492 39924 24544 39933
rect 46388 39924 46440 39976
rect 47400 39992 47452 40044
rect 23020 39856 23072 39908
rect 23664 39788 23716 39840
rect 48320 39788 48372 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 14648 39584 14700 39636
rect 23848 39584 23900 39636
rect 23756 39516 23808 39568
rect 16028 39448 16080 39500
rect 23020 39448 23072 39500
rect 46848 39491 46900 39500
rect 46848 39457 46857 39491
rect 46857 39457 46891 39491
rect 46891 39457 46900 39491
rect 46848 39448 46900 39457
rect 48320 39491 48372 39500
rect 48320 39457 48329 39491
rect 48329 39457 48363 39491
rect 48363 39457 48372 39491
rect 48320 39448 48372 39457
rect 13084 39423 13136 39432
rect 13084 39389 13093 39423
rect 13093 39389 13127 39423
rect 13127 39389 13136 39423
rect 13084 39380 13136 39389
rect 21732 39423 21784 39432
rect 21732 39389 21741 39423
rect 21741 39389 21775 39423
rect 21775 39389 21784 39423
rect 21732 39380 21784 39389
rect 22376 39423 22428 39432
rect 22376 39389 22385 39423
rect 22385 39389 22419 39423
rect 22419 39389 22428 39423
rect 22376 39380 22428 39389
rect 23664 39423 23716 39432
rect 22192 39312 22244 39364
rect 23664 39389 23673 39423
rect 23673 39389 23707 39423
rect 23707 39389 23716 39423
rect 23664 39380 23716 39389
rect 23756 39423 23808 39432
rect 23756 39389 23765 39423
rect 23765 39389 23799 39423
rect 23799 39389 23808 39423
rect 23756 39380 23808 39389
rect 24032 39380 24084 39432
rect 24492 39380 24544 39432
rect 25596 39423 25648 39432
rect 25596 39389 25605 39423
rect 25605 39389 25639 39423
rect 25639 39389 25648 39423
rect 25596 39380 25648 39389
rect 24952 39355 25004 39364
rect 24952 39321 24961 39355
rect 24961 39321 24995 39355
rect 24995 39321 25004 39355
rect 24952 39312 25004 39321
rect 47860 39312 47912 39364
rect 23572 39244 23624 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 47860 39083 47912 39092
rect 47860 39049 47869 39083
rect 47869 39049 47903 39083
rect 47903 39049 47912 39083
rect 47860 39040 47912 39049
rect 20904 39015 20956 39024
rect 20904 38981 20913 39015
rect 20913 38981 20947 39015
rect 20947 38981 20956 39015
rect 20904 38972 20956 38981
rect 23756 38972 23808 39024
rect 25596 38972 25648 39024
rect 1676 38947 1728 38956
rect 1676 38913 1685 38947
rect 1685 38913 1719 38947
rect 1719 38913 1728 38947
rect 1676 38904 1728 38913
rect 14740 38947 14792 38956
rect 14740 38913 14749 38947
rect 14749 38913 14783 38947
rect 14783 38913 14792 38947
rect 14740 38904 14792 38913
rect 14924 38947 14976 38956
rect 14924 38913 14933 38947
rect 14933 38913 14967 38947
rect 14967 38913 14976 38947
rect 14924 38904 14976 38913
rect 16028 38947 16080 38956
rect 14832 38836 14884 38888
rect 16028 38913 16037 38947
rect 16037 38913 16071 38947
rect 16071 38913 16080 38947
rect 16028 38904 16080 38913
rect 16948 38904 17000 38956
rect 1860 38811 1912 38820
rect 1860 38777 1869 38811
rect 1869 38777 1903 38811
rect 1903 38777 1912 38811
rect 1860 38768 1912 38777
rect 15016 38700 15068 38752
rect 18052 38836 18104 38888
rect 18880 38904 18932 38956
rect 20628 38879 20680 38888
rect 20628 38845 20637 38879
rect 20637 38845 20671 38879
rect 20671 38845 20680 38879
rect 20628 38836 20680 38845
rect 21732 38836 21784 38888
rect 22192 38904 22244 38956
rect 22284 38947 22336 38956
rect 22284 38913 22293 38947
rect 22293 38913 22327 38947
rect 22327 38913 22336 38947
rect 23572 38947 23624 38956
rect 22284 38904 22336 38913
rect 23572 38913 23581 38947
rect 23581 38913 23615 38947
rect 23615 38913 23624 38947
rect 23572 38904 23624 38913
rect 24400 38947 24452 38956
rect 24400 38913 24409 38947
rect 24409 38913 24443 38947
rect 24443 38913 24452 38947
rect 24400 38904 24452 38913
rect 23480 38879 23532 38888
rect 23480 38845 23489 38879
rect 23489 38845 23523 38879
rect 23523 38845 23532 38879
rect 23480 38836 23532 38845
rect 19248 38768 19300 38820
rect 23572 38768 23624 38820
rect 23756 38768 23808 38820
rect 23940 38879 23992 38888
rect 23940 38845 23949 38879
rect 23949 38845 23983 38879
rect 23983 38845 23992 38879
rect 23940 38836 23992 38845
rect 24492 38836 24544 38888
rect 28448 38904 28500 38956
rect 35716 38904 35768 38956
rect 47584 38904 47636 38956
rect 15936 38700 15988 38752
rect 17960 38743 18012 38752
rect 17960 38709 17969 38743
rect 17969 38709 18003 38743
rect 18003 38709 18012 38743
rect 17960 38700 18012 38709
rect 23388 38700 23440 38752
rect 23940 38700 23992 38752
rect 24860 38700 24912 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 14280 38496 14332 38548
rect 14924 38496 14976 38548
rect 16948 38539 17000 38548
rect 16948 38505 16957 38539
rect 16957 38505 16991 38539
rect 16991 38505 17000 38539
rect 16948 38496 17000 38505
rect 18880 38539 18932 38548
rect 18880 38505 18889 38539
rect 18889 38505 18923 38539
rect 18923 38505 18932 38539
rect 18880 38496 18932 38505
rect 22376 38496 22428 38548
rect 23480 38496 23532 38548
rect 25596 38496 25648 38548
rect 15108 38471 15160 38480
rect 15108 38437 15117 38471
rect 15117 38437 15151 38471
rect 15151 38437 15160 38471
rect 15108 38428 15160 38437
rect 4804 38292 4856 38344
rect 8484 38292 8536 38344
rect 12900 38292 12952 38344
rect 15016 38292 15068 38344
rect 15660 38292 15712 38344
rect 22284 38292 22336 38344
rect 23572 38335 23624 38344
rect 23572 38301 23581 38335
rect 23581 38301 23615 38335
rect 23615 38301 23624 38335
rect 23572 38292 23624 38301
rect 24584 38335 24636 38344
rect 24584 38301 24593 38335
rect 24593 38301 24627 38335
rect 24627 38301 24636 38335
rect 24584 38292 24636 38301
rect 24860 38335 24912 38344
rect 24860 38301 24894 38335
rect 24894 38301 24912 38335
rect 24860 38292 24912 38301
rect 48320 38292 48372 38344
rect 12808 38224 12860 38276
rect 15844 38267 15896 38276
rect 15844 38233 15878 38267
rect 15878 38233 15896 38267
rect 6552 38199 6604 38208
rect 6552 38165 6561 38199
rect 6561 38165 6595 38199
rect 6595 38165 6604 38199
rect 6552 38156 6604 38165
rect 14832 38156 14884 38208
rect 15844 38224 15896 38233
rect 18696 38224 18748 38276
rect 23664 38224 23716 38276
rect 16948 38156 17000 38208
rect 23848 38156 23900 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 12808 37952 12860 38004
rect 4804 37859 4856 37868
rect 4804 37825 4813 37859
rect 4813 37825 4847 37859
rect 4847 37825 4856 37859
rect 4804 37816 4856 37825
rect 5816 37859 5868 37868
rect 5816 37825 5825 37859
rect 5825 37825 5859 37859
rect 5859 37825 5868 37859
rect 5816 37816 5868 37825
rect 6552 37859 6604 37868
rect 6552 37825 6561 37859
rect 6561 37825 6595 37859
rect 6595 37825 6604 37859
rect 6552 37816 6604 37825
rect 8116 37816 8168 37868
rect 8484 37859 8536 37868
rect 8484 37825 8493 37859
rect 8493 37825 8527 37859
rect 8527 37825 8536 37859
rect 8484 37816 8536 37825
rect 14740 37884 14792 37936
rect 15844 37952 15896 38004
rect 18696 37995 18748 38004
rect 18696 37961 18705 37995
rect 18705 37961 18739 37995
rect 18739 37961 18748 37995
rect 18696 37952 18748 37961
rect 24492 37995 24544 38004
rect 24492 37961 24501 37995
rect 24501 37961 24535 37995
rect 24535 37961 24544 37995
rect 24492 37952 24544 37961
rect 14832 37816 14884 37868
rect 16948 37884 17000 37936
rect 18880 37884 18932 37936
rect 18972 37884 19024 37936
rect 15108 37816 15160 37868
rect 15936 37859 15988 37868
rect 15936 37825 15945 37859
rect 15945 37825 15979 37859
rect 15979 37825 15988 37859
rect 15936 37816 15988 37825
rect 13820 37748 13872 37800
rect 14280 37791 14332 37800
rect 14280 37757 14289 37791
rect 14289 37757 14323 37791
rect 14323 37757 14332 37791
rect 14280 37748 14332 37757
rect 17960 37816 18012 37868
rect 18236 37816 18288 37868
rect 18604 37748 18656 37800
rect 18144 37680 18196 37732
rect 19248 37816 19300 37868
rect 24584 37884 24636 37936
rect 23388 37859 23440 37868
rect 23388 37825 23422 37859
rect 23422 37825 23440 37859
rect 23388 37816 23440 37825
rect 46940 37816 46992 37868
rect 48044 37816 48096 37868
rect 20628 37748 20680 37800
rect 20720 37680 20772 37732
rect 4804 37655 4856 37664
rect 4804 37621 4813 37655
rect 4813 37621 4847 37655
rect 4847 37621 4856 37655
rect 4804 37612 4856 37621
rect 7932 37655 7984 37664
rect 7932 37621 7941 37655
rect 7941 37621 7975 37655
rect 7975 37621 7984 37655
rect 7932 37612 7984 37621
rect 8484 37655 8536 37664
rect 8484 37621 8493 37655
rect 8493 37621 8527 37655
rect 8527 37621 8536 37655
rect 8484 37612 8536 37621
rect 15108 37612 15160 37664
rect 19432 37612 19484 37664
rect 19800 37612 19852 37664
rect 22284 37612 22336 37664
rect 48136 37612 48188 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 7932 37451 7984 37460
rect 7932 37417 7941 37451
rect 7941 37417 7975 37451
rect 7975 37417 7984 37451
rect 7932 37408 7984 37417
rect 18236 37451 18288 37460
rect 18236 37417 18245 37451
rect 18245 37417 18279 37451
rect 18279 37417 18288 37451
rect 18236 37408 18288 37417
rect 20628 37451 20680 37460
rect 20628 37417 20637 37451
rect 20637 37417 20671 37451
rect 20671 37417 20680 37451
rect 20628 37408 20680 37417
rect 5816 37340 5868 37392
rect 16948 37340 17000 37392
rect 2688 37272 2740 37324
rect 4804 37315 4856 37324
rect 4804 37281 4813 37315
rect 4813 37281 4847 37315
rect 4847 37281 4856 37315
rect 4804 37272 4856 37281
rect 13820 37272 13872 37324
rect 14556 37272 14608 37324
rect 17960 37272 18012 37324
rect 18972 37272 19024 37324
rect 4896 37204 4948 37256
rect 7104 37247 7156 37256
rect 7104 37213 7113 37247
rect 7113 37213 7147 37247
rect 7147 37213 7156 37247
rect 7104 37204 7156 37213
rect 1676 37179 1728 37188
rect 1676 37145 1685 37179
rect 1685 37145 1719 37179
rect 1719 37145 1728 37179
rect 1676 37136 1728 37145
rect 14740 37204 14792 37256
rect 14924 37247 14976 37256
rect 14924 37213 14933 37247
rect 14933 37213 14967 37247
rect 14967 37213 14976 37247
rect 14924 37204 14976 37213
rect 15016 37204 15068 37256
rect 18604 37247 18656 37256
rect 15108 37136 15160 37188
rect 17040 37136 17092 37188
rect 18604 37213 18613 37247
rect 18613 37213 18647 37247
rect 18647 37213 18656 37247
rect 18604 37204 18656 37213
rect 19340 37204 19392 37256
rect 19800 37247 19852 37256
rect 19800 37213 19809 37247
rect 19809 37213 19843 37247
rect 19843 37213 19852 37247
rect 19800 37204 19852 37213
rect 20812 37204 20864 37256
rect 23848 37204 23900 37256
rect 24584 37204 24636 37256
rect 27712 37204 27764 37256
rect 9128 37111 9180 37120
rect 9128 37077 9137 37111
rect 9137 37077 9171 37111
rect 9171 37077 9180 37111
rect 9128 37068 9180 37077
rect 13176 37068 13228 37120
rect 14924 37068 14976 37120
rect 18604 37068 18656 37120
rect 20904 37136 20956 37188
rect 22468 37136 22520 37188
rect 23940 37136 23992 37188
rect 28448 37315 28500 37324
rect 28448 37281 28457 37315
rect 28457 37281 28491 37315
rect 28491 37281 28500 37315
rect 28448 37272 28500 37281
rect 48136 37315 48188 37324
rect 48136 37281 48145 37315
rect 48145 37281 48179 37315
rect 48179 37281 48188 37315
rect 48136 37272 48188 37281
rect 28080 37247 28132 37256
rect 28080 37213 28089 37247
rect 28089 37213 28123 37247
rect 28123 37213 28132 37247
rect 28080 37204 28132 37213
rect 28172 37247 28224 37256
rect 28172 37213 28181 37247
rect 28181 37213 28215 37247
rect 28215 37213 28224 37247
rect 46480 37247 46532 37256
rect 28172 37204 28224 37213
rect 46480 37213 46489 37247
rect 46489 37213 46523 37247
rect 46523 37213 46532 37247
rect 46480 37204 46532 37213
rect 48320 37247 48372 37256
rect 48320 37213 48329 37247
rect 48329 37213 48363 37247
rect 48363 37213 48372 37247
rect 48320 37204 48372 37213
rect 24768 37068 24820 37120
rect 26056 37111 26108 37120
rect 26056 37077 26065 37111
rect 26065 37077 26099 37111
rect 26099 37077 26108 37111
rect 26056 37068 26108 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 13820 36864 13872 36916
rect 20904 36907 20956 36916
rect 20904 36873 20913 36907
rect 20913 36873 20947 36907
rect 20947 36873 20956 36907
rect 20904 36864 20956 36873
rect 22192 36864 22244 36916
rect 28172 36864 28224 36916
rect 9128 36796 9180 36848
rect 13176 36839 13228 36848
rect 13176 36805 13210 36839
rect 13210 36805 13228 36839
rect 13176 36796 13228 36805
rect 14740 36796 14792 36848
rect 20628 36839 20680 36848
rect 20628 36805 20637 36839
rect 20637 36805 20671 36839
rect 20671 36805 20680 36839
rect 20628 36796 20680 36805
rect 21732 36796 21784 36848
rect 6000 36728 6052 36780
rect 8484 36728 8536 36780
rect 12900 36771 12952 36780
rect 12900 36737 12909 36771
rect 12909 36737 12943 36771
rect 12943 36737 12952 36771
rect 12900 36728 12952 36737
rect 14924 36728 14976 36780
rect 18236 36728 18288 36780
rect 19340 36728 19392 36780
rect 19524 36771 19576 36780
rect 19524 36737 19533 36771
rect 19533 36737 19567 36771
rect 19567 36737 19576 36771
rect 19524 36728 19576 36737
rect 4068 36660 4120 36712
rect 16488 36660 16540 36712
rect 19432 36703 19484 36712
rect 19432 36669 19441 36703
rect 19441 36669 19475 36703
rect 19475 36669 19484 36703
rect 19432 36660 19484 36669
rect 20720 36771 20772 36780
rect 14740 36592 14792 36644
rect 17316 36592 17368 36644
rect 20352 36592 20404 36644
rect 20720 36737 20729 36771
rect 20729 36737 20763 36771
rect 20763 36737 20772 36771
rect 20720 36728 20772 36737
rect 21548 36728 21600 36780
rect 22284 36771 22336 36780
rect 22284 36737 22293 36771
rect 22293 36737 22327 36771
rect 22327 36737 22336 36771
rect 22284 36728 22336 36737
rect 24952 36771 25004 36780
rect 22468 36660 22520 36712
rect 24952 36737 24961 36771
rect 24961 36737 24995 36771
rect 24995 36737 25004 36771
rect 24952 36728 25004 36737
rect 25596 36771 25648 36780
rect 24860 36660 24912 36712
rect 25596 36737 25605 36771
rect 25605 36737 25639 36771
rect 25639 36737 25648 36771
rect 25596 36728 25648 36737
rect 27712 36771 27764 36780
rect 27712 36737 27721 36771
rect 27721 36737 27755 36771
rect 27755 36737 27764 36771
rect 27712 36728 27764 36737
rect 27988 36771 28040 36780
rect 27988 36737 28022 36771
rect 28022 36737 28040 36771
rect 27988 36728 28040 36737
rect 25688 36592 25740 36644
rect 5448 36524 5500 36576
rect 9220 36567 9272 36576
rect 9220 36533 9229 36567
rect 9229 36533 9263 36567
rect 9263 36533 9272 36567
rect 9220 36524 9272 36533
rect 23940 36524 23992 36576
rect 24768 36524 24820 36576
rect 27712 36524 27764 36576
rect 48320 36524 48372 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 4068 36320 4120 36372
rect 4896 36320 4948 36372
rect 5448 36363 5500 36372
rect 5448 36329 5457 36363
rect 5457 36329 5491 36363
rect 5491 36329 5500 36363
rect 5448 36320 5500 36329
rect 6000 36363 6052 36372
rect 6000 36329 6009 36363
rect 6009 36329 6043 36363
rect 6043 36329 6052 36363
rect 6000 36320 6052 36329
rect 9220 36363 9272 36372
rect 9220 36329 9229 36363
rect 9229 36329 9263 36363
rect 9263 36329 9272 36363
rect 9220 36320 9272 36329
rect 17316 36363 17368 36372
rect 17316 36329 17325 36363
rect 17325 36329 17359 36363
rect 17359 36329 17368 36363
rect 17316 36320 17368 36329
rect 19524 36320 19576 36372
rect 24860 36320 24912 36372
rect 26332 36320 26384 36372
rect 27988 36363 28040 36372
rect 27988 36329 27997 36363
rect 27997 36329 28031 36363
rect 28031 36329 28040 36363
rect 27988 36320 28040 36329
rect 4896 36184 4948 36236
rect 5356 36184 5408 36236
rect 21732 36227 21784 36236
rect 4988 36116 5040 36168
rect 6184 36159 6236 36168
rect 6184 36125 6193 36159
rect 6193 36125 6227 36159
rect 6227 36125 6236 36159
rect 6184 36116 6236 36125
rect 8116 36159 8168 36168
rect 8116 36125 8125 36159
rect 8125 36125 8159 36159
rect 8159 36125 8168 36159
rect 8116 36116 8168 36125
rect 7104 36048 7156 36100
rect 9220 36116 9272 36168
rect 21732 36193 21741 36227
rect 21741 36193 21775 36227
rect 21775 36193 21784 36227
rect 21732 36184 21784 36193
rect 17040 36159 17092 36168
rect 17040 36125 17049 36159
rect 17049 36125 17083 36159
rect 17083 36125 17092 36159
rect 17040 36116 17092 36125
rect 21548 36159 21600 36168
rect 21548 36125 21557 36159
rect 21557 36125 21591 36159
rect 21591 36125 21600 36159
rect 21548 36116 21600 36125
rect 23480 36116 23532 36168
rect 28080 36252 28132 36304
rect 46848 36227 46900 36236
rect 46848 36193 46857 36227
rect 46857 36193 46891 36227
rect 46891 36193 46900 36227
rect 46848 36184 46900 36193
rect 48320 36227 48372 36236
rect 48320 36193 48329 36227
rect 48329 36193 48363 36227
rect 48363 36193 48372 36227
rect 48320 36184 48372 36193
rect 9588 36048 9640 36100
rect 27436 36159 27488 36168
rect 27436 36125 27445 36159
rect 27445 36125 27479 36159
rect 27479 36125 27488 36159
rect 27436 36116 27488 36125
rect 27712 36159 27764 36168
rect 27712 36125 27721 36159
rect 27721 36125 27755 36159
rect 27755 36125 27764 36159
rect 27712 36116 27764 36125
rect 28448 36116 28500 36168
rect 10048 36023 10100 36032
rect 10048 35989 10057 36023
rect 10057 35989 10091 36023
rect 10091 35989 10100 36023
rect 10048 35980 10100 35989
rect 25228 36048 25280 36100
rect 26148 36048 26200 36100
rect 48136 36091 48188 36100
rect 25044 35980 25096 36032
rect 26056 35980 26108 36032
rect 26516 36023 26568 36032
rect 26516 35989 26541 36023
rect 26541 35989 26568 36023
rect 48136 36057 48145 36091
rect 48145 36057 48179 36091
rect 48179 36057 48188 36091
rect 48136 36048 48188 36057
rect 26516 35980 26568 35989
rect 27804 35980 27856 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 6184 35776 6236 35828
rect 14096 35819 14148 35828
rect 14096 35785 14105 35819
rect 14105 35785 14139 35819
rect 14139 35785 14148 35819
rect 14096 35776 14148 35785
rect 21732 35776 21784 35828
rect 24032 35776 24084 35828
rect 24768 35776 24820 35828
rect 24860 35776 24912 35828
rect 25228 35776 25280 35828
rect 28724 35776 28776 35828
rect 48136 35776 48188 35828
rect 10048 35708 10100 35760
rect 5172 35683 5224 35692
rect 5172 35649 5181 35683
rect 5181 35649 5215 35683
rect 5215 35649 5224 35683
rect 5172 35640 5224 35649
rect 9588 35683 9640 35692
rect 9588 35649 9597 35683
rect 9597 35649 9631 35683
rect 9631 35649 9640 35683
rect 9588 35640 9640 35649
rect 15936 35708 15988 35760
rect 14556 35683 14608 35692
rect 14556 35649 14565 35683
rect 14565 35649 14599 35683
rect 14599 35649 14608 35683
rect 14556 35640 14608 35649
rect 19248 35640 19300 35692
rect 22008 35640 22060 35692
rect 25780 35708 25832 35760
rect 23480 35640 23532 35692
rect 24952 35640 25004 35692
rect 25596 35640 25648 35692
rect 26148 35683 26200 35692
rect 26148 35649 26157 35683
rect 26157 35649 26191 35683
rect 26191 35649 26200 35683
rect 26148 35640 26200 35649
rect 26332 35683 26384 35692
rect 26332 35649 26341 35683
rect 26341 35649 26375 35683
rect 26375 35649 26384 35683
rect 26332 35640 26384 35649
rect 26516 35708 26568 35760
rect 27344 35640 27396 35692
rect 32404 35640 32456 35692
rect 33048 35640 33100 35692
rect 34796 35640 34848 35692
rect 17960 35572 18012 35624
rect 23204 35615 23256 35624
rect 23204 35581 23213 35615
rect 23213 35581 23247 35615
rect 23247 35581 23256 35615
rect 23204 35572 23256 35581
rect 17684 35504 17736 35556
rect 24124 35572 24176 35624
rect 27068 35572 27120 35624
rect 34704 35572 34756 35624
rect 47124 35640 47176 35692
rect 24768 35504 24820 35556
rect 24952 35504 25004 35556
rect 26056 35504 26108 35556
rect 5448 35479 5500 35488
rect 5448 35445 5457 35479
rect 5457 35445 5491 35479
rect 5491 35445 5500 35479
rect 5448 35436 5500 35445
rect 8116 35436 8168 35488
rect 14004 35436 14056 35488
rect 14464 35479 14516 35488
rect 14464 35445 14473 35479
rect 14473 35445 14507 35479
rect 14507 35445 14516 35479
rect 14464 35436 14516 35445
rect 18052 35436 18104 35488
rect 21456 35436 21508 35488
rect 23756 35436 23808 35488
rect 25136 35436 25188 35488
rect 27712 35436 27764 35488
rect 28632 35436 28684 35488
rect 33508 35436 33560 35488
rect 35440 35436 35492 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 5448 35232 5500 35284
rect 21548 35232 21600 35284
rect 23204 35232 23256 35284
rect 25044 35275 25096 35284
rect 8300 35164 8352 35216
rect 17960 35164 18012 35216
rect 25044 35241 25053 35275
rect 25053 35241 25087 35275
rect 25087 35241 25096 35275
rect 25044 35232 25096 35241
rect 25136 35275 25188 35284
rect 25136 35241 25145 35275
rect 25145 35241 25179 35275
rect 25179 35241 25188 35275
rect 25780 35275 25832 35284
rect 25136 35232 25188 35241
rect 25780 35241 25789 35275
rect 25789 35241 25823 35275
rect 25823 35241 25832 35275
rect 25780 35232 25832 35241
rect 27436 35232 27488 35284
rect 33048 35275 33100 35284
rect 33048 35241 33057 35275
rect 33057 35241 33091 35275
rect 33091 35241 33100 35275
rect 33048 35232 33100 35241
rect 15660 35139 15712 35148
rect 15660 35105 15669 35139
rect 15669 35105 15703 35139
rect 15703 35105 15712 35139
rect 15660 35096 15712 35105
rect 17500 35096 17552 35148
rect 20812 35139 20864 35148
rect 20812 35105 20821 35139
rect 20821 35105 20855 35139
rect 20855 35105 20864 35139
rect 20812 35096 20864 35105
rect 4344 35071 4396 35080
rect 4344 35037 4353 35071
rect 4353 35037 4387 35071
rect 4387 35037 4396 35071
rect 4344 35028 4396 35037
rect 8116 35028 8168 35080
rect 16672 35028 16724 35080
rect 17684 35071 17736 35080
rect 17684 35037 17693 35071
rect 17693 35037 17727 35071
rect 17727 35037 17736 35071
rect 17684 35028 17736 35037
rect 5724 34960 5776 35012
rect 16856 34960 16908 35012
rect 7104 34892 7156 34944
rect 16580 34892 16632 34944
rect 17224 34960 17276 35012
rect 18052 35028 18104 35080
rect 21456 35096 21508 35148
rect 26148 35139 26200 35148
rect 26148 35105 26157 35139
rect 26157 35105 26191 35139
rect 26191 35105 26200 35139
rect 26148 35096 26200 35105
rect 27620 35139 27672 35148
rect 27620 35105 27629 35139
rect 27629 35105 27663 35139
rect 27663 35105 27672 35139
rect 27620 35096 27672 35105
rect 20904 34960 20956 35012
rect 17132 34892 17184 34944
rect 20720 34935 20772 34944
rect 20720 34901 20729 34935
rect 20729 34901 20763 34935
rect 20763 34901 20772 34935
rect 20720 34892 20772 34901
rect 21548 34935 21600 34944
rect 21548 34901 21557 34935
rect 21557 34901 21591 34935
rect 21591 34901 21600 34935
rect 21548 34892 21600 34901
rect 23480 34960 23532 35012
rect 23664 35003 23716 35012
rect 23664 34969 23682 35003
rect 23682 34969 23716 35003
rect 23664 34960 23716 34969
rect 23848 35028 23900 35080
rect 25872 35028 25924 35080
rect 24860 34892 24912 34944
rect 26240 35071 26292 35080
rect 26240 35037 26249 35071
rect 26249 35037 26283 35071
rect 26283 35037 26292 35071
rect 26240 35028 26292 35037
rect 27528 35028 27580 35080
rect 32312 35164 32364 35216
rect 28632 35139 28684 35148
rect 28632 35105 28641 35139
rect 28641 35105 28675 35139
rect 28675 35105 28684 35139
rect 28632 35096 28684 35105
rect 33508 35139 33560 35148
rect 28724 35071 28776 35080
rect 28724 35037 28733 35071
rect 28733 35037 28767 35071
rect 28767 35037 28776 35071
rect 28724 35028 28776 35037
rect 29736 35028 29788 35080
rect 30472 35028 30524 35080
rect 29368 34960 29420 35012
rect 30196 34960 30248 35012
rect 32312 35028 32364 35080
rect 33508 35105 33517 35139
rect 33517 35105 33551 35139
rect 33551 35105 33560 35139
rect 33508 35096 33560 35105
rect 35348 35096 35400 35148
rect 27160 34892 27212 34944
rect 31208 34935 31260 34944
rect 31208 34901 31217 34935
rect 31217 34901 31251 34935
rect 31251 34901 31260 34935
rect 31208 34892 31260 34901
rect 32680 34960 32732 35012
rect 35808 35028 35860 35080
rect 35992 35028 36044 35080
rect 37004 35028 37056 35080
rect 38660 35028 38712 35080
rect 39028 35028 39080 35080
rect 39212 35071 39264 35080
rect 39212 35037 39221 35071
rect 39221 35037 39255 35071
rect 39255 35037 39264 35071
rect 39212 35028 39264 35037
rect 34704 34960 34756 35012
rect 35624 35003 35676 35012
rect 35624 34969 35633 35003
rect 35633 34969 35667 35003
rect 35667 34969 35676 35003
rect 35624 34960 35676 34969
rect 36820 34960 36872 35012
rect 36912 34960 36964 35012
rect 34428 34892 34480 34944
rect 35532 34935 35584 34944
rect 35532 34901 35541 34935
rect 35541 34901 35575 34935
rect 35575 34901 35584 34935
rect 35532 34892 35584 34901
rect 36268 34935 36320 34944
rect 36268 34901 36277 34935
rect 36277 34901 36311 34935
rect 36311 34901 36320 34935
rect 36268 34892 36320 34901
rect 37648 34892 37700 34944
rect 38936 34892 38988 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 1952 34688 2004 34740
rect 4344 34688 4396 34740
rect 5724 34731 5776 34740
rect 5724 34697 5733 34731
rect 5733 34697 5767 34731
rect 5767 34697 5776 34731
rect 5724 34688 5776 34697
rect 7748 34688 7800 34740
rect 8024 34688 8076 34740
rect 1584 34595 1636 34604
rect 1584 34561 1593 34595
rect 1593 34561 1627 34595
rect 1627 34561 1636 34595
rect 1584 34552 1636 34561
rect 4804 34552 4856 34604
rect 4988 34552 5040 34604
rect 5908 34595 5960 34604
rect 5908 34561 5917 34595
rect 5917 34561 5951 34595
rect 5951 34561 5960 34595
rect 5908 34552 5960 34561
rect 4988 34416 5040 34468
rect 5172 34484 5224 34536
rect 7748 34552 7800 34604
rect 7288 34527 7340 34536
rect 7288 34493 7297 34527
rect 7297 34493 7331 34527
rect 7331 34493 7340 34527
rect 7288 34484 7340 34493
rect 8116 34484 8168 34536
rect 9680 34688 9732 34740
rect 14464 34688 14516 34740
rect 13728 34620 13780 34672
rect 14004 34595 14056 34604
rect 14004 34561 14022 34595
rect 14022 34561 14056 34595
rect 14004 34552 14056 34561
rect 9772 34484 9824 34536
rect 16580 34688 16632 34740
rect 16856 34731 16908 34740
rect 16856 34697 16865 34731
rect 16865 34697 16899 34731
rect 16899 34697 16908 34731
rect 16856 34688 16908 34697
rect 20904 34731 20956 34740
rect 20904 34697 20913 34731
rect 20913 34697 20947 34731
rect 20947 34697 20956 34731
rect 20904 34688 20956 34697
rect 23480 34688 23532 34740
rect 23664 34731 23716 34740
rect 23664 34697 23673 34731
rect 23673 34697 23707 34731
rect 23707 34697 23716 34731
rect 23664 34688 23716 34697
rect 24952 34688 25004 34740
rect 26332 34688 26384 34740
rect 29368 34731 29420 34740
rect 29368 34697 29377 34731
rect 29377 34697 29411 34731
rect 29411 34697 29420 34731
rect 29368 34688 29420 34697
rect 35992 34731 36044 34740
rect 17500 34620 17552 34672
rect 16672 34552 16724 34604
rect 17132 34595 17184 34604
rect 17132 34561 17141 34595
rect 17141 34561 17175 34595
rect 17175 34561 17184 34595
rect 17132 34552 17184 34561
rect 18144 34552 18196 34604
rect 18420 34595 18472 34604
rect 18420 34561 18429 34595
rect 18429 34561 18463 34595
rect 18463 34561 18472 34595
rect 18420 34552 18472 34561
rect 18604 34552 18656 34604
rect 18788 34552 18840 34604
rect 19248 34552 19300 34604
rect 21548 34620 21600 34672
rect 23940 34663 23992 34672
rect 23940 34629 23949 34663
rect 23949 34629 23983 34663
rect 23983 34629 23992 34663
rect 23940 34620 23992 34629
rect 24032 34663 24084 34672
rect 24032 34629 24041 34663
rect 24041 34629 24075 34663
rect 24075 34629 24084 34663
rect 24032 34620 24084 34629
rect 25780 34620 25832 34672
rect 32312 34620 32364 34672
rect 33508 34620 33560 34672
rect 20812 34552 20864 34604
rect 21824 34552 21876 34604
rect 23756 34552 23808 34604
rect 24768 34595 24820 34604
rect 24768 34561 24777 34595
rect 24777 34561 24811 34595
rect 24811 34561 24820 34595
rect 24768 34552 24820 34561
rect 24860 34552 24912 34604
rect 27068 34552 27120 34604
rect 27160 34552 27212 34604
rect 27528 34595 27580 34604
rect 27528 34561 27537 34595
rect 27537 34561 27571 34595
rect 27571 34561 27580 34595
rect 27528 34552 27580 34561
rect 30472 34595 30524 34604
rect 30472 34561 30481 34595
rect 30481 34561 30515 34595
rect 30515 34561 30524 34595
rect 30472 34552 30524 34561
rect 30748 34595 30800 34604
rect 30748 34561 30757 34595
rect 30757 34561 30791 34595
rect 30791 34561 30800 34595
rect 30748 34552 30800 34561
rect 30932 34595 30984 34604
rect 30932 34561 30941 34595
rect 30941 34561 30975 34595
rect 30975 34561 30984 34595
rect 30932 34552 30984 34561
rect 32496 34552 32548 34604
rect 33416 34552 33468 34604
rect 33784 34552 33836 34604
rect 35992 34697 36001 34731
rect 36001 34697 36035 34731
rect 36035 34697 36044 34731
rect 35992 34688 36044 34697
rect 36912 34731 36964 34740
rect 36912 34697 36921 34731
rect 36921 34697 36955 34731
rect 36955 34697 36964 34731
rect 36912 34688 36964 34697
rect 37004 34688 37056 34740
rect 34796 34620 34848 34672
rect 35808 34663 35860 34672
rect 35808 34629 35817 34663
rect 35817 34629 35851 34663
rect 35851 34629 35860 34663
rect 35808 34620 35860 34629
rect 33968 34552 34020 34604
rect 34428 34552 34480 34604
rect 35624 34595 35676 34604
rect 9220 34416 9272 34468
rect 5172 34391 5224 34400
rect 5172 34357 5181 34391
rect 5181 34357 5215 34391
rect 5215 34357 5224 34391
rect 5172 34348 5224 34357
rect 7012 34348 7064 34400
rect 9404 34348 9456 34400
rect 12440 34348 12492 34400
rect 15384 34484 15436 34536
rect 15660 34484 15712 34536
rect 17960 34484 18012 34536
rect 18880 34484 18932 34536
rect 22008 34527 22060 34536
rect 22008 34493 22017 34527
rect 22017 34493 22051 34527
rect 22051 34493 22060 34527
rect 22008 34484 22060 34493
rect 20720 34416 20772 34468
rect 23204 34484 23256 34536
rect 26240 34484 26292 34536
rect 31024 34484 31076 34536
rect 31208 34484 31260 34536
rect 32404 34484 32456 34536
rect 35348 34484 35400 34536
rect 35624 34561 35633 34595
rect 35633 34561 35667 34595
rect 35667 34561 35676 34595
rect 35624 34552 35676 34561
rect 38752 34620 38804 34672
rect 36820 34552 36872 34604
rect 37648 34595 37700 34604
rect 37648 34561 37657 34595
rect 37657 34561 37691 34595
rect 37691 34561 37700 34595
rect 37648 34552 37700 34561
rect 34704 34459 34756 34468
rect 34704 34425 34713 34459
rect 34713 34425 34747 34459
rect 34747 34425 34756 34459
rect 34704 34416 34756 34425
rect 37556 34484 37608 34536
rect 39120 34552 39172 34604
rect 38016 34484 38068 34536
rect 18420 34391 18472 34400
rect 18420 34357 18429 34391
rect 18429 34357 18463 34391
rect 18463 34357 18472 34391
rect 18420 34348 18472 34357
rect 27252 34348 27304 34400
rect 30196 34348 30248 34400
rect 39672 34391 39724 34400
rect 39672 34357 39681 34391
rect 39681 34357 39715 34391
rect 39715 34357 39724 34391
rect 39672 34348 39724 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 14096 34144 14148 34196
rect 17500 34144 17552 34196
rect 18880 34144 18932 34196
rect 20720 34144 20772 34196
rect 27252 34187 27304 34196
rect 5172 34008 5224 34060
rect 9404 34051 9456 34060
rect 9404 34017 9413 34051
rect 9413 34017 9447 34051
rect 9447 34017 9456 34051
rect 9404 34008 9456 34017
rect 15384 34051 15436 34060
rect 15384 34017 15393 34051
rect 15393 34017 15427 34051
rect 15427 34017 15436 34051
rect 15384 34008 15436 34017
rect 4160 33983 4212 33992
rect 4160 33949 4169 33983
rect 4169 33949 4203 33983
rect 4203 33949 4212 33983
rect 4160 33940 4212 33949
rect 7012 33983 7064 33992
rect 7012 33949 7021 33983
rect 7021 33949 7055 33983
rect 7055 33949 7064 33983
rect 7012 33940 7064 33949
rect 7288 33983 7340 33992
rect 7288 33949 7297 33983
rect 7297 33949 7331 33983
rect 7331 33949 7340 33983
rect 7288 33940 7340 33949
rect 8024 33983 8076 33992
rect 8024 33949 8033 33983
rect 8033 33949 8067 33983
rect 8067 33949 8076 33983
rect 8024 33940 8076 33949
rect 9680 33983 9732 33992
rect 9680 33949 9714 33983
rect 9714 33949 9732 33983
rect 9680 33940 9732 33949
rect 12072 33983 12124 33992
rect 12072 33949 12081 33983
rect 12081 33949 12115 33983
rect 12115 33949 12124 33983
rect 12072 33940 12124 33949
rect 12440 33940 12492 33992
rect 17776 34076 17828 34128
rect 18144 34076 18196 34128
rect 19248 34076 19300 34128
rect 18420 34008 18472 34060
rect 19340 34008 19392 34060
rect 7748 33872 7800 33924
rect 17500 33983 17552 33992
rect 17500 33949 17509 33983
rect 17509 33949 17543 33983
rect 17543 33949 17552 33983
rect 17500 33940 17552 33949
rect 17776 33940 17828 33992
rect 18512 33983 18564 33992
rect 5264 33804 5316 33856
rect 6828 33847 6880 33856
rect 6828 33813 6837 33847
rect 6837 33813 6871 33847
rect 6871 33813 6880 33847
rect 6828 33804 6880 33813
rect 7380 33804 7432 33856
rect 10324 33804 10376 33856
rect 12256 33847 12308 33856
rect 12256 33813 12265 33847
rect 12265 33813 12299 33847
rect 12299 33813 12308 33847
rect 12256 33804 12308 33813
rect 12348 33804 12400 33856
rect 17316 33872 17368 33924
rect 18512 33949 18521 33983
rect 18521 33949 18555 33983
rect 18555 33949 18564 33983
rect 18512 33940 18564 33949
rect 18788 33983 18840 33992
rect 18788 33949 18797 33983
rect 18797 33949 18831 33983
rect 18831 33949 18840 33983
rect 18788 33940 18840 33949
rect 19432 33983 19484 33992
rect 19432 33949 19441 33983
rect 19441 33949 19475 33983
rect 19475 33949 19484 33983
rect 19432 33940 19484 33949
rect 27252 34153 27261 34187
rect 27261 34153 27295 34187
rect 27295 34153 27304 34187
rect 27252 34144 27304 34153
rect 27620 34187 27672 34196
rect 27620 34153 27629 34187
rect 27629 34153 27663 34187
rect 27663 34153 27672 34187
rect 27620 34144 27672 34153
rect 31208 34144 31260 34196
rect 25688 34076 25740 34128
rect 27804 34076 27856 34128
rect 35440 34119 35492 34128
rect 35440 34085 35449 34119
rect 35449 34085 35483 34119
rect 35483 34085 35492 34119
rect 35440 34076 35492 34085
rect 35532 34076 35584 34128
rect 36268 34144 36320 34196
rect 37556 34144 37608 34196
rect 39212 34144 39264 34196
rect 40316 34144 40368 34196
rect 20168 33940 20220 33992
rect 22008 33940 22060 33992
rect 23480 33940 23532 33992
rect 26608 34008 26660 34060
rect 27252 34008 27304 34060
rect 32404 34051 32456 34060
rect 32404 34017 32413 34051
rect 32413 34017 32447 34051
rect 32447 34017 32456 34051
rect 32404 34008 32456 34017
rect 27160 33983 27212 33992
rect 27160 33949 27169 33983
rect 27169 33949 27203 33983
rect 27203 33949 27212 33983
rect 27160 33940 27212 33949
rect 27436 33983 27488 33992
rect 27436 33949 27445 33983
rect 27445 33949 27479 33983
rect 27479 33949 27488 33983
rect 27436 33940 27488 33949
rect 30104 33983 30156 33992
rect 30104 33949 30113 33983
rect 30113 33949 30147 33983
rect 30147 33949 30156 33983
rect 30104 33940 30156 33949
rect 30196 33940 30248 33992
rect 30380 33983 30432 33992
rect 30380 33949 30389 33983
rect 30389 33949 30423 33983
rect 30423 33949 30432 33983
rect 30380 33940 30432 33949
rect 34796 33940 34848 33992
rect 37004 34008 37056 34060
rect 36268 33983 36320 33992
rect 21180 33915 21232 33924
rect 17776 33804 17828 33856
rect 18696 33847 18748 33856
rect 18696 33813 18705 33847
rect 18705 33813 18739 33847
rect 18739 33813 18748 33847
rect 18696 33804 18748 33813
rect 21180 33881 21189 33915
rect 21189 33881 21223 33915
rect 21223 33881 21232 33915
rect 21180 33872 21232 33881
rect 32772 33872 32824 33924
rect 36268 33949 36277 33983
rect 36277 33949 36311 33983
rect 36311 33949 36320 33983
rect 36268 33940 36320 33949
rect 39028 34076 39080 34128
rect 39948 34076 40000 34128
rect 38752 34051 38804 34060
rect 38752 34017 38761 34051
rect 38761 34017 38795 34051
rect 38795 34017 38804 34051
rect 38752 34008 38804 34017
rect 39212 34051 39264 34060
rect 39212 34017 39221 34051
rect 39221 34017 39255 34051
rect 39255 34017 39264 34051
rect 39212 34008 39264 34017
rect 39672 34008 39724 34060
rect 38936 33983 38988 33992
rect 36176 33872 36228 33924
rect 20996 33847 21048 33856
rect 20996 33813 21023 33847
rect 21023 33813 21048 33847
rect 20996 33804 21048 33813
rect 25596 33804 25648 33856
rect 30012 33804 30064 33856
rect 33416 33804 33468 33856
rect 36544 33847 36596 33856
rect 36544 33813 36553 33847
rect 36553 33813 36587 33847
rect 36587 33813 36596 33847
rect 36544 33804 36596 33813
rect 37372 33872 37424 33924
rect 38936 33949 38945 33983
rect 38945 33949 38979 33983
rect 38979 33949 38988 33983
rect 38936 33940 38988 33949
rect 39120 33983 39172 33992
rect 39120 33949 39129 33983
rect 39129 33949 39163 33983
rect 39163 33949 39172 33983
rect 39120 33940 39172 33949
rect 40408 33940 40460 33992
rect 37740 33804 37792 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 4160 33600 4212 33652
rect 5908 33600 5960 33652
rect 9772 33600 9824 33652
rect 18788 33600 18840 33652
rect 21180 33643 21232 33652
rect 21180 33609 21189 33643
rect 21189 33609 21223 33643
rect 21223 33609 21232 33643
rect 21180 33600 21232 33609
rect 27160 33600 27212 33652
rect 27436 33600 27488 33652
rect 30104 33600 30156 33652
rect 32772 33643 32824 33652
rect 32772 33609 32781 33643
rect 32781 33609 32815 33643
rect 32815 33609 32824 33643
rect 32772 33600 32824 33609
rect 7748 33532 7800 33584
rect 12256 33532 12308 33584
rect 17776 33575 17828 33584
rect 4804 33464 4856 33516
rect 4988 33507 5040 33516
rect 4988 33473 4997 33507
rect 4997 33473 5031 33507
rect 5031 33473 5040 33507
rect 4988 33464 5040 33473
rect 7196 33464 7248 33516
rect 7380 33507 7432 33516
rect 7380 33473 7389 33507
rect 7389 33473 7423 33507
rect 7423 33473 7432 33507
rect 7380 33464 7432 33473
rect 9220 33507 9272 33516
rect 9220 33473 9229 33507
rect 9229 33473 9263 33507
rect 9263 33473 9272 33507
rect 9220 33464 9272 33473
rect 10324 33507 10376 33516
rect 10324 33473 10333 33507
rect 10333 33473 10367 33507
rect 10367 33473 10376 33507
rect 10324 33464 10376 33473
rect 13176 33464 13228 33516
rect 13728 33464 13780 33516
rect 17776 33541 17785 33575
rect 17785 33541 17819 33575
rect 17819 33541 17828 33575
rect 17776 33532 17828 33541
rect 18144 33532 18196 33584
rect 18052 33464 18104 33516
rect 18512 33464 18564 33516
rect 20996 33532 21048 33584
rect 25596 33575 25648 33584
rect 25596 33541 25605 33575
rect 25605 33541 25639 33575
rect 25639 33541 25648 33575
rect 25596 33532 25648 33541
rect 25688 33575 25740 33584
rect 25688 33541 25697 33575
rect 25697 33541 25731 33575
rect 25731 33541 25740 33575
rect 25688 33532 25740 33541
rect 17684 33396 17736 33448
rect 19340 33464 19392 33516
rect 19708 33507 19760 33516
rect 19708 33473 19717 33507
rect 19717 33473 19751 33507
rect 19751 33473 19760 33507
rect 20168 33507 20220 33516
rect 19708 33464 19760 33473
rect 20168 33473 20177 33507
rect 20177 33473 20211 33507
rect 20211 33473 20220 33507
rect 20168 33464 20220 33473
rect 20444 33464 20496 33516
rect 21088 33507 21140 33516
rect 21088 33473 21097 33507
rect 21097 33473 21131 33507
rect 21131 33473 21140 33507
rect 21088 33464 21140 33473
rect 21272 33507 21324 33516
rect 21272 33473 21281 33507
rect 21281 33473 21315 33507
rect 21315 33473 21324 33507
rect 21272 33464 21324 33473
rect 24860 33464 24912 33516
rect 25780 33507 25832 33516
rect 20904 33396 20956 33448
rect 23848 33439 23900 33448
rect 23848 33405 23857 33439
rect 23857 33405 23891 33439
rect 23891 33405 23900 33439
rect 23848 33396 23900 33405
rect 17960 33328 18012 33380
rect 18512 33328 18564 33380
rect 18696 33328 18748 33380
rect 24676 33328 24728 33380
rect 25780 33473 25815 33507
rect 25815 33473 25832 33507
rect 25780 33464 25832 33473
rect 25688 33396 25740 33448
rect 26608 33507 26660 33516
rect 26608 33473 26617 33507
rect 26617 33473 26651 33507
rect 26651 33473 26660 33507
rect 26608 33464 26660 33473
rect 27252 33464 27304 33516
rect 28724 33532 28776 33584
rect 30748 33532 30800 33584
rect 26332 33396 26384 33448
rect 5264 33303 5316 33312
rect 5264 33269 5273 33303
rect 5273 33269 5307 33303
rect 5307 33269 5316 33303
rect 5264 33260 5316 33269
rect 11704 33303 11756 33312
rect 11704 33269 11713 33303
rect 11713 33269 11747 33303
rect 11747 33269 11756 33303
rect 11704 33260 11756 33269
rect 17224 33303 17276 33312
rect 17224 33269 17233 33303
rect 17233 33269 17267 33303
rect 17267 33269 17276 33303
rect 17224 33260 17276 33269
rect 18144 33303 18196 33312
rect 18144 33269 18153 33303
rect 18153 33269 18187 33303
rect 18187 33269 18196 33303
rect 18144 33260 18196 33269
rect 25228 33260 25280 33312
rect 29092 33328 29144 33380
rect 30472 33464 30524 33516
rect 31208 33464 31260 33516
rect 32956 33507 33008 33516
rect 32956 33473 32965 33507
rect 32965 33473 32999 33507
rect 32999 33473 33008 33507
rect 32956 33464 33008 33473
rect 35440 33532 35492 33584
rect 46940 33507 46992 33516
rect 46940 33473 46949 33507
rect 46949 33473 46983 33507
rect 46983 33473 46992 33507
rect 46940 33464 46992 33473
rect 36544 33396 36596 33448
rect 34612 33328 34664 33380
rect 27528 33303 27580 33312
rect 27528 33269 27537 33303
rect 27537 33269 27571 33303
rect 27571 33269 27580 33303
rect 27528 33260 27580 33269
rect 29644 33260 29696 33312
rect 46940 33328 46992 33380
rect 47032 33303 47084 33312
rect 47032 33269 47041 33303
rect 47041 33269 47075 33303
rect 47075 33269 47084 33303
rect 47032 33260 47084 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 2688 33056 2740 33108
rect 4988 32988 5040 33040
rect 3792 32852 3844 32904
rect 6000 32895 6052 32904
rect 6000 32861 6009 32895
rect 6009 32861 6043 32895
rect 6043 32861 6052 32895
rect 6000 32852 6052 32861
rect 6828 32852 6880 32904
rect 5448 32827 5500 32836
rect 5448 32793 5457 32827
rect 5457 32793 5491 32827
rect 5491 32793 5500 32827
rect 5448 32784 5500 32793
rect 21088 33056 21140 33108
rect 26332 33099 26384 33108
rect 26332 33065 26341 33099
rect 26341 33065 26375 33099
rect 26375 33065 26384 33099
rect 26332 33056 26384 33065
rect 27160 33056 27212 33108
rect 30380 33056 30432 33108
rect 31392 33056 31444 33108
rect 7196 32988 7248 33040
rect 9404 32920 9456 32972
rect 9220 32852 9272 32904
rect 11704 32852 11756 32904
rect 14280 32852 14332 32904
rect 15384 32920 15436 32972
rect 15568 32852 15620 32904
rect 19248 32852 19300 32904
rect 21272 32920 21324 32972
rect 14832 32784 14884 32836
rect 18328 32784 18380 32836
rect 19708 32784 19760 32836
rect 21180 32852 21232 32904
rect 21824 32895 21876 32904
rect 21824 32861 21833 32895
rect 21833 32861 21867 32895
rect 21867 32861 21876 32895
rect 21824 32852 21876 32861
rect 23848 32920 23900 32972
rect 24032 32852 24084 32904
rect 25228 32895 25280 32904
rect 25228 32861 25262 32895
rect 25262 32861 25280 32895
rect 25228 32852 25280 32861
rect 27436 32920 27488 32972
rect 28356 32920 28408 32972
rect 29736 32963 29788 32972
rect 29736 32929 29745 32963
rect 29745 32929 29779 32963
rect 29779 32929 29788 32963
rect 29736 32920 29788 32929
rect 32956 33056 33008 33108
rect 40408 33099 40460 33108
rect 40408 33065 40417 33099
rect 40417 33065 40451 33099
rect 40451 33065 40460 33099
rect 40408 33056 40460 33065
rect 35256 32920 35308 32972
rect 27528 32895 27580 32904
rect 27528 32861 27537 32895
rect 27537 32861 27571 32895
rect 27571 32861 27580 32895
rect 27528 32852 27580 32861
rect 30012 32895 30064 32904
rect 30012 32861 30046 32895
rect 30046 32861 30064 32895
rect 30012 32852 30064 32861
rect 33416 32895 33468 32904
rect 33416 32861 33425 32895
rect 33425 32861 33459 32895
rect 33459 32861 33468 32895
rect 33416 32852 33468 32861
rect 23388 32784 23440 32836
rect 31576 32784 31628 32836
rect 33140 32784 33192 32836
rect 36176 32852 36228 32904
rect 38936 32895 38988 32904
rect 38936 32861 38945 32895
rect 38945 32861 38979 32895
rect 38979 32861 38988 32895
rect 38936 32852 38988 32861
rect 39120 32895 39172 32904
rect 39120 32861 39129 32895
rect 39129 32861 39163 32895
rect 39163 32861 39172 32895
rect 39120 32852 39172 32861
rect 40224 32895 40276 32904
rect 40224 32861 40233 32895
rect 40233 32861 40267 32895
rect 40267 32861 40276 32895
rect 40224 32852 40276 32861
rect 41328 32852 41380 32904
rect 46756 32988 46808 33040
rect 47124 32988 47176 33040
rect 47032 32920 47084 32972
rect 46480 32895 46532 32904
rect 46480 32861 46489 32895
rect 46489 32861 46523 32895
rect 46523 32861 46532 32895
rect 46480 32852 46532 32861
rect 36360 32784 36412 32836
rect 48320 32827 48372 32836
rect 48320 32793 48329 32827
rect 48329 32793 48363 32827
rect 48363 32793 48372 32827
rect 48320 32784 48372 32793
rect 9772 32759 9824 32768
rect 9772 32725 9781 32759
rect 9781 32725 9815 32759
rect 9815 32725 9824 32759
rect 9772 32716 9824 32725
rect 10324 32716 10376 32768
rect 12164 32759 12216 32768
rect 12164 32725 12173 32759
rect 12173 32725 12207 32759
rect 12207 32725 12216 32759
rect 12164 32716 12216 32725
rect 13544 32759 13596 32768
rect 13544 32725 13553 32759
rect 13553 32725 13587 32759
rect 13587 32725 13596 32759
rect 13544 32716 13596 32725
rect 20444 32716 20496 32768
rect 22192 32716 22244 32768
rect 24124 32716 24176 32768
rect 25228 32716 25280 32768
rect 33048 32716 33100 32768
rect 33600 32716 33652 32768
rect 35532 32716 35584 32768
rect 37832 32716 37884 32768
rect 40132 32716 40184 32768
rect 45560 32716 45612 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 5448 32512 5500 32564
rect 6000 32512 6052 32564
rect 10324 32555 10376 32564
rect 10324 32521 10333 32555
rect 10333 32521 10367 32555
rect 10367 32521 10376 32555
rect 10324 32512 10376 32521
rect 12072 32512 12124 32564
rect 14556 32555 14608 32564
rect 14556 32521 14565 32555
rect 14565 32521 14599 32555
rect 14599 32521 14608 32555
rect 14556 32512 14608 32521
rect 17408 32512 17460 32564
rect 18052 32555 18104 32564
rect 18052 32521 18061 32555
rect 18061 32521 18095 32555
rect 18095 32521 18104 32555
rect 18052 32512 18104 32521
rect 24032 32512 24084 32564
rect 26240 32555 26292 32564
rect 26240 32521 26249 32555
rect 26249 32521 26283 32555
rect 26283 32521 26292 32555
rect 26240 32512 26292 32521
rect 28724 32512 28776 32564
rect 33140 32555 33192 32564
rect 33140 32521 33149 32555
rect 33149 32521 33183 32555
rect 33183 32521 33192 32555
rect 33140 32512 33192 32521
rect 33600 32555 33652 32564
rect 33600 32521 33609 32555
rect 33609 32521 33643 32555
rect 33643 32521 33652 32555
rect 33600 32512 33652 32521
rect 34612 32512 34664 32564
rect 13544 32444 13596 32496
rect 20260 32444 20312 32496
rect 1584 32419 1636 32428
rect 1584 32385 1593 32419
rect 1593 32385 1627 32419
rect 1627 32385 1636 32419
rect 1584 32376 1636 32385
rect 3792 32419 3844 32428
rect 3792 32385 3801 32419
rect 3801 32385 3835 32419
rect 3835 32385 3844 32419
rect 3792 32376 3844 32385
rect 6920 32376 6972 32428
rect 11060 32376 11112 32428
rect 13176 32419 13228 32428
rect 13176 32385 13185 32419
rect 13185 32385 13219 32419
rect 13219 32385 13228 32419
rect 13176 32376 13228 32385
rect 17224 32376 17276 32428
rect 18144 32419 18196 32428
rect 18144 32385 18153 32419
rect 18153 32385 18187 32419
rect 18187 32385 18196 32419
rect 18144 32376 18196 32385
rect 19248 32376 19300 32428
rect 3976 32351 4028 32360
rect 3976 32317 3985 32351
rect 3985 32317 4019 32351
rect 4019 32317 4028 32351
rect 3976 32308 4028 32317
rect 4068 32308 4120 32360
rect 8944 32351 8996 32360
rect 8944 32317 8953 32351
rect 8953 32317 8987 32351
rect 8987 32317 8996 32351
rect 8944 32308 8996 32317
rect 11888 32308 11940 32360
rect 15568 32351 15620 32360
rect 15568 32317 15577 32351
rect 15577 32317 15611 32351
rect 15611 32317 15620 32351
rect 15568 32308 15620 32317
rect 17592 32308 17644 32360
rect 19340 32308 19392 32360
rect 12164 32283 12216 32292
rect 12164 32249 12173 32283
rect 12173 32249 12207 32283
rect 12207 32249 12216 32283
rect 12164 32240 12216 32249
rect 15016 32215 15068 32224
rect 15016 32181 15025 32215
rect 15025 32181 15059 32215
rect 15059 32181 15068 32215
rect 15016 32172 15068 32181
rect 20168 32240 20220 32292
rect 21272 32376 21324 32428
rect 23848 32444 23900 32496
rect 22100 32376 22152 32428
rect 25044 32419 25096 32428
rect 22008 32351 22060 32360
rect 22008 32317 22017 32351
rect 22017 32317 22051 32351
rect 22051 32317 22060 32351
rect 22008 32308 22060 32317
rect 25044 32385 25053 32419
rect 25053 32385 25087 32419
rect 25087 32385 25096 32419
rect 25044 32376 25096 32385
rect 26148 32419 26200 32428
rect 26148 32385 26157 32419
rect 26157 32385 26191 32419
rect 26191 32385 26200 32419
rect 26148 32376 26200 32385
rect 26516 32376 26568 32428
rect 28356 32444 28408 32496
rect 31024 32444 31076 32496
rect 25872 32308 25924 32360
rect 31392 32419 31444 32428
rect 31392 32385 31401 32419
rect 31401 32385 31435 32419
rect 31435 32385 31444 32419
rect 31392 32376 31444 32385
rect 31668 32376 31720 32428
rect 32864 32444 32916 32496
rect 33048 32419 33100 32428
rect 33048 32385 33057 32419
rect 33057 32385 33091 32419
rect 33091 32385 33100 32419
rect 33048 32376 33100 32385
rect 34796 32376 34848 32428
rect 35256 32376 35308 32428
rect 37924 32512 37976 32564
rect 40224 32512 40276 32564
rect 36360 32487 36412 32496
rect 36360 32453 36369 32487
rect 36369 32453 36403 32487
rect 36403 32453 36412 32487
rect 36360 32444 36412 32453
rect 47768 32512 47820 32564
rect 45560 32487 45612 32496
rect 45560 32453 45569 32487
rect 45569 32453 45603 32487
rect 45603 32453 45612 32487
rect 45560 32444 45612 32453
rect 46480 32444 46532 32496
rect 35992 32376 36044 32428
rect 36176 32376 36228 32428
rect 38016 32419 38068 32428
rect 38016 32385 38025 32419
rect 38025 32385 38059 32419
rect 38059 32385 38068 32419
rect 38016 32376 38068 32385
rect 38292 32419 38344 32428
rect 38292 32385 38326 32419
rect 38326 32385 38344 32419
rect 39856 32419 39908 32428
rect 38292 32376 38344 32385
rect 39856 32385 39865 32419
rect 39865 32385 39899 32419
rect 39899 32385 39908 32419
rect 39856 32376 39908 32385
rect 40040 32419 40092 32428
rect 40040 32385 40049 32419
rect 40049 32385 40083 32419
rect 40083 32385 40092 32419
rect 40040 32376 40092 32385
rect 40316 32419 40368 32428
rect 40316 32385 40325 32419
rect 40325 32385 40359 32419
rect 40359 32385 40368 32419
rect 40316 32376 40368 32385
rect 44640 32376 44692 32428
rect 47308 32444 47360 32496
rect 31576 32308 31628 32360
rect 31760 32308 31812 32360
rect 19984 32172 20036 32224
rect 20444 32172 20496 32224
rect 34704 32308 34756 32360
rect 35624 32308 35676 32360
rect 45376 32351 45428 32360
rect 45376 32317 45385 32351
rect 45385 32317 45419 32351
rect 45419 32317 45428 32351
rect 45376 32308 45428 32317
rect 36912 32240 36964 32292
rect 21272 32215 21324 32224
rect 21272 32181 21281 32215
rect 21281 32181 21315 32215
rect 21315 32181 21324 32215
rect 21272 32172 21324 32181
rect 23388 32215 23440 32224
rect 23388 32181 23397 32215
rect 23397 32181 23431 32215
rect 23431 32181 23440 32215
rect 23388 32172 23440 32181
rect 35440 32172 35492 32224
rect 36176 32215 36228 32224
rect 36176 32181 36185 32215
rect 36185 32181 36219 32215
rect 36219 32181 36228 32215
rect 36176 32172 36228 32181
rect 39396 32215 39448 32224
rect 39396 32181 39405 32215
rect 39405 32181 39439 32215
rect 39439 32181 39448 32215
rect 39396 32172 39448 32181
rect 46020 32172 46072 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 3976 31968 4028 32020
rect 8944 31968 8996 32020
rect 11060 32011 11112 32020
rect 11060 31977 11069 32011
rect 11069 31977 11103 32011
rect 11103 31977 11112 32011
rect 11060 31968 11112 31977
rect 14280 32011 14332 32020
rect 14280 31977 14289 32011
rect 14289 31977 14323 32011
rect 14323 31977 14332 32011
rect 14280 31968 14332 31977
rect 9404 31900 9456 31952
rect 6736 31832 6788 31884
rect 7012 31875 7064 31884
rect 7012 31841 7021 31875
rect 7021 31841 7055 31875
rect 7055 31841 7064 31875
rect 7012 31832 7064 31841
rect 15016 31900 15068 31952
rect 15384 31968 15436 32020
rect 19340 31968 19392 32020
rect 20444 31968 20496 32020
rect 22100 31968 22152 32020
rect 31024 31968 31076 32020
rect 17592 31875 17644 31884
rect 17592 31841 17601 31875
rect 17601 31841 17635 31875
rect 17635 31841 17644 31875
rect 17592 31832 17644 31841
rect 22008 31832 22060 31884
rect 31300 31900 31352 31952
rect 22468 31875 22520 31884
rect 22468 31841 22477 31875
rect 22477 31841 22511 31875
rect 22511 31841 22520 31875
rect 22468 31832 22520 31841
rect 23388 31832 23440 31884
rect 31760 31875 31812 31884
rect 5448 31764 5500 31816
rect 7104 31807 7156 31816
rect 7104 31773 7113 31807
rect 7113 31773 7147 31807
rect 7147 31773 7156 31807
rect 7104 31764 7156 31773
rect 9220 31807 9272 31816
rect 9220 31773 9229 31807
rect 9229 31773 9263 31807
rect 9263 31773 9272 31807
rect 9220 31764 9272 31773
rect 10600 31807 10652 31816
rect 10600 31773 10609 31807
rect 10609 31773 10643 31807
rect 10643 31773 10652 31807
rect 10600 31764 10652 31773
rect 11888 31764 11940 31816
rect 15292 31764 15344 31816
rect 14556 31696 14608 31748
rect 15660 31696 15712 31748
rect 20168 31696 20220 31748
rect 22192 31807 22244 31816
rect 22192 31773 22201 31807
rect 22201 31773 22235 31807
rect 22235 31773 22244 31807
rect 22192 31764 22244 31773
rect 23940 31764 23992 31816
rect 25044 31807 25096 31816
rect 25044 31773 25053 31807
rect 25053 31773 25087 31807
rect 25087 31773 25096 31807
rect 25044 31764 25096 31773
rect 25780 31764 25832 31816
rect 22376 31696 22428 31748
rect 6552 31628 6604 31680
rect 16580 31671 16632 31680
rect 16580 31637 16589 31671
rect 16589 31637 16623 31671
rect 16623 31637 16632 31671
rect 17040 31671 17092 31680
rect 16580 31628 16632 31637
rect 17040 31637 17049 31671
rect 17049 31637 17083 31671
rect 17083 31637 17092 31671
rect 17040 31628 17092 31637
rect 17960 31628 18012 31680
rect 29736 31696 29788 31748
rect 31024 31764 31076 31816
rect 31760 31841 31769 31875
rect 31769 31841 31803 31875
rect 31803 31841 31812 31875
rect 31760 31832 31812 31841
rect 35624 31968 35676 32020
rect 38292 32011 38344 32020
rect 38292 31977 38301 32011
rect 38301 31977 38335 32011
rect 38335 31977 38344 32011
rect 38292 31968 38344 31977
rect 39120 31968 39172 32020
rect 41328 31968 41380 32020
rect 35348 31875 35400 31884
rect 35348 31841 35357 31875
rect 35357 31841 35391 31875
rect 35391 31841 35400 31875
rect 35348 31832 35400 31841
rect 37924 31875 37976 31884
rect 37924 31841 37933 31875
rect 37933 31841 37967 31875
rect 37967 31841 37976 31875
rect 37924 31832 37976 31841
rect 38016 31832 38068 31884
rect 40040 31875 40092 31884
rect 40040 31841 40049 31875
rect 40049 31841 40083 31875
rect 40083 31841 40092 31875
rect 40040 31832 40092 31841
rect 46020 31875 46072 31884
rect 46020 31841 46029 31875
rect 46029 31841 46063 31875
rect 46063 31841 46072 31875
rect 46020 31832 46072 31841
rect 47952 31832 48004 31884
rect 31668 31764 31720 31816
rect 35440 31764 35492 31816
rect 37556 31807 37608 31816
rect 37556 31773 37565 31807
rect 37565 31773 37599 31807
rect 37599 31773 37608 31807
rect 37556 31764 37608 31773
rect 37648 31764 37700 31816
rect 35808 31696 35860 31748
rect 25136 31628 25188 31680
rect 25688 31671 25740 31680
rect 25688 31637 25697 31671
rect 25697 31637 25731 31671
rect 25731 31637 25740 31671
rect 25688 31628 25740 31637
rect 25872 31628 25924 31680
rect 31576 31671 31628 31680
rect 31576 31637 31585 31671
rect 31585 31637 31619 31671
rect 31619 31637 31628 31671
rect 31576 31628 31628 31637
rect 34704 31628 34756 31680
rect 36084 31628 36136 31680
rect 39396 31764 39448 31816
rect 40132 31764 40184 31816
rect 45836 31807 45888 31816
rect 45836 31773 45845 31807
rect 45845 31773 45879 31807
rect 45879 31773 45888 31807
rect 45836 31764 45888 31773
rect 38016 31696 38068 31748
rect 39212 31696 39264 31748
rect 37924 31628 37976 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 6920 31356 6972 31408
rect 8024 31356 8076 31408
rect 6552 31331 6604 31340
rect 6552 31297 6561 31331
rect 6561 31297 6595 31331
rect 6595 31297 6604 31331
rect 6552 31288 6604 31297
rect 9220 31356 9272 31408
rect 11704 31288 11756 31340
rect 16580 31424 16632 31476
rect 20168 31467 20220 31476
rect 20168 31433 20177 31467
rect 20177 31433 20211 31467
rect 20211 31433 20220 31467
rect 20168 31424 20220 31433
rect 24952 31424 25004 31476
rect 25780 31467 25832 31476
rect 25780 31433 25789 31467
rect 25789 31433 25823 31467
rect 25823 31433 25832 31467
rect 25780 31424 25832 31433
rect 34796 31424 34848 31476
rect 35992 31467 36044 31476
rect 35992 31433 36001 31467
rect 36001 31433 36035 31467
rect 36035 31433 36044 31467
rect 35992 31424 36044 31433
rect 44456 31424 44508 31476
rect 45376 31424 45428 31476
rect 15292 31356 15344 31408
rect 21272 31356 21324 31408
rect 16488 31288 16540 31340
rect 17960 31288 18012 31340
rect 6092 31220 6144 31272
rect 6460 31220 6512 31272
rect 8208 31263 8260 31272
rect 8208 31229 8217 31263
rect 8217 31229 8251 31263
rect 8251 31229 8260 31263
rect 8208 31220 8260 31229
rect 13544 31263 13596 31272
rect 13544 31229 13553 31263
rect 13553 31229 13587 31263
rect 13587 31229 13596 31263
rect 13544 31220 13596 31229
rect 19340 31288 19392 31340
rect 12532 31152 12584 31204
rect 17040 31152 17092 31204
rect 17500 31152 17552 31204
rect 19984 31331 20036 31340
rect 19984 31297 19993 31331
rect 19993 31297 20027 31331
rect 20027 31297 20036 31331
rect 19984 31288 20036 31297
rect 20352 31220 20404 31272
rect 24768 31331 24820 31340
rect 24768 31297 24777 31331
rect 24777 31297 24811 31331
rect 24811 31297 24820 31331
rect 24768 31288 24820 31297
rect 25596 31288 25648 31340
rect 25688 31331 25740 31340
rect 25688 31297 25697 31331
rect 25697 31297 25731 31331
rect 25731 31297 25740 31331
rect 25688 31288 25740 31297
rect 25872 31331 25924 31340
rect 25872 31297 25881 31331
rect 25881 31297 25915 31331
rect 25915 31297 25924 31331
rect 28356 31331 28408 31340
rect 25872 31288 25924 31297
rect 28356 31297 28365 31331
rect 28365 31297 28399 31331
rect 28399 31297 28408 31331
rect 28356 31288 28408 31297
rect 28908 31288 28960 31340
rect 31024 31356 31076 31408
rect 31300 31331 31352 31340
rect 25504 31220 25556 31272
rect 22468 31152 22520 31204
rect 9220 31127 9272 31136
rect 9220 31093 9229 31127
rect 9229 31093 9263 31127
rect 9263 31093 9272 31127
rect 9220 31084 9272 31093
rect 10324 31127 10376 31136
rect 10324 31093 10333 31127
rect 10333 31093 10367 31127
rect 10367 31093 10376 31127
rect 10324 31084 10376 31093
rect 10784 31084 10836 31136
rect 15936 31127 15988 31136
rect 15936 31093 15945 31127
rect 15945 31093 15979 31127
rect 15979 31093 15988 31127
rect 15936 31084 15988 31093
rect 17868 31127 17920 31136
rect 17868 31093 17877 31127
rect 17877 31093 17911 31127
rect 17911 31093 17920 31127
rect 17868 31084 17920 31093
rect 25228 31152 25280 31204
rect 31300 31297 31309 31331
rect 31309 31297 31343 31331
rect 31343 31297 31352 31331
rect 31300 31288 31352 31297
rect 31576 31288 31628 31340
rect 35348 31356 35400 31408
rect 36176 31356 36228 31408
rect 33968 31331 34020 31340
rect 33968 31297 34002 31331
rect 34002 31297 34020 31331
rect 35532 31331 35584 31340
rect 33968 31288 34020 31297
rect 35532 31297 35541 31331
rect 35541 31297 35575 31331
rect 35575 31297 35584 31331
rect 35532 31288 35584 31297
rect 35808 31331 35860 31340
rect 35808 31297 35817 31331
rect 35817 31297 35851 31331
rect 35851 31297 35860 31331
rect 37924 31356 37976 31408
rect 37832 31331 37884 31340
rect 35808 31288 35860 31297
rect 37832 31297 37841 31331
rect 37841 31297 37875 31331
rect 37875 31297 37884 31331
rect 37832 31288 37884 31297
rect 38384 31288 38436 31340
rect 39396 31356 39448 31408
rect 39212 31331 39264 31340
rect 39212 31297 39221 31331
rect 39221 31297 39255 31331
rect 39255 31297 39264 31331
rect 39212 31288 39264 31297
rect 42616 31288 42668 31340
rect 44732 31331 44784 31340
rect 44732 31297 44741 31331
rect 44741 31297 44775 31331
rect 44775 31297 44784 31331
rect 44732 31288 44784 31297
rect 37648 31220 37700 31272
rect 37740 31263 37792 31272
rect 37740 31229 37749 31263
rect 37749 31229 37783 31263
rect 37783 31229 37792 31263
rect 42892 31263 42944 31272
rect 37740 31220 37792 31229
rect 42892 31229 42901 31263
rect 42901 31229 42935 31263
rect 42935 31229 42944 31263
rect 42892 31220 42944 31229
rect 25412 31084 25464 31136
rect 29736 31127 29788 31136
rect 29736 31093 29745 31127
rect 29745 31093 29779 31127
rect 29779 31093 29788 31127
rect 29736 31084 29788 31093
rect 30288 31127 30340 31136
rect 30288 31093 30297 31127
rect 30297 31093 30331 31127
rect 30331 31093 30340 31127
rect 30288 31084 30340 31093
rect 33048 31084 33100 31136
rect 37464 31084 37516 31136
rect 39120 31127 39172 31136
rect 39120 31093 39129 31127
rect 39129 31093 39163 31127
rect 39163 31093 39172 31127
rect 39120 31084 39172 31093
rect 44916 31127 44968 31136
rect 44916 31093 44925 31127
rect 44925 31093 44959 31127
rect 44959 31093 44968 31127
rect 44916 31084 44968 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 13544 30880 13596 30932
rect 15660 30923 15712 30932
rect 15660 30889 15669 30923
rect 15669 30889 15703 30923
rect 15703 30889 15712 30923
rect 15660 30880 15712 30889
rect 28908 30923 28960 30932
rect 28908 30889 28917 30923
rect 28917 30889 28951 30923
rect 28951 30889 28960 30923
rect 28908 30880 28960 30889
rect 37556 30880 37608 30932
rect 42616 30923 42668 30932
rect 42616 30889 42625 30923
rect 42625 30889 42659 30923
rect 42659 30889 42668 30923
rect 42616 30880 42668 30889
rect 45836 30880 45888 30932
rect 42892 30812 42944 30864
rect 44088 30812 44140 30864
rect 6920 30744 6972 30796
rect 7104 30676 7156 30728
rect 9772 30744 9824 30796
rect 12348 30787 12400 30796
rect 12348 30753 12357 30787
rect 12357 30753 12391 30787
rect 12391 30753 12400 30787
rect 12348 30744 12400 30753
rect 9312 30676 9364 30728
rect 10784 30719 10836 30728
rect 10784 30685 10818 30719
rect 10818 30685 10836 30719
rect 10784 30676 10836 30685
rect 15936 30676 15988 30728
rect 17868 30676 17920 30728
rect 18420 30676 18472 30728
rect 25412 30719 25464 30728
rect 25412 30685 25421 30719
rect 25421 30685 25455 30719
rect 25455 30685 25464 30719
rect 25412 30676 25464 30685
rect 27344 30744 27396 30796
rect 34704 30744 34756 30796
rect 25964 30676 26016 30728
rect 12440 30608 12492 30660
rect 12900 30608 12952 30660
rect 25136 30608 25188 30660
rect 8392 30583 8444 30592
rect 8392 30549 8401 30583
rect 8401 30549 8435 30583
rect 8435 30549 8444 30583
rect 8392 30540 8444 30549
rect 12164 30540 12216 30592
rect 16580 30583 16632 30592
rect 16580 30549 16589 30583
rect 16589 30549 16623 30583
rect 16623 30549 16632 30583
rect 16580 30540 16632 30549
rect 23572 30540 23624 30592
rect 26240 30540 26292 30592
rect 36912 30676 36964 30728
rect 37188 30719 37240 30728
rect 37188 30685 37197 30719
rect 37197 30685 37231 30719
rect 37231 30685 37240 30719
rect 37188 30676 37240 30685
rect 37464 30719 37516 30728
rect 36084 30651 36136 30660
rect 36084 30617 36093 30651
rect 36093 30617 36127 30651
rect 36127 30617 36136 30651
rect 36084 30608 36136 30617
rect 36268 30651 36320 30660
rect 36268 30617 36277 30651
rect 36277 30617 36311 30651
rect 36311 30617 36320 30651
rect 36268 30608 36320 30617
rect 37464 30685 37473 30719
rect 37473 30685 37507 30719
rect 37507 30685 37516 30719
rect 37464 30676 37516 30685
rect 44456 30719 44508 30728
rect 37924 30608 37976 30660
rect 29828 30540 29880 30592
rect 30196 30583 30248 30592
rect 30196 30549 30205 30583
rect 30205 30549 30239 30583
rect 30239 30549 30248 30583
rect 30196 30540 30248 30549
rect 37832 30540 37884 30592
rect 41236 30540 41288 30592
rect 42800 30540 42852 30592
rect 44456 30685 44465 30719
rect 44465 30685 44499 30719
rect 44499 30685 44508 30719
rect 44456 30676 44508 30685
rect 44180 30608 44232 30660
rect 44548 30608 44600 30660
rect 44916 30676 44968 30728
rect 45836 30608 45888 30660
rect 43536 30583 43588 30592
rect 43536 30549 43545 30583
rect 43545 30549 43579 30583
rect 43579 30549 43588 30583
rect 43536 30540 43588 30549
rect 43720 30540 43772 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 11704 30379 11756 30388
rect 11704 30345 11713 30379
rect 11713 30345 11747 30379
rect 11747 30345 11756 30379
rect 11704 30336 11756 30345
rect 12900 30379 12952 30388
rect 12900 30345 12909 30379
rect 12909 30345 12943 30379
rect 12943 30345 12952 30379
rect 12900 30336 12952 30345
rect 9220 30200 9272 30252
rect 10324 30268 10376 30320
rect 13084 30243 13136 30252
rect 6552 30132 6604 30184
rect 12164 30175 12216 30184
rect 12164 30141 12173 30175
rect 12173 30141 12207 30175
rect 12207 30141 12216 30175
rect 12164 30132 12216 30141
rect 13084 30209 13093 30243
rect 13093 30209 13127 30243
rect 13127 30209 13136 30243
rect 13084 30200 13136 30209
rect 15476 30200 15528 30252
rect 18328 30268 18380 30320
rect 30196 30336 30248 30388
rect 40132 30379 40184 30388
rect 40132 30345 40147 30379
rect 40147 30345 40181 30379
rect 40181 30345 40184 30379
rect 40132 30336 40184 30345
rect 44180 30379 44232 30388
rect 44180 30345 44189 30379
rect 44189 30345 44223 30379
rect 44223 30345 44232 30379
rect 44180 30336 44232 30345
rect 22100 30200 22152 30252
rect 10600 30064 10652 30116
rect 16580 30132 16632 30184
rect 17868 30132 17920 30184
rect 18420 30175 18472 30184
rect 18420 30141 18429 30175
rect 18429 30141 18463 30175
rect 18463 30141 18472 30175
rect 18420 30132 18472 30141
rect 22008 30132 22060 30184
rect 23296 30243 23348 30252
rect 23296 30209 23330 30243
rect 23330 30209 23348 30243
rect 23296 30200 23348 30209
rect 22468 30175 22520 30184
rect 22468 30141 22477 30175
rect 22477 30141 22511 30175
rect 22511 30141 22520 30175
rect 25780 30243 25832 30252
rect 25780 30209 25789 30243
rect 25789 30209 25823 30243
rect 25823 30209 25832 30243
rect 25780 30200 25832 30209
rect 27344 30243 27396 30252
rect 27344 30209 27353 30243
rect 27353 30209 27387 30243
rect 27387 30209 27396 30243
rect 27344 30200 27396 30209
rect 29736 30200 29788 30252
rect 32496 30243 32548 30252
rect 32496 30209 32505 30243
rect 32505 30209 32539 30243
rect 32539 30209 32548 30243
rect 32496 30200 32548 30209
rect 32680 30200 32732 30252
rect 34336 30243 34388 30252
rect 34336 30209 34345 30243
rect 34345 30209 34379 30243
rect 34379 30209 34388 30243
rect 34336 30200 34388 30209
rect 34612 30243 34664 30252
rect 34612 30209 34621 30243
rect 34621 30209 34655 30243
rect 34655 30209 34664 30243
rect 34612 30200 34664 30209
rect 22468 30132 22520 30141
rect 25964 30132 26016 30184
rect 27528 30175 27580 30184
rect 27528 30141 27537 30175
rect 27537 30141 27571 30175
rect 27571 30141 27580 30175
rect 27528 30132 27580 30141
rect 30288 30132 30340 30184
rect 31944 30132 31996 30184
rect 32772 30175 32824 30184
rect 32772 30141 32781 30175
rect 32781 30141 32815 30175
rect 32815 30141 32824 30175
rect 32772 30132 32824 30141
rect 34796 30243 34848 30252
rect 34796 30209 34805 30243
rect 34805 30209 34839 30243
rect 34839 30209 34848 30243
rect 34796 30200 34848 30209
rect 35440 30243 35492 30252
rect 35440 30209 35449 30243
rect 35449 30209 35483 30243
rect 35483 30209 35492 30243
rect 35440 30200 35492 30209
rect 6736 29996 6788 30048
rect 9312 29996 9364 30048
rect 12440 30064 12492 30116
rect 18328 30064 18380 30116
rect 15384 30039 15436 30048
rect 15384 30005 15393 30039
rect 15393 30005 15427 30039
rect 15427 30005 15436 30039
rect 15384 29996 15436 30005
rect 21548 29996 21600 30048
rect 22376 30039 22428 30048
rect 22376 30005 22385 30039
rect 22385 30005 22419 30039
rect 22419 30005 22428 30039
rect 22376 29996 22428 30005
rect 24860 30064 24912 30116
rect 25780 30064 25832 30116
rect 29000 30064 29052 30116
rect 31576 30064 31628 30116
rect 33232 30064 33284 30116
rect 34612 30064 34664 30116
rect 36452 30200 36504 30252
rect 37740 30200 37792 30252
rect 38292 30200 38344 30252
rect 39120 30268 39172 30320
rect 38844 30200 38896 30252
rect 38384 30175 38436 30184
rect 38384 30141 38393 30175
rect 38393 30141 38427 30175
rect 38427 30141 38436 30175
rect 38384 30132 38436 30141
rect 39212 30132 39264 30184
rect 39488 30175 39540 30184
rect 39488 30141 39497 30175
rect 39497 30141 39531 30175
rect 39531 30141 39540 30175
rect 39488 30132 39540 30141
rect 40684 30200 40736 30252
rect 40776 30243 40828 30252
rect 40776 30209 40785 30243
rect 40785 30209 40819 30243
rect 40819 30209 40828 30243
rect 40776 30200 40828 30209
rect 40592 30132 40644 30184
rect 41328 30200 41380 30252
rect 44548 30311 44600 30320
rect 44548 30277 44557 30311
rect 44557 30277 44591 30311
rect 44591 30277 44600 30311
rect 44548 30268 44600 30277
rect 43352 30243 43404 30252
rect 43352 30209 43361 30243
rect 43361 30209 43395 30243
rect 43395 30209 43404 30243
rect 43352 30200 43404 30209
rect 44180 30200 44232 30252
rect 47768 30243 47820 30252
rect 47768 30209 47777 30243
rect 47777 30209 47811 30243
rect 47811 30209 47820 30243
rect 47768 30200 47820 30209
rect 43444 30132 43496 30184
rect 24768 29996 24820 30048
rect 25412 29996 25464 30048
rect 32312 30039 32364 30048
rect 32312 30005 32321 30039
rect 32321 30005 32355 30039
rect 32355 30005 32364 30039
rect 32312 29996 32364 30005
rect 34060 29996 34112 30048
rect 34704 29996 34756 30048
rect 36636 29996 36688 30048
rect 38844 30039 38896 30048
rect 38844 30005 38853 30039
rect 38853 30005 38887 30039
rect 38887 30005 38896 30039
rect 38844 29996 38896 30005
rect 38936 29996 38988 30048
rect 40224 30064 40276 30116
rect 43168 30064 43220 30116
rect 43352 30064 43404 30116
rect 43260 29996 43312 30048
rect 43904 29996 43956 30048
rect 46480 29996 46532 30048
rect 47860 30039 47912 30048
rect 47860 30005 47869 30039
rect 47869 30005 47903 30039
rect 47903 30005 47912 30039
rect 47860 29996 47912 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 5172 29792 5224 29844
rect 6828 29792 6880 29844
rect 204 29724 256 29776
rect 13084 29767 13136 29776
rect 6736 29699 6788 29708
rect 6736 29665 6745 29699
rect 6745 29665 6779 29699
rect 6779 29665 6788 29699
rect 6736 29656 6788 29665
rect 13084 29733 13093 29767
rect 13093 29733 13127 29767
rect 13127 29733 13136 29767
rect 13084 29724 13136 29733
rect 17500 29767 17552 29776
rect 17500 29733 17509 29767
rect 17509 29733 17543 29767
rect 17543 29733 17552 29767
rect 17500 29724 17552 29733
rect 23296 29767 23348 29776
rect 23296 29733 23305 29767
rect 23305 29733 23339 29767
rect 23339 29733 23348 29767
rect 23296 29724 23348 29733
rect 12164 29656 12216 29708
rect 12440 29699 12492 29708
rect 12440 29665 12449 29699
rect 12449 29665 12483 29699
rect 12483 29665 12492 29699
rect 12440 29656 12492 29665
rect 17776 29656 17828 29708
rect 19248 29656 19300 29708
rect 10600 29588 10652 29640
rect 14280 29631 14332 29640
rect 14280 29597 14289 29631
rect 14289 29597 14323 29631
rect 14323 29597 14332 29631
rect 14280 29588 14332 29597
rect 14740 29588 14792 29640
rect 18420 29588 18472 29640
rect 18604 29588 18656 29640
rect 20904 29656 20956 29708
rect 22468 29656 22520 29708
rect 24952 29656 25004 29708
rect 25504 29724 25556 29776
rect 27344 29767 27396 29776
rect 27344 29733 27353 29767
rect 27353 29733 27387 29767
rect 27387 29733 27396 29767
rect 27344 29724 27396 29733
rect 32864 29767 32916 29776
rect 32864 29733 32873 29767
rect 32873 29733 32907 29767
rect 32907 29733 32916 29767
rect 32864 29724 32916 29733
rect 33968 29724 34020 29776
rect 44732 29792 44784 29844
rect 44640 29724 44692 29776
rect 25412 29699 25464 29708
rect 25412 29665 25421 29699
rect 25421 29665 25455 29699
rect 25455 29665 25464 29699
rect 25412 29656 25464 29665
rect 25964 29699 26016 29708
rect 25964 29665 25973 29699
rect 25973 29665 26007 29699
rect 26007 29665 26016 29699
rect 25964 29656 26016 29665
rect 29644 29656 29696 29708
rect 20628 29588 20680 29640
rect 22008 29588 22060 29640
rect 23480 29631 23532 29640
rect 23480 29597 23489 29631
rect 23489 29597 23523 29631
rect 23523 29597 23532 29631
rect 23480 29588 23532 29597
rect 24768 29588 24820 29640
rect 25780 29588 25832 29640
rect 26240 29631 26292 29640
rect 26240 29597 26274 29631
rect 26274 29597 26292 29631
rect 26240 29588 26292 29597
rect 29828 29588 29880 29640
rect 30104 29588 30156 29640
rect 31024 29588 31076 29640
rect 35348 29656 35400 29708
rect 34060 29631 34112 29640
rect 34060 29597 34069 29631
rect 34069 29597 34103 29631
rect 34103 29597 34112 29631
rect 34060 29588 34112 29597
rect 6920 29563 6972 29572
rect 6920 29529 6929 29563
rect 6929 29529 6963 29563
rect 6963 29529 6972 29563
rect 6920 29520 6972 29529
rect 10232 29452 10284 29504
rect 12624 29495 12676 29504
rect 12624 29461 12633 29495
rect 12633 29461 12667 29495
rect 12667 29461 12676 29495
rect 12624 29452 12676 29461
rect 14464 29495 14516 29504
rect 14464 29461 14473 29495
rect 14473 29461 14507 29495
rect 14507 29461 14516 29495
rect 14464 29452 14516 29461
rect 15384 29520 15436 29572
rect 17868 29563 17920 29572
rect 17868 29529 17877 29563
rect 17877 29529 17911 29563
rect 17911 29529 17920 29563
rect 17868 29520 17920 29529
rect 21548 29563 21600 29572
rect 17224 29452 17276 29504
rect 19984 29452 20036 29504
rect 21548 29529 21582 29563
rect 21582 29529 21600 29563
rect 21548 29520 21600 29529
rect 23572 29452 23624 29504
rect 23848 29452 23900 29504
rect 25044 29452 25096 29504
rect 27620 29452 27672 29504
rect 29092 29452 29144 29504
rect 30472 29452 30524 29504
rect 32312 29520 32364 29572
rect 33508 29520 33560 29572
rect 34336 29631 34388 29640
rect 34336 29597 34345 29631
rect 34345 29597 34379 29631
rect 34379 29597 34388 29631
rect 37372 29656 37424 29708
rect 40040 29699 40092 29708
rect 34336 29588 34388 29597
rect 36452 29588 36504 29640
rect 37832 29631 37884 29640
rect 37832 29597 37841 29631
rect 37841 29597 37875 29631
rect 37875 29597 37884 29631
rect 37832 29588 37884 29597
rect 38016 29631 38068 29640
rect 38016 29597 38025 29631
rect 38025 29597 38059 29631
rect 38059 29597 38068 29631
rect 38016 29588 38068 29597
rect 38936 29588 38988 29640
rect 39120 29631 39172 29640
rect 39120 29597 39129 29631
rect 39129 29597 39163 29631
rect 39163 29597 39172 29631
rect 39120 29588 39172 29597
rect 39488 29588 39540 29640
rect 40040 29665 40049 29699
rect 40049 29665 40083 29699
rect 40083 29665 40092 29699
rect 40040 29656 40092 29665
rect 42984 29656 43036 29708
rect 43536 29656 43588 29708
rect 46480 29699 46532 29708
rect 46480 29665 46489 29699
rect 46489 29665 46523 29699
rect 46523 29665 46532 29699
rect 46480 29656 46532 29665
rect 47860 29656 47912 29708
rect 40776 29588 40828 29640
rect 42892 29631 42944 29640
rect 34796 29520 34848 29572
rect 33324 29452 33376 29504
rect 33416 29452 33468 29504
rect 38660 29452 38712 29504
rect 38844 29452 38896 29504
rect 40500 29452 40552 29504
rect 42892 29597 42901 29631
rect 42901 29597 42935 29631
rect 42935 29597 42944 29631
rect 42892 29588 42944 29597
rect 43444 29588 43496 29640
rect 43904 29631 43956 29640
rect 43904 29597 43913 29631
rect 43913 29597 43947 29631
rect 43947 29597 43956 29631
rect 43904 29588 43956 29597
rect 44180 29520 44232 29572
rect 48320 29563 48372 29572
rect 48320 29529 48329 29563
rect 48329 29529 48363 29563
rect 48363 29529 48372 29563
rect 48320 29520 48372 29529
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 6920 29248 6972 29300
rect 13268 29248 13320 29300
rect 15476 29291 15528 29300
rect 8392 29223 8444 29232
rect 8392 29189 8426 29223
rect 8426 29189 8444 29223
rect 8392 29180 8444 29189
rect 14464 29223 14516 29232
rect 14464 29189 14482 29223
rect 14482 29189 14516 29223
rect 15476 29257 15485 29291
rect 15485 29257 15519 29291
rect 15519 29257 15528 29291
rect 15476 29248 15528 29257
rect 15660 29248 15712 29300
rect 29644 29248 29696 29300
rect 29828 29291 29880 29300
rect 29828 29257 29837 29291
rect 29837 29257 29871 29291
rect 29871 29257 29880 29291
rect 29828 29248 29880 29257
rect 33324 29248 33376 29300
rect 34152 29248 34204 29300
rect 14464 29180 14516 29189
rect 5632 29155 5684 29164
rect 5632 29121 5641 29155
rect 5641 29121 5675 29155
rect 5675 29121 5684 29155
rect 5632 29112 5684 29121
rect 6828 29112 6880 29164
rect 15660 29155 15712 29164
rect 15660 29121 15669 29155
rect 15669 29121 15703 29155
rect 15703 29121 15712 29155
rect 15660 29112 15712 29121
rect 16856 29112 16908 29164
rect 19432 29180 19484 29232
rect 8116 29087 8168 29096
rect 8116 29053 8125 29087
rect 8125 29053 8159 29087
rect 8159 29053 8168 29087
rect 8116 29044 8168 29053
rect 14740 29087 14792 29096
rect 14740 29053 14749 29087
rect 14749 29053 14783 29087
rect 14783 29053 14792 29087
rect 14740 29044 14792 29053
rect 6920 28976 6972 29028
rect 12716 28976 12768 29028
rect 9496 28951 9548 28960
rect 9496 28917 9505 28951
rect 9505 28917 9539 28951
rect 9539 28917 9548 28951
rect 9496 28908 9548 28917
rect 13544 28908 13596 28960
rect 19340 29155 19392 29164
rect 19340 29121 19349 29155
rect 19349 29121 19383 29155
rect 19383 29121 19392 29155
rect 19340 29112 19392 29121
rect 32036 29180 32088 29232
rect 32404 29180 32456 29232
rect 20076 29155 20128 29164
rect 20076 29121 20110 29155
rect 20110 29121 20128 29155
rect 20076 29112 20128 29121
rect 20628 29112 20680 29164
rect 22100 29112 22152 29164
rect 22560 29112 22612 29164
rect 23572 29112 23624 29164
rect 24768 29112 24820 29164
rect 22928 29044 22980 29096
rect 24400 29087 24452 29096
rect 24400 29053 24409 29087
rect 24409 29053 24443 29087
rect 24443 29053 24452 29087
rect 24400 29044 24452 29053
rect 24860 29044 24912 29096
rect 25504 29112 25556 29164
rect 27528 29155 27580 29164
rect 25780 29044 25832 29096
rect 27528 29121 27537 29155
rect 27537 29121 27571 29155
rect 27571 29121 27580 29155
rect 27528 29112 27580 29121
rect 30472 29155 30524 29164
rect 30472 29121 30481 29155
rect 30481 29121 30515 29155
rect 30515 29121 30524 29155
rect 30472 29112 30524 29121
rect 30932 29112 30984 29164
rect 31024 29112 31076 29164
rect 32680 29112 32732 29164
rect 27344 29044 27396 29096
rect 30656 29087 30708 29096
rect 23756 28976 23808 29028
rect 25596 29019 25648 29028
rect 25596 28985 25605 29019
rect 25605 28985 25639 29019
rect 25639 28985 25648 29019
rect 25596 28976 25648 28985
rect 18328 28908 18380 28960
rect 18604 28908 18656 28960
rect 21180 28951 21232 28960
rect 21180 28917 21189 28951
rect 21189 28917 21223 28951
rect 21223 28917 21232 28951
rect 21180 28908 21232 28917
rect 30656 29053 30665 29087
rect 30665 29053 30699 29087
rect 30699 29053 30708 29087
rect 30656 29044 30708 29053
rect 32956 29155 33008 29164
rect 32956 29121 32965 29155
rect 32965 29121 32999 29155
rect 32999 29121 33008 29155
rect 33508 29155 33560 29164
rect 32956 29112 33008 29121
rect 33508 29121 33517 29155
rect 33517 29121 33551 29155
rect 33551 29121 33560 29155
rect 33508 29112 33560 29121
rect 35348 29180 35400 29232
rect 37280 29180 37332 29232
rect 38016 29180 38068 29232
rect 40224 29180 40276 29232
rect 40684 29223 40736 29232
rect 40684 29189 40693 29223
rect 40693 29189 40727 29223
rect 40727 29189 40736 29223
rect 40684 29180 40736 29189
rect 43536 29180 43588 29232
rect 30104 28976 30156 29028
rect 33232 29044 33284 29096
rect 33416 29087 33468 29096
rect 33416 29053 33425 29087
rect 33425 29053 33459 29087
rect 33459 29053 33468 29087
rect 33416 29044 33468 29053
rect 31576 28976 31628 29028
rect 35440 29112 35492 29164
rect 36636 29155 36688 29164
rect 36636 29121 36645 29155
rect 36645 29121 36679 29155
rect 36679 29121 36688 29155
rect 36636 29112 36688 29121
rect 36268 29044 36320 29096
rect 38292 29112 38344 29164
rect 38660 29112 38712 29164
rect 40592 29155 40644 29164
rect 28816 28908 28868 28960
rect 32496 28908 32548 28960
rect 37924 28976 37976 29028
rect 38292 28976 38344 29028
rect 38384 28976 38436 29028
rect 40592 29121 40601 29155
rect 40601 29121 40635 29155
rect 40635 29121 40644 29155
rect 40592 29112 40644 29121
rect 40776 29155 40828 29164
rect 40776 29121 40785 29155
rect 40785 29121 40819 29155
rect 40819 29121 40828 29155
rect 40776 29112 40828 29121
rect 42800 29112 42852 29164
rect 43720 29155 43772 29164
rect 43720 29121 43729 29155
rect 43729 29121 43763 29155
rect 43763 29121 43772 29155
rect 43720 29112 43772 29121
rect 47308 29112 47360 29164
rect 39212 29044 39264 29096
rect 43168 29044 43220 29096
rect 43260 29044 43312 29096
rect 43904 29044 43956 29096
rect 40224 28976 40276 29028
rect 40684 28976 40736 29028
rect 43352 29019 43404 29028
rect 43352 28985 43361 29019
rect 43361 28985 43395 29019
rect 43395 28985 43404 29019
rect 43352 28976 43404 28985
rect 44640 28976 44692 29028
rect 46204 28976 46256 29028
rect 48320 28976 48372 29028
rect 38476 28908 38528 28960
rect 39120 28908 39172 28960
rect 46480 28908 46532 28960
rect 47124 28951 47176 28960
rect 47124 28917 47133 28951
rect 47133 28917 47167 28951
rect 47167 28917 47176 28951
rect 47124 28908 47176 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 8116 28747 8168 28756
rect 8116 28713 8125 28747
rect 8125 28713 8159 28747
rect 8159 28713 8168 28747
rect 8116 28704 8168 28713
rect 14280 28704 14332 28756
rect 16856 28747 16908 28756
rect 16856 28713 16865 28747
rect 16865 28713 16899 28747
rect 16899 28713 16908 28747
rect 16856 28704 16908 28713
rect 12164 28679 12216 28688
rect 12164 28645 12173 28679
rect 12173 28645 12207 28679
rect 12207 28645 12216 28679
rect 12164 28636 12216 28645
rect 5540 28611 5592 28620
rect 5540 28577 5549 28611
rect 5549 28577 5583 28611
rect 5583 28577 5592 28611
rect 5540 28568 5592 28577
rect 6920 28611 6972 28620
rect 6920 28577 6929 28611
rect 6929 28577 6963 28611
rect 6963 28577 6972 28611
rect 6920 28568 6972 28577
rect 7104 28611 7156 28620
rect 7104 28577 7113 28611
rect 7113 28577 7147 28611
rect 7147 28577 7156 28611
rect 7104 28568 7156 28577
rect 9496 28568 9548 28620
rect 8024 28500 8076 28552
rect 9312 28500 9364 28552
rect 13728 28568 13780 28620
rect 17776 28704 17828 28756
rect 19432 28747 19484 28756
rect 19432 28713 19441 28747
rect 19441 28713 19475 28747
rect 19475 28713 19484 28747
rect 19432 28704 19484 28713
rect 20444 28704 20496 28756
rect 22376 28704 22428 28756
rect 23480 28704 23532 28756
rect 24400 28704 24452 28756
rect 31484 28704 31536 28756
rect 32220 28704 32272 28756
rect 33416 28704 33468 28756
rect 17776 28568 17828 28620
rect 11888 28432 11940 28484
rect 13544 28475 13596 28484
rect 13544 28441 13553 28475
rect 13553 28441 13587 28475
rect 13587 28441 13596 28475
rect 13544 28432 13596 28441
rect 14648 28500 14700 28552
rect 17224 28543 17276 28552
rect 17224 28509 17233 28543
rect 17233 28509 17267 28543
rect 17267 28509 17276 28543
rect 17224 28500 17276 28509
rect 18236 28543 18288 28552
rect 18236 28509 18245 28543
rect 18245 28509 18279 28543
rect 18279 28509 18288 28543
rect 18236 28500 18288 28509
rect 18328 28543 18380 28552
rect 18328 28509 18337 28543
rect 18337 28509 18371 28543
rect 18371 28509 18380 28543
rect 18604 28543 18656 28552
rect 18328 28500 18380 28509
rect 18604 28509 18613 28543
rect 18613 28509 18647 28543
rect 18647 28509 18656 28543
rect 18604 28500 18656 28509
rect 19984 28568 20036 28620
rect 20904 28568 20956 28620
rect 22560 28568 22612 28620
rect 18420 28475 18472 28484
rect 9128 28407 9180 28416
rect 9128 28373 9137 28407
rect 9137 28373 9171 28407
rect 9171 28373 9180 28407
rect 9128 28364 9180 28373
rect 12716 28364 12768 28416
rect 12900 28407 12952 28416
rect 12900 28373 12909 28407
rect 12909 28373 12943 28407
rect 12943 28373 12952 28407
rect 12900 28364 12952 28373
rect 18420 28441 18429 28475
rect 18429 28441 18463 28475
rect 18463 28441 18472 28475
rect 18420 28432 18472 28441
rect 19432 28432 19484 28484
rect 20628 28500 20680 28552
rect 23756 28611 23808 28620
rect 23756 28577 23765 28611
rect 23765 28577 23799 28611
rect 23799 28577 23808 28611
rect 23756 28568 23808 28577
rect 21180 28500 21232 28552
rect 22376 28543 22428 28552
rect 22376 28509 22385 28543
rect 22385 28509 22419 28543
rect 22419 28509 22428 28543
rect 22376 28500 22428 28509
rect 22652 28543 22704 28552
rect 22652 28509 22661 28543
rect 22661 28509 22695 28543
rect 22695 28509 22704 28543
rect 22652 28500 22704 28509
rect 23572 28500 23624 28552
rect 24124 28500 24176 28552
rect 25872 28568 25924 28620
rect 29092 28568 29144 28620
rect 24860 28500 24912 28552
rect 29920 28543 29972 28552
rect 29920 28509 29929 28543
rect 29929 28509 29963 28543
rect 29963 28509 29972 28543
rect 29920 28500 29972 28509
rect 30656 28568 30708 28620
rect 31576 28568 31628 28620
rect 35348 28704 35400 28756
rect 36452 28747 36504 28756
rect 36452 28713 36461 28747
rect 36461 28713 36495 28747
rect 36495 28713 36504 28747
rect 36452 28704 36504 28713
rect 38292 28747 38344 28756
rect 38292 28713 38301 28747
rect 38301 28713 38335 28747
rect 38335 28713 38344 28747
rect 38292 28704 38344 28713
rect 38660 28704 38712 28756
rect 37188 28636 37240 28688
rect 40316 28679 40368 28688
rect 40316 28645 40325 28679
rect 40325 28645 40359 28679
rect 40359 28645 40368 28679
rect 40316 28636 40368 28645
rect 31484 28500 31536 28552
rect 33048 28543 33100 28552
rect 32220 28432 32272 28484
rect 33048 28509 33057 28543
rect 33057 28509 33091 28543
rect 33091 28509 33100 28543
rect 33048 28500 33100 28509
rect 33232 28500 33284 28552
rect 37372 28543 37424 28552
rect 33324 28475 33376 28484
rect 18052 28407 18104 28416
rect 18052 28373 18061 28407
rect 18061 28373 18095 28407
rect 18095 28373 18104 28407
rect 18052 28364 18104 28373
rect 20260 28364 20312 28416
rect 22284 28364 22336 28416
rect 23388 28364 23440 28416
rect 29736 28407 29788 28416
rect 29736 28373 29745 28407
rect 29745 28373 29779 28407
rect 29779 28373 29788 28407
rect 29736 28364 29788 28373
rect 33324 28441 33333 28475
rect 33333 28441 33367 28475
rect 33367 28441 33376 28475
rect 33324 28432 33376 28441
rect 33416 28475 33468 28484
rect 33416 28441 33425 28475
rect 33425 28441 33459 28475
rect 33459 28441 33468 28475
rect 33416 28432 33468 28441
rect 34980 28432 35032 28484
rect 37372 28509 37381 28543
rect 37381 28509 37415 28543
rect 37415 28509 37424 28543
rect 37372 28500 37424 28509
rect 38476 28543 38528 28552
rect 38476 28509 38489 28543
rect 38489 28509 38523 28543
rect 38523 28509 38528 28543
rect 38476 28500 38528 28509
rect 37464 28432 37516 28484
rect 38660 28509 38669 28530
rect 38669 28509 38703 28530
rect 38703 28509 38712 28530
rect 38660 28478 38712 28509
rect 39120 28500 39172 28552
rect 40132 28568 40184 28620
rect 42064 28568 42116 28620
rect 43352 28568 43404 28620
rect 46480 28611 46532 28620
rect 46480 28577 46489 28611
rect 46489 28577 46523 28611
rect 46523 28577 46532 28611
rect 46480 28568 46532 28577
rect 47124 28568 47176 28620
rect 48228 28611 48280 28620
rect 48228 28577 48237 28611
rect 48237 28577 48271 28611
rect 48271 28577 48280 28611
rect 48228 28568 48280 28577
rect 40224 28500 40276 28552
rect 40408 28500 40460 28552
rect 40500 28432 40552 28484
rect 42800 28500 42852 28552
rect 43720 28500 43772 28552
rect 43904 28543 43956 28552
rect 43904 28509 43913 28543
rect 43913 28509 43947 28543
rect 43947 28509 43956 28543
rect 43904 28500 43956 28509
rect 43812 28432 43864 28484
rect 37556 28407 37608 28416
rect 37556 28373 37565 28407
rect 37565 28373 37599 28407
rect 37599 28373 37608 28407
rect 37556 28364 37608 28373
rect 41788 28364 41840 28416
rect 43536 28364 43588 28416
rect 43996 28364 44048 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 12624 28160 12676 28212
rect 17132 28160 17184 28212
rect 18604 28160 18656 28212
rect 20076 28203 20128 28212
rect 20076 28169 20085 28203
rect 20085 28169 20119 28203
rect 20119 28169 20128 28203
rect 20076 28160 20128 28169
rect 23388 28203 23440 28212
rect 23388 28169 23397 28203
rect 23397 28169 23431 28203
rect 23431 28169 23440 28203
rect 23388 28160 23440 28169
rect 30380 28160 30432 28212
rect 33416 28160 33468 28212
rect 34980 28203 35032 28212
rect 34980 28169 34989 28203
rect 34989 28169 35023 28203
rect 35023 28169 35032 28203
rect 34980 28160 35032 28169
rect 42800 28203 42852 28212
rect 42800 28169 42809 28203
rect 42809 28169 42843 28203
rect 42843 28169 42852 28203
rect 42800 28160 42852 28169
rect 43168 28203 43220 28212
rect 43168 28169 43177 28203
rect 43177 28169 43211 28203
rect 43211 28169 43220 28203
rect 43168 28160 43220 28169
rect 43812 28160 43864 28212
rect 12900 28135 12952 28144
rect 12900 28101 12918 28135
rect 12918 28101 12952 28135
rect 12900 28092 12952 28101
rect 18420 28092 18472 28144
rect 7196 28024 7248 28076
rect 9128 28067 9180 28076
rect 9128 28033 9137 28067
rect 9137 28033 9171 28067
rect 9171 28033 9180 28067
rect 9128 28024 9180 28033
rect 9220 28024 9272 28076
rect 14740 28024 14792 28076
rect 17408 28024 17460 28076
rect 20260 28067 20312 28076
rect 20260 28033 20269 28067
rect 20269 28033 20303 28067
rect 20303 28033 20312 28067
rect 20260 28024 20312 28033
rect 20444 28067 20496 28076
rect 20444 28033 20453 28067
rect 20453 28033 20487 28067
rect 20487 28033 20496 28067
rect 20444 28024 20496 28033
rect 22284 28067 22336 28076
rect 22284 28033 22318 28067
rect 22318 28033 22336 28067
rect 22284 28024 22336 28033
rect 22652 28092 22704 28144
rect 25044 28024 25096 28076
rect 25412 28067 25464 28076
rect 25412 28033 25421 28067
rect 25421 28033 25455 28067
rect 25455 28033 25464 28067
rect 25412 28024 25464 28033
rect 27804 28024 27856 28076
rect 29736 28092 29788 28144
rect 37556 28092 37608 28144
rect 39212 28092 39264 28144
rect 40040 28092 40092 28144
rect 40684 28135 40736 28144
rect 40684 28101 40693 28135
rect 40693 28101 40727 28135
rect 40727 28101 40736 28135
rect 40684 28092 40736 28101
rect 30932 28024 30984 28076
rect 34704 28024 34756 28076
rect 40132 28024 40184 28076
rect 42064 28024 42116 28076
rect 7012 27956 7064 28008
rect 10600 27999 10652 28008
rect 10600 27965 10609 27999
rect 10609 27965 10643 27999
rect 10643 27965 10652 27999
rect 10600 27956 10652 27965
rect 20352 27956 20404 28008
rect 22008 27999 22060 28008
rect 8208 27888 8260 27940
rect 9036 27820 9088 27872
rect 11796 27863 11848 27872
rect 11796 27829 11805 27863
rect 11805 27829 11839 27863
rect 11839 27829 11848 27863
rect 11796 27820 11848 27829
rect 22008 27965 22017 27999
rect 22017 27965 22051 27999
rect 22051 27965 22060 27999
rect 22008 27956 22060 27965
rect 27620 27999 27672 28008
rect 27620 27965 27629 27999
rect 27629 27965 27663 27999
rect 27663 27965 27672 27999
rect 27620 27956 27672 27965
rect 28816 27999 28868 28008
rect 28816 27965 28825 27999
rect 28825 27965 28859 27999
rect 28859 27965 28868 27999
rect 28816 27956 28868 27965
rect 34520 27999 34572 28008
rect 34520 27965 34529 27999
rect 34529 27965 34563 27999
rect 34563 27965 34572 27999
rect 34520 27956 34572 27965
rect 39856 27956 39908 28008
rect 26240 27888 26292 27940
rect 31668 27888 31720 27940
rect 37096 27888 37148 27940
rect 37464 27888 37516 27940
rect 41420 27888 41472 27940
rect 42800 27956 42852 28008
rect 43260 28024 43312 28076
rect 43720 28024 43772 28076
rect 44088 28024 44140 28076
rect 44732 28024 44784 28076
rect 47768 28067 47820 28076
rect 47768 28033 47777 28067
rect 47777 28033 47811 28067
rect 47811 28033 47820 28067
rect 47768 28024 47820 28033
rect 43536 27956 43588 28008
rect 23940 27820 23992 27872
rect 25228 27863 25280 27872
rect 25228 27829 25237 27863
rect 25237 27829 25271 27863
rect 25271 27829 25280 27863
rect 25228 27820 25280 27829
rect 27160 27863 27212 27872
rect 27160 27829 27169 27863
rect 27169 27829 27203 27863
rect 27203 27829 27212 27863
rect 27160 27820 27212 27829
rect 33324 27820 33376 27872
rect 39028 27820 39080 27872
rect 42064 27820 42116 27872
rect 44364 27888 44416 27940
rect 42984 27820 43036 27872
rect 43904 27820 43956 27872
rect 46480 27820 46532 27872
rect 48136 27820 48188 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 12164 27659 12216 27668
rect 12164 27625 12173 27659
rect 12173 27625 12207 27659
rect 12207 27625 12216 27659
rect 12164 27616 12216 27625
rect 17408 27659 17460 27668
rect 17408 27625 17417 27659
rect 17417 27625 17451 27659
rect 17451 27625 17460 27659
rect 17408 27616 17460 27625
rect 7196 27591 7248 27600
rect 7196 27557 7205 27591
rect 7205 27557 7239 27591
rect 7239 27557 7248 27591
rect 7196 27548 7248 27557
rect 9220 27548 9272 27600
rect 10600 27591 10652 27600
rect 10600 27557 10609 27591
rect 10609 27557 10643 27591
rect 10643 27557 10652 27591
rect 10600 27548 10652 27557
rect 14832 27548 14884 27600
rect 17592 27548 17644 27600
rect 22376 27616 22428 27668
rect 25780 27616 25832 27668
rect 29920 27616 29972 27668
rect 38384 27659 38436 27668
rect 38384 27625 38393 27659
rect 38393 27625 38427 27659
rect 38427 27625 38436 27659
rect 38384 27616 38436 27625
rect 39120 27616 39172 27668
rect 40684 27616 40736 27668
rect 19432 27548 19484 27600
rect 22560 27548 22612 27600
rect 23020 27548 23072 27600
rect 25964 27548 26016 27600
rect 40316 27591 40368 27600
rect 40316 27557 40325 27591
rect 40325 27557 40359 27591
rect 40359 27557 40368 27591
rect 40316 27548 40368 27557
rect 7932 27523 7984 27532
rect 7932 27489 7941 27523
rect 7941 27489 7975 27523
rect 7975 27489 7984 27523
rect 7932 27480 7984 27489
rect 9956 27480 10008 27532
rect 12532 27480 12584 27532
rect 13728 27480 13780 27532
rect 15016 27480 15068 27532
rect 17224 27480 17276 27532
rect 18052 27480 18104 27532
rect 22008 27480 22060 27532
rect 6092 27387 6144 27396
rect 6092 27353 6126 27387
rect 6126 27353 6144 27387
rect 10232 27455 10284 27464
rect 10232 27421 10241 27455
rect 10241 27421 10275 27455
rect 10275 27421 10284 27455
rect 10232 27412 10284 27421
rect 14556 27412 14608 27464
rect 14832 27412 14884 27464
rect 17592 27455 17644 27464
rect 17592 27421 17601 27455
rect 17601 27421 17635 27455
rect 17635 27421 17644 27455
rect 17592 27412 17644 27421
rect 17776 27455 17828 27464
rect 17776 27421 17785 27455
rect 17785 27421 17819 27455
rect 17819 27421 17828 27455
rect 17776 27412 17828 27421
rect 22928 27412 22980 27464
rect 23020 27412 23072 27464
rect 23388 27412 23440 27464
rect 30012 27480 30064 27532
rect 43904 27616 43956 27668
rect 44088 27480 44140 27532
rect 28816 27412 28868 27464
rect 29644 27412 29696 27464
rect 30104 27412 30156 27464
rect 30380 27455 30432 27464
rect 30380 27421 30389 27455
rect 30389 27421 30423 27455
rect 30423 27421 30432 27455
rect 30380 27412 30432 27421
rect 32864 27455 32916 27464
rect 32864 27421 32873 27455
rect 32873 27421 32907 27455
rect 32907 27421 32916 27455
rect 32864 27412 32916 27421
rect 33140 27455 33192 27464
rect 33140 27421 33149 27455
rect 33149 27421 33183 27455
rect 33183 27421 33192 27455
rect 33140 27412 33192 27421
rect 36360 27455 36412 27464
rect 36360 27421 36369 27455
rect 36369 27421 36403 27455
rect 36403 27421 36412 27455
rect 36360 27412 36412 27421
rect 36544 27455 36596 27464
rect 36544 27421 36553 27455
rect 36553 27421 36587 27455
rect 36587 27421 36596 27455
rect 36544 27412 36596 27421
rect 38016 27455 38068 27464
rect 38016 27421 38025 27455
rect 38025 27421 38059 27455
rect 38059 27421 38068 27455
rect 38016 27412 38068 27421
rect 40224 27412 40276 27464
rect 41788 27455 41840 27464
rect 41788 27421 41797 27455
rect 41797 27421 41831 27455
rect 41831 27421 41840 27455
rect 41788 27412 41840 27421
rect 43352 27412 43404 27464
rect 44732 27616 44784 27668
rect 46848 27523 46900 27532
rect 46848 27489 46857 27523
rect 46857 27489 46891 27523
rect 46891 27489 46900 27523
rect 46848 27480 46900 27489
rect 48136 27523 48188 27532
rect 48136 27489 48145 27523
rect 48145 27489 48179 27523
rect 48179 27489 48188 27523
rect 48136 27480 48188 27489
rect 48320 27523 48372 27532
rect 48320 27489 48329 27523
rect 48329 27489 48363 27523
rect 48363 27489 48372 27523
rect 48320 27480 48372 27489
rect 44364 27412 44416 27464
rect 6092 27344 6144 27353
rect 8024 27344 8076 27396
rect 11796 27344 11848 27396
rect 15016 27344 15068 27396
rect 23756 27344 23808 27396
rect 25228 27344 25280 27396
rect 27160 27344 27212 27396
rect 41236 27344 41288 27396
rect 41512 27344 41564 27396
rect 43996 27344 44048 27396
rect 1860 27276 1912 27328
rect 12900 27276 12952 27328
rect 14372 27276 14424 27328
rect 27528 27276 27580 27328
rect 32680 27319 32732 27328
rect 32680 27285 32689 27319
rect 32689 27285 32723 27319
rect 32723 27285 32732 27319
rect 32680 27276 32732 27285
rect 39672 27276 39724 27328
rect 42800 27276 42852 27328
rect 47492 27276 47544 27328
rect 47676 27276 47728 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 6092 27072 6144 27124
rect 11796 27072 11848 27124
rect 17592 27072 17644 27124
rect 21180 27072 21232 27124
rect 25412 27072 25464 27124
rect 27804 27115 27856 27124
rect 7932 26936 7984 26988
rect 8024 26979 8076 26988
rect 8024 26945 8033 26979
rect 8033 26945 8067 26979
rect 8067 26945 8076 26979
rect 8024 26936 8076 26945
rect 9312 27004 9364 27056
rect 9036 26979 9088 26988
rect 9036 26945 9070 26979
rect 9070 26945 9088 26979
rect 9036 26936 9088 26945
rect 14372 26979 14424 26988
rect 14372 26945 14406 26979
rect 14406 26945 14424 26979
rect 14372 26936 14424 26945
rect 16212 26936 16264 26988
rect 18144 26936 18196 26988
rect 13636 26868 13688 26920
rect 17132 26911 17184 26920
rect 17132 26877 17141 26911
rect 17141 26877 17175 26911
rect 17175 26877 17184 26911
rect 17132 26868 17184 26877
rect 17868 26868 17920 26920
rect 24676 26936 24728 26988
rect 25964 26979 26016 26988
rect 20996 26868 21048 26920
rect 21364 26911 21416 26920
rect 21364 26877 21373 26911
rect 21373 26877 21407 26911
rect 21407 26877 21416 26911
rect 21364 26868 21416 26877
rect 25964 26945 25973 26979
rect 25973 26945 26007 26979
rect 26007 26945 26016 26979
rect 25964 26936 26016 26945
rect 27528 27004 27580 27056
rect 27804 27081 27813 27115
rect 27813 27081 27847 27115
rect 27847 27081 27856 27115
rect 27804 27072 27856 27081
rect 33140 27072 33192 27124
rect 36544 27072 36596 27124
rect 38016 27072 38068 27124
rect 32680 27004 32732 27056
rect 33416 27004 33468 27056
rect 34152 27004 34204 27056
rect 36360 27004 36412 27056
rect 26884 26868 26936 26920
rect 35440 26936 35492 26988
rect 36544 26936 36596 26988
rect 40224 27004 40276 27056
rect 38568 26936 38620 26988
rect 32036 26868 32088 26920
rect 36268 26911 36320 26920
rect 36268 26877 36277 26911
rect 36277 26877 36311 26911
rect 36311 26877 36320 26911
rect 36268 26868 36320 26877
rect 36452 26911 36504 26920
rect 36452 26877 36461 26911
rect 36461 26877 36495 26911
rect 36495 26877 36504 26911
rect 36452 26868 36504 26877
rect 37372 26868 37424 26920
rect 38844 26868 38896 26920
rect 39672 26911 39724 26920
rect 39672 26877 39681 26911
rect 39681 26877 39715 26911
rect 39715 26877 39724 26911
rect 41420 26979 41472 26988
rect 41420 26945 41429 26979
rect 41429 26945 41463 26979
rect 41463 26945 41472 26979
rect 41420 26936 41472 26945
rect 42892 26936 42944 26988
rect 43996 26936 44048 26988
rect 44180 26979 44232 26988
rect 44180 26945 44214 26979
rect 44214 26945 44232 26979
rect 44180 26936 44232 26945
rect 46756 26936 46808 26988
rect 47124 26936 47176 26988
rect 47400 26936 47452 26988
rect 47768 26979 47820 26988
rect 47768 26945 47777 26979
rect 47777 26945 47811 26979
rect 47811 26945 47820 26979
rect 47768 26936 47820 26945
rect 42064 26911 42116 26920
rect 39672 26868 39724 26877
rect 42064 26877 42073 26911
rect 42073 26877 42107 26911
rect 42107 26877 42116 26911
rect 42064 26868 42116 26877
rect 42984 26868 43036 26920
rect 10140 26775 10192 26784
rect 10140 26741 10149 26775
rect 10149 26741 10183 26775
rect 10183 26741 10192 26775
rect 10140 26732 10192 26741
rect 15200 26732 15252 26784
rect 20812 26732 20864 26784
rect 23572 26732 23624 26784
rect 24860 26732 24912 26784
rect 35348 26732 35400 26784
rect 35808 26775 35860 26784
rect 35808 26741 35817 26775
rect 35817 26741 35851 26775
rect 35851 26741 35860 26775
rect 35808 26732 35860 26741
rect 40500 26775 40552 26784
rect 40500 26741 40509 26775
rect 40509 26741 40543 26775
rect 40543 26741 40552 26775
rect 40500 26732 40552 26741
rect 45284 26775 45336 26784
rect 45284 26741 45293 26775
rect 45293 26741 45327 26775
rect 45327 26741 45336 26775
rect 45284 26732 45336 26741
rect 46664 26732 46716 26784
rect 48136 26732 48188 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 9956 26571 10008 26580
rect 9956 26537 9965 26571
rect 9965 26537 9999 26571
rect 9999 26537 10008 26571
rect 9956 26528 10008 26537
rect 14556 26571 14608 26580
rect 14556 26537 14565 26571
rect 14565 26537 14599 26571
rect 14599 26537 14608 26571
rect 14556 26528 14608 26537
rect 17776 26528 17828 26580
rect 10140 26392 10192 26444
rect 9588 26367 9640 26376
rect 9588 26333 9597 26367
rect 9597 26333 9631 26367
rect 9631 26333 9640 26367
rect 9588 26324 9640 26333
rect 12256 26367 12308 26376
rect 12256 26333 12265 26367
rect 12265 26333 12299 26367
rect 12299 26333 12308 26367
rect 12256 26324 12308 26333
rect 14556 26324 14608 26376
rect 14924 26324 14976 26376
rect 15200 26367 15252 26376
rect 15200 26333 15209 26367
rect 15209 26333 15243 26367
rect 15243 26333 15252 26367
rect 15200 26324 15252 26333
rect 16212 26324 16264 26376
rect 17776 26392 17828 26444
rect 18144 26392 18196 26444
rect 17132 26367 17184 26376
rect 17132 26333 17141 26367
rect 17141 26333 17175 26367
rect 17175 26333 17184 26367
rect 17132 26324 17184 26333
rect 17868 26324 17920 26376
rect 21364 26460 21416 26512
rect 23572 26528 23624 26580
rect 23756 26571 23808 26580
rect 23756 26537 23765 26571
rect 23765 26537 23799 26571
rect 23799 26537 23808 26571
rect 26240 26571 26292 26580
rect 23756 26528 23808 26537
rect 26240 26537 26249 26571
rect 26249 26537 26283 26571
rect 26283 26537 26292 26571
rect 26240 26528 26292 26537
rect 26976 26528 27028 26580
rect 33416 26571 33468 26580
rect 33416 26537 33425 26571
rect 33425 26537 33459 26571
rect 33459 26537 33468 26571
rect 33416 26528 33468 26537
rect 36268 26528 36320 26580
rect 22376 26392 22428 26444
rect 24032 26460 24084 26512
rect 20812 26367 20864 26376
rect 20812 26333 20821 26367
rect 20821 26333 20855 26367
rect 20855 26333 20864 26367
rect 20812 26324 20864 26333
rect 31944 26460 31996 26512
rect 32036 26435 32088 26444
rect 23940 26324 23992 26376
rect 25228 26367 25280 26376
rect 24676 26256 24728 26308
rect 25228 26333 25237 26367
rect 25237 26333 25271 26367
rect 25271 26333 25280 26367
rect 25228 26324 25280 26333
rect 26148 26324 26200 26376
rect 26884 26256 26936 26308
rect 12072 26231 12124 26240
rect 12072 26197 12081 26231
rect 12081 26197 12115 26231
rect 12115 26197 12124 26231
rect 12072 26188 12124 26197
rect 17040 26188 17092 26240
rect 19984 26231 20036 26240
rect 19984 26197 19993 26231
rect 19993 26197 20027 26231
rect 20027 26197 20036 26231
rect 19984 26188 20036 26197
rect 21456 26188 21508 26240
rect 23388 26231 23440 26240
rect 23388 26197 23397 26231
rect 23397 26197 23431 26231
rect 23431 26197 23440 26231
rect 23388 26188 23440 26197
rect 31116 26188 31168 26240
rect 32036 26401 32045 26435
rect 32045 26401 32079 26435
rect 32079 26401 32088 26435
rect 32036 26392 32088 26401
rect 44180 26571 44232 26580
rect 44180 26537 44189 26571
rect 44189 26537 44223 26571
rect 44223 26537 44232 26571
rect 44180 26528 44232 26537
rect 38384 26460 38436 26512
rect 34244 26324 34296 26376
rect 38016 26392 38068 26444
rect 38844 26324 38896 26376
rect 39672 26392 39724 26444
rect 40224 26392 40276 26444
rect 46480 26435 46532 26444
rect 46480 26401 46489 26435
rect 46489 26401 46523 26435
rect 46523 26401 46532 26435
rect 46480 26392 46532 26401
rect 46664 26435 46716 26444
rect 46664 26401 46673 26435
rect 46673 26401 46707 26435
rect 46707 26401 46716 26435
rect 46664 26392 46716 26401
rect 47952 26435 48004 26444
rect 47952 26401 47961 26435
rect 47961 26401 47995 26435
rect 47995 26401 48004 26435
rect 47952 26392 48004 26401
rect 40868 26324 40920 26376
rect 43996 26367 44048 26376
rect 43996 26333 44005 26367
rect 44005 26333 44039 26367
rect 44039 26333 44048 26367
rect 43996 26324 44048 26333
rect 32312 26299 32364 26308
rect 32312 26265 32346 26299
rect 32346 26265 32364 26299
rect 32312 26256 32364 26265
rect 35348 26256 35400 26308
rect 38568 26256 38620 26308
rect 40224 26256 40276 26308
rect 36360 26188 36412 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 7932 26027 7984 26036
rect 7932 25993 7941 26027
rect 7941 25993 7975 26027
rect 7975 25993 7984 26027
rect 7932 25984 7984 25993
rect 21456 26027 21508 26036
rect 21456 25993 21465 26027
rect 21465 25993 21499 26027
rect 21499 25993 21508 26027
rect 21456 25984 21508 25993
rect 22008 25984 22060 26036
rect 12072 25916 12124 25968
rect 18512 25916 18564 25968
rect 7104 25848 7156 25900
rect 17868 25848 17920 25900
rect 6460 25780 6512 25832
rect 3424 25644 3476 25696
rect 18144 25712 18196 25764
rect 18880 25848 18932 25900
rect 19984 25916 20036 25968
rect 23388 25916 23440 25968
rect 19524 25755 19576 25764
rect 19524 25721 19533 25755
rect 19533 25721 19567 25755
rect 19567 25721 19576 25755
rect 19524 25712 19576 25721
rect 12440 25644 12492 25696
rect 13084 25687 13136 25696
rect 13084 25653 13093 25687
rect 13093 25653 13127 25687
rect 13127 25653 13136 25687
rect 13084 25644 13136 25653
rect 18604 25644 18656 25696
rect 19616 25687 19668 25696
rect 19616 25653 19625 25687
rect 19625 25653 19659 25687
rect 19659 25653 19668 25687
rect 19616 25644 19668 25653
rect 25228 25984 25280 26036
rect 21640 25780 21692 25832
rect 24952 25848 25004 25900
rect 25688 25848 25740 25900
rect 26516 25916 26568 25968
rect 27160 25848 27212 25900
rect 31208 25848 31260 25900
rect 31668 25984 31720 26036
rect 32864 25984 32916 26036
rect 35440 26027 35492 26036
rect 35440 25993 35449 26027
rect 35449 25993 35483 26027
rect 35483 25993 35492 26027
rect 35440 25984 35492 25993
rect 35808 25984 35860 26036
rect 40500 25984 40552 26036
rect 43996 25984 44048 26036
rect 31760 25916 31812 25968
rect 40132 25916 40184 25968
rect 32588 25891 32640 25900
rect 25596 25823 25648 25832
rect 25596 25789 25605 25823
rect 25605 25789 25639 25823
rect 25639 25789 25648 25823
rect 25596 25780 25648 25789
rect 31116 25780 31168 25832
rect 31576 25780 31628 25832
rect 32588 25857 32597 25891
rect 32597 25857 32631 25891
rect 32631 25857 32640 25891
rect 32588 25848 32640 25857
rect 32864 25891 32916 25900
rect 32864 25857 32873 25891
rect 32873 25857 32907 25891
rect 32907 25857 32916 25891
rect 32864 25848 32916 25857
rect 33140 25848 33192 25900
rect 34796 25848 34848 25900
rect 36360 25848 36412 25900
rect 38016 25891 38068 25900
rect 38016 25857 38025 25891
rect 38025 25857 38059 25891
rect 38059 25857 38068 25891
rect 38016 25848 38068 25857
rect 38844 25891 38896 25900
rect 32680 25780 32732 25832
rect 34244 25780 34296 25832
rect 36636 25780 36688 25832
rect 37188 25780 37240 25832
rect 38844 25857 38853 25891
rect 38853 25857 38887 25891
rect 38887 25857 38896 25891
rect 38844 25848 38896 25857
rect 39028 25891 39080 25900
rect 39028 25857 39037 25891
rect 39037 25857 39071 25891
rect 39071 25857 39080 25891
rect 39028 25848 39080 25857
rect 38384 25780 38436 25832
rect 38568 25712 38620 25764
rect 38660 25712 38712 25764
rect 40316 25891 40368 25900
rect 40316 25857 40325 25891
rect 40325 25857 40359 25891
rect 40359 25857 40368 25891
rect 40316 25848 40368 25857
rect 45192 25848 45244 25900
rect 40224 25780 40276 25832
rect 43076 25780 43128 25832
rect 43996 25780 44048 25832
rect 44456 25823 44508 25832
rect 44456 25789 44465 25823
rect 44465 25789 44499 25823
rect 44499 25789 44508 25823
rect 44456 25780 44508 25789
rect 45284 25780 45336 25832
rect 46756 25823 46808 25832
rect 46756 25789 46765 25823
rect 46765 25789 46799 25823
rect 46799 25789 46808 25823
rect 46756 25780 46808 25789
rect 47032 25823 47084 25832
rect 47032 25789 47041 25823
rect 47041 25789 47075 25823
rect 47075 25789 47084 25823
rect 47032 25780 47084 25789
rect 47216 25823 47268 25832
rect 47216 25789 47225 25823
rect 47225 25789 47259 25823
rect 47259 25789 47268 25823
rect 47216 25780 47268 25789
rect 20352 25644 20404 25696
rect 26424 25687 26476 25696
rect 26424 25653 26433 25687
rect 26433 25653 26467 25687
rect 26467 25653 26476 25687
rect 26424 25644 26476 25653
rect 29552 25687 29604 25696
rect 29552 25653 29561 25687
rect 29561 25653 29595 25687
rect 29595 25653 29604 25687
rect 29552 25644 29604 25653
rect 30196 25644 30248 25696
rect 33692 25644 33744 25696
rect 38292 25644 38344 25696
rect 48320 25644 48372 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 6460 25483 6512 25492
rect 6460 25449 6469 25483
rect 6469 25449 6503 25483
rect 6503 25449 6512 25483
rect 6460 25440 6512 25449
rect 7104 25483 7156 25492
rect 7104 25449 7113 25483
rect 7113 25449 7147 25483
rect 7147 25449 7156 25483
rect 7104 25440 7156 25449
rect 12256 25440 12308 25492
rect 18604 25483 18656 25492
rect 18604 25449 18613 25483
rect 18613 25449 18647 25483
rect 18647 25449 18656 25483
rect 18604 25440 18656 25449
rect 19524 25440 19576 25492
rect 24952 25483 25004 25492
rect 24952 25449 24961 25483
rect 24961 25449 24995 25483
rect 24995 25449 25004 25483
rect 24952 25440 25004 25449
rect 29644 25440 29696 25492
rect 31208 25483 31260 25492
rect 31208 25449 31217 25483
rect 31217 25449 31251 25483
rect 31251 25449 31260 25483
rect 31208 25440 31260 25449
rect 32312 25440 32364 25492
rect 32588 25440 32640 25492
rect 33784 25440 33836 25492
rect 43076 25483 43128 25492
rect 43076 25449 43085 25483
rect 43085 25449 43119 25483
rect 43119 25449 43128 25483
rect 43076 25440 43128 25449
rect 43536 25440 43588 25492
rect 44456 25440 44508 25492
rect 45192 25483 45244 25492
rect 45192 25449 45201 25483
rect 45201 25449 45235 25483
rect 45235 25449 45244 25483
rect 45192 25440 45244 25449
rect 9312 25372 9364 25424
rect 18512 25415 18564 25424
rect 3424 25347 3476 25356
rect 3424 25313 3433 25347
rect 3433 25313 3467 25347
rect 3467 25313 3476 25347
rect 3424 25304 3476 25313
rect 8024 25304 8076 25356
rect 9588 25347 9640 25356
rect 1584 25279 1636 25288
rect 1584 25245 1593 25279
rect 1593 25245 1627 25279
rect 1627 25245 1636 25279
rect 1584 25236 1636 25245
rect 9588 25313 9597 25347
rect 9597 25313 9631 25347
rect 9631 25313 9640 25347
rect 9588 25304 9640 25313
rect 18512 25381 18521 25415
rect 18521 25381 18555 25415
rect 18555 25381 18564 25415
rect 18512 25372 18564 25381
rect 12532 25304 12584 25356
rect 17040 25347 17092 25356
rect 17040 25313 17049 25347
rect 17049 25313 17083 25347
rect 17083 25313 17092 25347
rect 17040 25304 17092 25313
rect 20996 25415 21048 25424
rect 20996 25381 21005 25415
rect 21005 25381 21039 25415
rect 21039 25381 21048 25415
rect 20996 25372 21048 25381
rect 3240 25211 3292 25220
rect 3240 25177 3249 25211
rect 3249 25177 3283 25211
rect 3283 25177 3292 25211
rect 3240 25168 3292 25177
rect 8024 25168 8076 25220
rect 13084 25236 13136 25288
rect 15292 25236 15344 25288
rect 15936 25279 15988 25288
rect 15936 25245 15945 25279
rect 15945 25245 15979 25279
rect 15979 25245 15988 25279
rect 15936 25236 15988 25245
rect 16212 25279 16264 25288
rect 16212 25245 16221 25279
rect 16221 25245 16255 25279
rect 16255 25245 16264 25279
rect 16212 25236 16264 25245
rect 16948 25236 17000 25288
rect 17868 25236 17920 25288
rect 19616 25304 19668 25356
rect 23848 25304 23900 25356
rect 18880 25279 18932 25288
rect 18880 25245 18889 25279
rect 18889 25245 18923 25279
rect 18923 25245 18932 25279
rect 20628 25279 20680 25288
rect 18880 25236 18932 25245
rect 20628 25245 20637 25279
rect 20637 25245 20671 25279
rect 20671 25245 20680 25279
rect 20628 25236 20680 25245
rect 21456 25279 21508 25288
rect 21456 25245 21465 25279
rect 21465 25245 21499 25279
rect 21499 25245 21508 25279
rect 21456 25236 21508 25245
rect 21640 25279 21692 25288
rect 21640 25245 21649 25279
rect 21649 25245 21683 25279
rect 21683 25245 21692 25279
rect 21640 25236 21692 25245
rect 23664 25279 23716 25288
rect 23664 25245 23673 25279
rect 23673 25245 23707 25279
rect 23707 25245 23716 25279
rect 23664 25236 23716 25245
rect 8576 25211 8628 25220
rect 8576 25177 8585 25211
rect 8585 25177 8619 25211
rect 8619 25177 8628 25211
rect 8576 25168 8628 25177
rect 11612 25211 11664 25220
rect 11612 25177 11621 25211
rect 11621 25177 11655 25211
rect 11655 25177 11664 25211
rect 11612 25168 11664 25177
rect 16120 25211 16172 25220
rect 16120 25177 16129 25211
rect 16129 25177 16163 25211
rect 16163 25177 16172 25211
rect 16120 25168 16172 25177
rect 18236 25168 18288 25220
rect 25596 25304 25648 25356
rect 24124 25236 24176 25288
rect 26424 25236 26476 25288
rect 12624 25100 12676 25152
rect 14832 25143 14884 25152
rect 14832 25109 14841 25143
rect 14841 25109 14875 25143
rect 14875 25109 14884 25143
rect 14832 25100 14884 25109
rect 17316 25100 17368 25152
rect 17500 25143 17552 25152
rect 17500 25109 17509 25143
rect 17509 25109 17543 25143
rect 17543 25109 17552 25143
rect 17500 25100 17552 25109
rect 18144 25143 18196 25152
rect 18144 25109 18153 25143
rect 18153 25109 18187 25143
rect 18187 25109 18196 25143
rect 18144 25100 18196 25109
rect 23756 25100 23808 25152
rect 25872 25168 25924 25220
rect 29552 25236 29604 25288
rect 38384 25372 38436 25424
rect 41788 25372 41840 25424
rect 43352 25372 43404 25424
rect 30288 25279 30340 25288
rect 30288 25245 30297 25279
rect 30297 25245 30331 25279
rect 30331 25245 30340 25279
rect 30288 25236 30340 25245
rect 26240 25100 26292 25152
rect 27344 25100 27396 25152
rect 30196 25168 30248 25220
rect 30472 25100 30524 25152
rect 30564 25100 30616 25152
rect 31576 25279 31628 25288
rect 31576 25245 31585 25279
rect 31585 25245 31619 25279
rect 31619 25245 31628 25279
rect 31576 25236 31628 25245
rect 32680 25279 32732 25288
rect 32680 25245 32689 25279
rect 32689 25245 32723 25279
rect 32723 25245 32732 25279
rect 33692 25279 33744 25288
rect 32680 25236 32732 25245
rect 33692 25245 33701 25279
rect 33701 25245 33735 25279
rect 33735 25245 33744 25279
rect 33692 25236 33744 25245
rect 33968 25279 34020 25288
rect 33968 25245 33977 25279
rect 33977 25245 34011 25279
rect 34011 25245 34020 25279
rect 33968 25236 34020 25245
rect 34152 25279 34204 25288
rect 34152 25245 34161 25279
rect 34161 25245 34195 25279
rect 34195 25245 34204 25279
rect 34152 25236 34204 25245
rect 40132 25279 40184 25288
rect 40132 25245 40141 25279
rect 40141 25245 40175 25279
rect 40175 25245 40184 25279
rect 40132 25236 40184 25245
rect 42340 25279 42392 25288
rect 42340 25245 42349 25279
rect 42349 25245 42383 25279
rect 42383 25245 42392 25279
rect 42340 25236 42392 25245
rect 40868 25211 40920 25220
rect 40868 25177 40877 25211
rect 40877 25177 40911 25211
rect 40911 25177 40920 25211
rect 40868 25168 40920 25177
rect 42064 25211 42116 25220
rect 42064 25177 42073 25211
rect 42073 25177 42107 25211
rect 42107 25177 42116 25211
rect 42064 25168 42116 25177
rect 46848 25347 46900 25356
rect 46848 25313 46857 25347
rect 46857 25313 46891 25347
rect 46891 25313 46900 25347
rect 46848 25304 46900 25313
rect 48136 25347 48188 25356
rect 48136 25313 48145 25347
rect 48145 25313 48179 25347
rect 48179 25313 48188 25347
rect 48136 25304 48188 25313
rect 48320 25347 48372 25356
rect 48320 25313 48329 25347
rect 48329 25313 48363 25347
rect 48363 25313 48372 25347
rect 48320 25304 48372 25313
rect 42892 25236 42944 25288
rect 43444 25279 43496 25288
rect 43444 25245 43453 25279
rect 43453 25245 43487 25279
rect 43487 25245 43496 25279
rect 43444 25236 43496 25245
rect 39488 25100 39540 25152
rect 41420 25100 41472 25152
rect 41972 25100 42024 25152
rect 45560 25211 45612 25220
rect 45560 25177 45569 25211
rect 45569 25177 45603 25211
rect 45603 25177 45612 25211
rect 45560 25168 45612 25177
rect 43076 25100 43128 25152
rect 43444 25100 43496 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 9588 24896 9640 24948
rect 11612 24896 11664 24948
rect 13544 24896 13596 24948
rect 2596 24803 2648 24812
rect 2596 24769 2605 24803
rect 2605 24769 2639 24803
rect 2639 24769 2648 24803
rect 2596 24760 2648 24769
rect 5264 24760 5316 24812
rect 8024 24760 8076 24812
rect 8852 24760 8904 24812
rect 10232 24803 10284 24812
rect 10232 24769 10241 24803
rect 10241 24769 10275 24803
rect 10275 24769 10284 24803
rect 10232 24760 10284 24769
rect 3240 24692 3292 24744
rect 9312 24692 9364 24744
rect 11152 24556 11204 24608
rect 12440 24828 12492 24880
rect 11796 24760 11848 24812
rect 12992 24760 13044 24812
rect 16120 24896 16172 24948
rect 17868 24939 17920 24948
rect 14832 24828 14884 24880
rect 17868 24905 17877 24939
rect 17877 24905 17911 24939
rect 17911 24905 17920 24939
rect 17868 24896 17920 24905
rect 20628 24896 20680 24948
rect 27344 24939 27396 24948
rect 27344 24905 27353 24939
rect 27353 24905 27387 24939
rect 27387 24905 27396 24939
rect 27344 24896 27396 24905
rect 30288 24896 30340 24948
rect 24860 24828 24912 24880
rect 17684 24803 17736 24812
rect 13636 24692 13688 24744
rect 16488 24692 16540 24744
rect 17684 24769 17693 24803
rect 17693 24769 17727 24803
rect 17727 24769 17736 24803
rect 17684 24760 17736 24769
rect 17316 24624 17368 24676
rect 19616 24760 19668 24812
rect 19064 24692 19116 24744
rect 23480 24760 23532 24812
rect 23572 24760 23624 24812
rect 25872 24803 25924 24812
rect 25872 24769 25881 24803
rect 25881 24769 25915 24803
rect 25915 24769 25924 24803
rect 25872 24760 25924 24769
rect 26240 24803 26292 24812
rect 26240 24769 26249 24803
rect 26249 24769 26283 24803
rect 26283 24769 26292 24803
rect 26240 24760 26292 24769
rect 19984 24735 20036 24744
rect 19984 24701 19993 24735
rect 19993 24701 20027 24735
rect 20027 24701 20036 24735
rect 23112 24735 23164 24744
rect 19984 24692 20036 24701
rect 12348 24556 12400 24608
rect 13912 24599 13964 24608
rect 13912 24565 13921 24599
rect 13921 24565 13955 24599
rect 13955 24565 13964 24599
rect 13912 24556 13964 24565
rect 17868 24556 17920 24608
rect 19340 24556 19392 24608
rect 20444 24556 20496 24608
rect 22008 24556 22060 24608
rect 23112 24701 23121 24735
rect 23121 24701 23155 24735
rect 23155 24701 23164 24735
rect 23112 24692 23164 24701
rect 23848 24692 23900 24744
rect 26148 24624 26200 24676
rect 27436 24803 27488 24812
rect 27436 24769 27445 24803
rect 27445 24769 27479 24803
rect 27479 24769 27488 24803
rect 27436 24760 27488 24769
rect 30748 24803 30800 24812
rect 27160 24667 27212 24676
rect 27160 24633 27169 24667
rect 27169 24633 27203 24667
rect 27203 24633 27212 24667
rect 27160 24624 27212 24633
rect 29000 24667 29052 24676
rect 29000 24633 29009 24667
rect 29009 24633 29043 24667
rect 29043 24633 29052 24667
rect 29000 24624 29052 24633
rect 30748 24769 30757 24803
rect 30757 24769 30791 24803
rect 30791 24769 30800 24803
rect 30748 24760 30800 24769
rect 31024 24760 31076 24812
rect 31208 24803 31260 24812
rect 31208 24769 31217 24803
rect 31217 24769 31251 24803
rect 31251 24769 31260 24803
rect 31208 24760 31260 24769
rect 32772 24896 32824 24948
rect 36452 24896 36504 24948
rect 41972 24939 42024 24948
rect 41972 24905 41981 24939
rect 41981 24905 42015 24939
rect 42015 24905 42024 24939
rect 41972 24896 42024 24905
rect 45560 24896 45612 24948
rect 33508 24828 33560 24880
rect 33968 24828 34020 24880
rect 31484 24760 31536 24812
rect 30472 24692 30524 24744
rect 32864 24760 32916 24812
rect 33600 24803 33652 24812
rect 33600 24769 33609 24803
rect 33609 24769 33643 24803
rect 33643 24769 33652 24803
rect 33600 24760 33652 24769
rect 33784 24803 33836 24812
rect 33784 24769 33793 24803
rect 33793 24769 33827 24803
rect 33827 24769 33836 24803
rect 33784 24760 33836 24769
rect 37740 24760 37792 24812
rect 34152 24692 34204 24744
rect 38660 24760 38712 24812
rect 38844 24760 38896 24812
rect 38108 24692 38160 24744
rect 38568 24692 38620 24744
rect 41788 24803 41840 24812
rect 41788 24769 41797 24803
rect 41797 24769 41831 24803
rect 41831 24769 41840 24803
rect 41788 24760 41840 24769
rect 43536 24828 43588 24880
rect 43168 24803 43220 24812
rect 43168 24769 43176 24803
rect 43176 24769 43210 24803
rect 43210 24769 43220 24803
rect 43168 24760 43220 24769
rect 43444 24760 43496 24812
rect 44548 24803 44600 24812
rect 44548 24769 44582 24803
rect 44582 24769 44600 24803
rect 44548 24760 44600 24769
rect 42892 24692 42944 24744
rect 43076 24735 43128 24744
rect 43076 24701 43085 24735
rect 43085 24701 43119 24735
rect 43119 24701 43128 24735
rect 43076 24692 43128 24701
rect 43260 24735 43312 24744
rect 43260 24701 43269 24735
rect 43269 24701 43303 24735
rect 43303 24701 43312 24735
rect 43260 24692 43312 24701
rect 43352 24735 43404 24744
rect 43352 24701 43361 24735
rect 43361 24701 43395 24735
rect 43395 24701 43404 24735
rect 47032 24760 47084 24812
rect 47216 24803 47268 24812
rect 47216 24769 47225 24803
rect 47225 24769 47259 24803
rect 47259 24769 47268 24803
rect 47216 24760 47268 24769
rect 48228 24803 48280 24812
rect 48228 24769 48237 24803
rect 48237 24769 48271 24803
rect 48271 24769 48280 24803
rect 48228 24760 48280 24769
rect 43352 24692 43404 24701
rect 47492 24692 47544 24744
rect 31760 24556 31812 24608
rect 31852 24556 31904 24608
rect 33232 24556 33284 24608
rect 34152 24556 34204 24608
rect 34704 24556 34756 24608
rect 36452 24556 36504 24608
rect 37832 24556 37884 24608
rect 38660 24556 38712 24608
rect 39212 24599 39264 24608
rect 39212 24565 39221 24599
rect 39221 24565 39255 24599
rect 39255 24565 39264 24599
rect 39212 24556 39264 24565
rect 41604 24599 41656 24608
rect 41604 24565 41613 24599
rect 41613 24565 41647 24599
rect 41647 24565 41656 24599
rect 41604 24556 41656 24565
rect 42708 24556 42760 24608
rect 43444 24556 43496 24608
rect 44180 24556 44232 24608
rect 47216 24624 47268 24676
rect 48044 24667 48096 24676
rect 48044 24633 48053 24667
rect 48053 24633 48087 24667
rect 48087 24633 48096 24667
rect 48044 24624 48096 24633
rect 45560 24556 45612 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 11796 24395 11848 24404
rect 11796 24361 11805 24395
rect 11805 24361 11839 24395
rect 11839 24361 11848 24395
rect 11796 24352 11848 24361
rect 12992 24395 13044 24404
rect 12992 24361 13001 24395
rect 13001 24361 13035 24395
rect 13035 24361 13044 24395
rect 12992 24352 13044 24361
rect 16672 24352 16724 24404
rect 17684 24352 17736 24404
rect 19616 24395 19668 24404
rect 19616 24361 19625 24395
rect 19625 24361 19659 24395
rect 19659 24361 19668 24395
rect 19616 24352 19668 24361
rect 20076 24352 20128 24404
rect 23020 24352 23072 24404
rect 26148 24352 26200 24404
rect 27436 24352 27488 24404
rect 8576 24216 8628 24268
rect 8208 24191 8260 24200
rect 8208 24157 8217 24191
rect 8217 24157 8251 24191
rect 8251 24157 8260 24191
rect 14556 24284 14608 24336
rect 12440 24259 12492 24268
rect 12440 24225 12449 24259
rect 12449 24225 12483 24259
rect 12483 24225 12492 24259
rect 12440 24216 12492 24225
rect 14740 24216 14792 24268
rect 15384 24284 15436 24336
rect 15936 24284 15988 24336
rect 16488 24284 16540 24336
rect 11152 24191 11204 24200
rect 8208 24148 8260 24157
rect 11152 24157 11161 24191
rect 11161 24157 11195 24191
rect 11195 24157 11204 24191
rect 11152 24148 11204 24157
rect 13912 24148 13964 24200
rect 14556 24191 14608 24200
rect 14556 24157 14565 24191
rect 14565 24157 14599 24191
rect 14599 24157 14608 24191
rect 14556 24148 14608 24157
rect 14924 24148 14976 24200
rect 15384 24148 15436 24200
rect 3332 24080 3384 24132
rect 6644 24080 6696 24132
rect 10140 24012 10192 24064
rect 12348 24080 12400 24132
rect 15292 24080 15344 24132
rect 14464 24012 14516 24064
rect 16396 24216 16448 24268
rect 16120 24148 16172 24200
rect 16948 24284 17000 24336
rect 17500 24216 17552 24268
rect 17592 24148 17644 24200
rect 21364 24216 21416 24268
rect 22008 24259 22060 24268
rect 22008 24225 22017 24259
rect 22017 24225 22051 24259
rect 22051 24225 22060 24259
rect 22008 24216 22060 24225
rect 22836 24259 22888 24268
rect 22836 24225 22845 24259
rect 22845 24225 22879 24259
rect 22879 24225 22888 24259
rect 22836 24216 22888 24225
rect 19800 24191 19852 24200
rect 19800 24157 19809 24191
rect 19809 24157 19843 24191
rect 19843 24157 19852 24191
rect 19800 24148 19852 24157
rect 20076 24191 20128 24200
rect 20076 24157 20085 24191
rect 20085 24157 20119 24191
rect 20119 24157 20128 24191
rect 20076 24148 20128 24157
rect 17132 24012 17184 24064
rect 25872 24148 25924 24200
rect 20628 24080 20680 24132
rect 27620 24216 27672 24268
rect 26792 24191 26844 24200
rect 26792 24157 26801 24191
rect 26801 24157 26835 24191
rect 26835 24157 26844 24191
rect 26792 24148 26844 24157
rect 19800 24012 19852 24064
rect 20168 24012 20220 24064
rect 20260 24012 20312 24064
rect 26056 24012 26108 24064
rect 26700 24055 26752 24064
rect 26700 24021 26709 24055
rect 26709 24021 26743 24055
rect 26743 24021 26752 24055
rect 26700 24012 26752 24021
rect 27620 24080 27672 24132
rect 28540 24191 28592 24200
rect 28540 24157 28549 24191
rect 28549 24157 28583 24191
rect 28583 24157 28592 24191
rect 28540 24148 28592 24157
rect 29000 24352 29052 24404
rect 32496 24352 32548 24404
rect 31208 24284 31260 24336
rect 31760 24284 31812 24336
rect 34520 24352 34572 24404
rect 38108 24395 38160 24404
rect 38108 24361 38117 24395
rect 38117 24361 38151 24395
rect 38151 24361 38160 24395
rect 38108 24352 38160 24361
rect 42064 24352 42116 24404
rect 43536 24395 43588 24404
rect 31116 24216 31168 24268
rect 28448 24080 28500 24132
rect 31484 24148 31536 24200
rect 33968 24216 34020 24268
rect 43536 24361 43545 24395
rect 43545 24361 43579 24395
rect 43579 24361 43588 24395
rect 43536 24352 43588 24361
rect 43168 24259 43220 24268
rect 30472 24080 30524 24132
rect 34244 24148 34296 24200
rect 43168 24225 43177 24259
rect 43177 24225 43211 24259
rect 43211 24225 43220 24259
rect 43168 24216 43220 24225
rect 43996 24259 44048 24268
rect 43996 24225 44005 24259
rect 44005 24225 44039 24259
rect 44039 24225 44048 24259
rect 43996 24216 44048 24225
rect 48136 24259 48188 24268
rect 48136 24225 48145 24259
rect 48145 24225 48179 24259
rect 48179 24225 48188 24259
rect 48136 24216 48188 24225
rect 31852 24123 31904 24132
rect 31852 24089 31861 24123
rect 31861 24089 31895 24123
rect 31895 24089 31904 24123
rect 31852 24080 31904 24089
rect 33140 24123 33192 24132
rect 33140 24089 33174 24123
rect 33174 24089 33192 24123
rect 33140 24080 33192 24089
rect 33784 24012 33836 24064
rect 34888 24012 34940 24064
rect 36176 24080 36228 24132
rect 38936 24148 38988 24200
rect 40868 24148 40920 24200
rect 42708 24148 42760 24200
rect 43352 24191 43404 24200
rect 43352 24157 43361 24191
rect 43361 24157 43395 24191
rect 43395 24157 43404 24191
rect 43352 24148 43404 24157
rect 44180 24191 44232 24200
rect 44180 24157 44189 24191
rect 44189 24157 44223 24191
rect 44223 24157 44232 24191
rect 44180 24148 44232 24157
rect 46480 24191 46532 24200
rect 46480 24157 46489 24191
rect 46489 24157 46523 24191
rect 46523 24157 46532 24191
rect 46480 24148 46532 24157
rect 36728 24012 36780 24064
rect 39120 24080 39172 24132
rect 39212 24123 39264 24132
rect 39212 24089 39230 24123
rect 39230 24089 39264 24123
rect 41604 24123 41656 24132
rect 39212 24080 39264 24089
rect 41604 24089 41638 24123
rect 41638 24089 41656 24123
rect 41604 24080 41656 24089
rect 42340 24080 42392 24132
rect 47860 24080 47912 24132
rect 42800 24012 42852 24064
rect 44272 24012 44324 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 6644 23851 6696 23860
rect 6644 23817 6653 23851
rect 6653 23817 6687 23851
rect 6687 23817 6696 23851
rect 6644 23808 6696 23817
rect 8852 23851 8904 23860
rect 8852 23817 8861 23851
rect 8861 23817 8895 23851
rect 8895 23817 8904 23851
rect 8852 23808 8904 23817
rect 10140 23851 10192 23860
rect 6552 23715 6604 23724
rect 6552 23681 6561 23715
rect 6561 23681 6595 23715
rect 6595 23681 6604 23715
rect 6552 23672 6604 23681
rect 10140 23817 10149 23851
rect 10149 23817 10183 23851
rect 10183 23817 10192 23851
rect 10140 23808 10192 23817
rect 15384 23851 15436 23860
rect 15384 23817 15393 23851
rect 15393 23817 15427 23851
rect 15427 23817 15436 23851
rect 15384 23808 15436 23817
rect 17132 23808 17184 23860
rect 20260 23808 20312 23860
rect 20628 23851 20680 23860
rect 20628 23817 20637 23851
rect 20637 23817 20671 23851
rect 20671 23817 20680 23851
rect 20628 23808 20680 23817
rect 23112 23808 23164 23860
rect 23572 23851 23624 23860
rect 23572 23817 23581 23851
rect 23581 23817 23615 23851
rect 23615 23817 23624 23851
rect 23572 23808 23624 23817
rect 23664 23808 23716 23860
rect 26332 23808 26384 23860
rect 11704 23672 11756 23724
rect 14280 23715 14332 23724
rect 14280 23681 14314 23715
rect 14314 23681 14332 23715
rect 20352 23740 20404 23792
rect 14280 23672 14332 23681
rect 19340 23672 19392 23724
rect 23204 23715 23256 23724
rect 9312 23604 9364 23656
rect 13084 23604 13136 23656
rect 13636 23604 13688 23656
rect 23204 23681 23213 23715
rect 23213 23681 23247 23715
rect 23247 23681 23256 23715
rect 23204 23672 23256 23681
rect 25504 23604 25556 23656
rect 28448 23808 28500 23860
rect 27712 23715 27764 23724
rect 27712 23681 27721 23715
rect 27721 23681 27755 23715
rect 27755 23681 27764 23715
rect 27712 23672 27764 23681
rect 27160 23604 27212 23656
rect 27620 23604 27672 23656
rect 23480 23536 23532 23588
rect 30748 23740 30800 23792
rect 32496 23808 32548 23860
rect 33048 23808 33100 23860
rect 36176 23808 36228 23860
rect 38844 23851 38896 23860
rect 38844 23817 38853 23851
rect 38853 23817 38887 23851
rect 38887 23817 38896 23851
rect 38844 23808 38896 23817
rect 39028 23808 39080 23860
rect 43628 23808 43680 23860
rect 44548 23808 44600 23860
rect 47860 23851 47912 23860
rect 47860 23817 47869 23851
rect 47869 23817 47903 23851
rect 47903 23817 47912 23851
rect 47860 23808 47912 23817
rect 47124 23740 47176 23792
rect 30380 23715 30432 23724
rect 30380 23681 30389 23715
rect 30389 23681 30423 23715
rect 30423 23681 30432 23715
rect 30380 23672 30432 23681
rect 30472 23672 30524 23724
rect 31116 23604 31168 23656
rect 33508 23672 33560 23724
rect 33784 23715 33836 23724
rect 33784 23681 33793 23715
rect 33793 23681 33827 23715
rect 33827 23681 33836 23715
rect 33784 23672 33836 23681
rect 34244 23715 34296 23724
rect 34244 23681 34253 23715
rect 34253 23681 34287 23715
rect 34287 23681 34296 23715
rect 34244 23672 34296 23681
rect 34796 23672 34848 23724
rect 34888 23672 34940 23724
rect 36636 23715 36688 23724
rect 36636 23681 36645 23715
rect 36645 23681 36679 23715
rect 36679 23681 36688 23715
rect 36636 23672 36688 23681
rect 37648 23672 37700 23724
rect 37740 23672 37792 23724
rect 39120 23672 39172 23724
rect 39488 23715 39540 23724
rect 33692 23604 33744 23656
rect 36452 23647 36504 23656
rect 36452 23613 36461 23647
rect 36461 23613 36495 23647
rect 36495 23613 36504 23647
rect 36452 23604 36504 23613
rect 36728 23604 36780 23656
rect 39488 23681 39497 23715
rect 39497 23681 39531 23715
rect 39531 23681 39540 23715
rect 39488 23672 39540 23681
rect 43260 23672 43312 23724
rect 44272 23715 44324 23724
rect 44272 23681 44281 23715
rect 44281 23681 44315 23715
rect 44315 23681 44324 23715
rect 44272 23672 44324 23681
rect 46480 23672 46532 23724
rect 39396 23604 39448 23656
rect 30288 23536 30340 23588
rect 20536 23468 20588 23520
rect 26608 23468 26660 23520
rect 27804 23468 27856 23520
rect 29276 23468 29328 23520
rect 31668 23511 31720 23520
rect 31668 23477 31677 23511
rect 31677 23477 31711 23511
rect 31711 23477 31720 23511
rect 31668 23468 31720 23477
rect 33232 23468 33284 23520
rect 39028 23536 39080 23588
rect 35624 23511 35676 23520
rect 35624 23477 35633 23511
rect 35633 23477 35667 23511
rect 35667 23477 35676 23511
rect 35624 23468 35676 23477
rect 36084 23468 36136 23520
rect 36636 23468 36688 23520
rect 40408 23511 40460 23520
rect 40408 23477 40417 23511
rect 40417 23477 40451 23511
rect 40451 23477 40460 23511
rect 40408 23468 40460 23477
rect 42800 23468 42852 23520
rect 42984 23468 43036 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 14280 23307 14332 23316
rect 14280 23273 14289 23307
rect 14289 23273 14323 23307
rect 14323 23273 14332 23307
rect 14280 23264 14332 23273
rect 21272 23264 21324 23316
rect 14648 23196 14700 23248
rect 26700 23264 26752 23316
rect 32588 23264 32640 23316
rect 33140 23264 33192 23316
rect 34796 23264 34848 23316
rect 37648 23307 37700 23316
rect 37648 23273 37657 23307
rect 37657 23273 37691 23307
rect 37691 23273 37700 23307
rect 37648 23264 37700 23273
rect 42340 23307 42392 23316
rect 42340 23273 42349 23307
rect 42349 23273 42383 23307
rect 42383 23273 42392 23307
rect 42340 23264 42392 23273
rect 11704 23060 11756 23112
rect 12440 23128 12492 23180
rect 19984 23128 20036 23180
rect 22376 23171 22428 23180
rect 22376 23137 22385 23171
rect 22385 23137 22419 23171
rect 22419 23137 22428 23171
rect 22376 23128 22428 23137
rect 23204 23128 23256 23180
rect 26976 23128 27028 23180
rect 14464 23103 14516 23112
rect 14464 23069 14473 23103
rect 14473 23069 14507 23103
rect 14507 23069 14516 23103
rect 14464 23060 14516 23069
rect 14648 23103 14700 23112
rect 14648 23069 14657 23103
rect 14657 23069 14691 23103
rect 14691 23069 14700 23103
rect 14648 23060 14700 23069
rect 15016 23060 15068 23112
rect 24768 23103 24820 23112
rect 24768 23069 24777 23103
rect 24777 23069 24811 23103
rect 24811 23069 24820 23103
rect 24768 23060 24820 23069
rect 25044 23103 25096 23112
rect 25044 23069 25053 23103
rect 25053 23069 25087 23103
rect 25087 23069 25096 23103
rect 25044 23060 25096 23069
rect 11612 22924 11664 22976
rect 12808 22924 12860 22976
rect 16212 22924 16264 22976
rect 17592 22924 17644 22976
rect 22652 22924 22704 22976
rect 22744 22924 22796 22976
rect 24584 22967 24636 22976
rect 24584 22933 24593 22967
rect 24593 22933 24627 22967
rect 24627 22933 24636 22967
rect 24584 22924 24636 22933
rect 27344 23060 27396 23112
rect 26608 22992 26660 23044
rect 27712 23196 27764 23248
rect 29276 23196 29328 23248
rect 32220 23196 32272 23248
rect 48044 23264 48096 23316
rect 43260 23196 43312 23248
rect 30104 23128 30156 23180
rect 31576 23128 31628 23180
rect 33600 23128 33652 23180
rect 35624 23128 35676 23180
rect 27620 23103 27672 23112
rect 27620 23069 27629 23103
rect 27629 23069 27663 23103
rect 27663 23069 27672 23103
rect 27620 23060 27672 23069
rect 28448 23103 28500 23112
rect 27804 23035 27856 23044
rect 27804 23001 27813 23035
rect 27813 23001 27847 23035
rect 27847 23001 27856 23035
rect 27804 22992 27856 23001
rect 28448 23069 28457 23103
rect 28457 23069 28491 23103
rect 28491 23069 28500 23103
rect 28448 23060 28500 23069
rect 28540 23060 28592 23112
rect 30288 23103 30340 23112
rect 30288 23069 30297 23103
rect 30297 23069 30331 23103
rect 30331 23069 30340 23103
rect 30288 23060 30340 23069
rect 30472 23103 30524 23112
rect 30472 23069 30481 23103
rect 30481 23069 30515 23103
rect 30515 23069 30524 23103
rect 30472 23060 30524 23069
rect 31668 23060 31720 23112
rect 33232 23103 33284 23112
rect 33232 23069 33241 23103
rect 33241 23069 33275 23103
rect 33275 23069 33284 23103
rect 33232 23060 33284 23069
rect 34704 23060 34756 23112
rect 36728 23103 36780 23112
rect 30380 22992 30432 23044
rect 32956 22992 33008 23044
rect 36728 23069 36737 23103
rect 36737 23069 36771 23103
rect 36771 23069 36780 23103
rect 36728 23060 36780 23069
rect 39856 23128 39908 23180
rect 40408 23128 40460 23180
rect 43168 23128 43220 23180
rect 37740 23103 37792 23112
rect 37740 23069 37749 23103
rect 37749 23069 37783 23103
rect 37783 23069 37792 23103
rect 37740 23060 37792 23069
rect 38660 22992 38712 23044
rect 43444 23060 43496 23112
rect 43076 22992 43128 23044
rect 30564 22924 30616 22976
rect 31300 22924 31352 22976
rect 36360 22967 36412 22976
rect 36360 22933 36369 22967
rect 36369 22933 36403 22967
rect 36403 22933 36412 22967
rect 36360 22924 36412 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 11704 22763 11756 22772
rect 11704 22729 11713 22763
rect 11713 22729 11747 22763
rect 11747 22729 11756 22763
rect 11704 22720 11756 22729
rect 23204 22720 23256 22772
rect 27528 22720 27580 22772
rect 27712 22720 27764 22772
rect 42800 22720 42852 22772
rect 42892 22720 42944 22772
rect 24584 22652 24636 22704
rect 26792 22652 26844 22704
rect 27344 22652 27396 22704
rect 28540 22652 28592 22704
rect 2596 22627 2648 22636
rect 2596 22593 2605 22627
rect 2605 22593 2639 22627
rect 2639 22593 2648 22627
rect 2596 22584 2648 22593
rect 7564 22584 7616 22636
rect 11428 22584 11480 22636
rect 16304 22627 16356 22636
rect 16304 22593 16313 22627
rect 16313 22593 16347 22627
rect 16347 22593 16356 22627
rect 16304 22584 16356 22593
rect 16396 22584 16448 22636
rect 17040 22627 17092 22636
rect 17040 22593 17049 22627
rect 17049 22593 17083 22627
rect 17083 22593 17092 22627
rect 17040 22584 17092 22593
rect 20996 22627 21048 22636
rect 20996 22593 21005 22627
rect 21005 22593 21039 22627
rect 21039 22593 21048 22627
rect 20996 22584 21048 22593
rect 21272 22627 21324 22636
rect 21272 22593 21281 22627
rect 21281 22593 21315 22627
rect 21315 22593 21324 22627
rect 21272 22584 21324 22593
rect 22560 22584 22612 22636
rect 24124 22627 24176 22636
rect 24124 22593 24133 22627
rect 24133 22593 24167 22627
rect 24167 22593 24176 22627
rect 24124 22584 24176 22593
rect 26608 22584 26660 22636
rect 27436 22627 27488 22636
rect 27436 22593 27445 22627
rect 27445 22593 27479 22627
rect 27479 22593 27488 22627
rect 27436 22584 27488 22593
rect 27712 22584 27764 22636
rect 28448 22627 28500 22636
rect 28448 22593 28457 22627
rect 28457 22593 28491 22627
rect 28491 22593 28500 22627
rect 28448 22584 28500 22593
rect 13084 22559 13136 22568
rect 13084 22525 13093 22559
rect 13093 22525 13127 22559
rect 13127 22525 13136 22559
rect 13084 22516 13136 22525
rect 15568 22559 15620 22568
rect 15568 22525 15577 22559
rect 15577 22525 15611 22559
rect 15611 22525 15620 22559
rect 15568 22516 15620 22525
rect 20352 22559 20404 22568
rect 20352 22525 20361 22559
rect 20361 22525 20395 22559
rect 20395 22525 20404 22559
rect 22008 22559 22060 22568
rect 20352 22516 20404 22525
rect 22008 22525 22017 22559
rect 22017 22525 22051 22559
rect 22051 22525 22060 22559
rect 22008 22516 22060 22525
rect 27344 22516 27396 22568
rect 30012 22652 30064 22704
rect 30840 22584 30892 22636
rect 31300 22627 31352 22636
rect 31300 22593 31309 22627
rect 31309 22593 31343 22627
rect 31343 22593 31352 22627
rect 31300 22584 31352 22593
rect 32956 22652 33008 22704
rect 34152 22652 34204 22704
rect 36360 22652 36412 22704
rect 33784 22627 33836 22636
rect 33784 22593 33793 22627
rect 33793 22593 33827 22627
rect 33827 22593 33836 22627
rect 33784 22584 33836 22593
rect 35624 22584 35676 22636
rect 36728 22584 36780 22636
rect 38936 22627 38988 22636
rect 36820 22516 36872 22568
rect 38936 22593 38945 22627
rect 38945 22593 38979 22627
rect 38979 22593 38988 22627
rect 38936 22584 38988 22593
rect 39028 22584 39080 22636
rect 41788 22584 41840 22636
rect 42800 22627 42852 22636
rect 41696 22559 41748 22568
rect 41696 22525 41705 22559
rect 41705 22525 41739 22559
rect 41739 22525 41748 22559
rect 41696 22516 41748 22525
rect 42800 22593 42809 22627
rect 42809 22593 42843 22627
rect 42843 22593 42852 22627
rect 42800 22584 42852 22593
rect 44180 22652 44232 22704
rect 43904 22627 43956 22636
rect 43904 22593 43913 22627
rect 43913 22593 43947 22627
rect 43947 22593 43956 22627
rect 43904 22584 43956 22593
rect 20720 22448 20772 22500
rect 33416 22448 33468 22500
rect 34060 22448 34112 22500
rect 42892 22448 42944 22500
rect 43444 22448 43496 22500
rect 3240 22380 3292 22432
rect 16764 22380 16816 22432
rect 18972 22423 19024 22432
rect 18972 22389 18981 22423
rect 18981 22389 19015 22423
rect 19015 22389 19024 22423
rect 18972 22380 19024 22389
rect 20444 22380 20496 22432
rect 25044 22380 25096 22432
rect 25504 22423 25556 22432
rect 25504 22389 25513 22423
rect 25513 22389 25547 22423
rect 25547 22389 25556 22423
rect 25504 22380 25556 22389
rect 28632 22423 28684 22432
rect 28632 22389 28641 22423
rect 28641 22389 28675 22423
rect 28675 22389 28684 22423
rect 28632 22380 28684 22389
rect 29092 22423 29144 22432
rect 29092 22389 29101 22423
rect 29101 22389 29135 22423
rect 29135 22389 29144 22423
rect 29092 22380 29144 22389
rect 29276 22423 29328 22432
rect 29276 22389 29285 22423
rect 29285 22389 29319 22423
rect 29319 22389 29328 22423
rect 29276 22380 29328 22389
rect 31208 22380 31260 22432
rect 34796 22380 34848 22432
rect 35440 22380 35492 22432
rect 37372 22380 37424 22432
rect 40316 22423 40368 22432
rect 40316 22389 40325 22423
rect 40325 22389 40359 22423
rect 40359 22389 40368 22423
rect 40316 22380 40368 22389
rect 42432 22380 42484 22432
rect 43260 22380 43312 22432
rect 44272 22380 44324 22432
rect 48320 22380 48372 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 14648 22219 14700 22228
rect 14648 22185 14657 22219
rect 14657 22185 14691 22219
rect 14691 22185 14700 22219
rect 14648 22176 14700 22185
rect 16488 22176 16540 22228
rect 18236 22176 18288 22228
rect 22560 22219 22612 22228
rect 22560 22185 22569 22219
rect 22569 22185 22603 22219
rect 22603 22185 22612 22219
rect 22560 22176 22612 22185
rect 22652 22176 22704 22228
rect 24768 22176 24820 22228
rect 24860 22176 24912 22228
rect 11612 22151 11664 22160
rect 11612 22117 11621 22151
rect 11621 22117 11655 22151
rect 11655 22117 11664 22151
rect 11612 22108 11664 22117
rect 3240 22083 3292 22092
rect 3240 22049 3249 22083
rect 3249 22049 3283 22083
rect 3283 22049 3292 22083
rect 3240 22040 3292 22049
rect 11428 22083 11480 22092
rect 11428 22049 11437 22083
rect 11437 22049 11471 22083
rect 11471 22049 11480 22083
rect 11428 22040 11480 22049
rect 11888 22083 11940 22092
rect 11888 22049 11897 22083
rect 11897 22049 11931 22083
rect 11931 22049 11940 22083
rect 11888 22040 11940 22049
rect 13084 22040 13136 22092
rect 15568 22040 15620 22092
rect 3424 22015 3476 22024
rect 3424 21981 3433 22015
rect 3433 21981 3467 22015
rect 3467 21981 3476 22015
rect 14464 22015 14516 22024
rect 3424 21972 3476 21981
rect 14464 21981 14473 22015
rect 14473 21981 14507 22015
rect 14507 21981 14516 22015
rect 14464 21972 14516 21981
rect 14740 22015 14792 22024
rect 14740 21981 14749 22015
rect 14749 21981 14783 22015
rect 14783 21981 14792 22015
rect 14740 21972 14792 21981
rect 17868 21972 17920 22024
rect 18328 22108 18380 22160
rect 18972 22040 19024 22092
rect 18328 22015 18380 22024
rect 18328 21981 18337 22015
rect 18337 21981 18371 22015
rect 18371 21981 18380 22015
rect 20996 22040 21048 22092
rect 22008 22083 22060 22092
rect 22008 22049 22017 22083
rect 22017 22049 22051 22083
rect 22051 22049 22060 22083
rect 22008 22040 22060 22049
rect 23572 22040 23624 22092
rect 23848 22108 23900 22160
rect 27252 22176 27304 22228
rect 27436 22176 27488 22228
rect 32220 22176 32272 22228
rect 33784 22176 33836 22228
rect 37740 22176 37792 22228
rect 39028 22219 39080 22228
rect 39028 22185 39037 22219
rect 39037 22185 39071 22219
rect 39071 22185 39080 22219
rect 39028 22176 39080 22185
rect 41788 22176 41840 22228
rect 42892 22176 42944 22228
rect 43168 22176 43220 22228
rect 43352 22176 43404 22228
rect 43904 22176 43956 22228
rect 44180 22219 44232 22228
rect 44180 22185 44189 22219
rect 44189 22185 44223 22219
rect 44223 22185 44232 22219
rect 44180 22176 44232 22185
rect 44272 22219 44324 22228
rect 44272 22185 44281 22219
rect 44281 22185 44315 22219
rect 44315 22185 44324 22219
rect 44272 22176 44324 22185
rect 27712 22108 27764 22160
rect 43444 22151 43496 22160
rect 43444 22117 43453 22151
rect 43453 22117 43487 22151
rect 43487 22117 43496 22151
rect 43444 22108 43496 22117
rect 26516 22040 26568 22092
rect 18328 21972 18380 21981
rect 22744 22015 22796 22024
rect 1584 21947 1636 21956
rect 1584 21913 1593 21947
rect 1593 21913 1627 21947
rect 1627 21913 1636 21947
rect 1584 21904 1636 21913
rect 16856 21904 16908 21956
rect 17040 21904 17092 21956
rect 22744 21981 22753 22015
rect 22753 21981 22787 22015
rect 22787 21981 22796 22015
rect 22744 21972 22796 21981
rect 33876 22040 33928 22092
rect 36084 22040 36136 22092
rect 36360 22083 36412 22092
rect 36360 22049 36369 22083
rect 36369 22049 36403 22083
rect 36403 22049 36412 22083
rect 36360 22040 36412 22049
rect 36820 22083 36872 22092
rect 36820 22049 36829 22083
rect 36829 22049 36863 22083
rect 36863 22049 36872 22083
rect 36820 22040 36872 22049
rect 37372 22083 37424 22092
rect 37372 22049 37381 22083
rect 37381 22049 37415 22083
rect 37415 22049 37424 22083
rect 37372 22040 37424 22049
rect 37924 22040 37976 22092
rect 43168 22083 43220 22092
rect 24124 21972 24176 22024
rect 24676 21972 24728 22024
rect 24952 21972 25004 22024
rect 25504 21972 25556 22024
rect 26240 21972 26292 22024
rect 26792 21972 26844 22024
rect 27528 22015 27580 22024
rect 27528 21981 27537 22015
rect 27537 21981 27571 22015
rect 27571 21981 27580 22015
rect 27528 21972 27580 21981
rect 27804 22015 27856 22024
rect 27804 21981 27813 22015
rect 27813 21981 27847 22015
rect 27847 21981 27856 22015
rect 27804 21972 27856 21981
rect 29092 21972 29144 22024
rect 29920 22015 29972 22024
rect 29920 21981 29929 22015
rect 29929 21981 29963 22015
rect 29963 21981 29972 22015
rect 29920 21972 29972 21981
rect 30104 22015 30156 22024
rect 30104 21981 30113 22015
rect 30113 21981 30147 22015
rect 30147 21981 30156 22015
rect 30104 21972 30156 21981
rect 30288 21972 30340 22024
rect 14280 21879 14332 21888
rect 14280 21845 14289 21879
rect 14289 21845 14323 21879
rect 14323 21845 14332 21879
rect 14280 21836 14332 21845
rect 16580 21836 16632 21888
rect 19984 21904 20036 21956
rect 20076 21904 20128 21956
rect 21180 21947 21232 21956
rect 21180 21913 21189 21947
rect 21189 21913 21223 21947
rect 21223 21913 21232 21947
rect 21180 21904 21232 21913
rect 28908 21904 28960 21956
rect 30840 21904 30892 21956
rect 31024 21972 31076 22024
rect 31208 22015 31260 22024
rect 31208 21981 31242 22015
rect 31242 21981 31260 22015
rect 31208 21972 31260 21981
rect 35256 22015 35308 22024
rect 17776 21836 17828 21888
rect 18236 21836 18288 21888
rect 22284 21836 22336 21888
rect 22376 21836 22428 21888
rect 23664 21879 23716 21888
rect 23664 21845 23673 21879
rect 23673 21845 23707 21879
rect 23707 21845 23716 21879
rect 26424 21879 26476 21888
rect 23664 21836 23716 21845
rect 26424 21845 26433 21879
rect 26433 21845 26467 21879
rect 26467 21845 26476 21879
rect 26424 21836 26476 21845
rect 26608 21879 26660 21888
rect 26608 21845 26617 21879
rect 26617 21845 26651 21879
rect 26651 21845 26660 21879
rect 26608 21836 26660 21845
rect 28080 21879 28132 21888
rect 28080 21845 28089 21879
rect 28089 21845 28123 21879
rect 28123 21845 28132 21879
rect 28080 21836 28132 21845
rect 29828 21836 29880 21888
rect 30932 21836 30984 21888
rect 31668 21836 31720 21888
rect 35256 21981 35265 22015
rect 35265 21981 35299 22015
rect 35299 21981 35308 22015
rect 35256 21972 35308 21981
rect 35440 22015 35492 22024
rect 35440 21981 35449 22015
rect 35449 21981 35483 22015
rect 35483 21981 35492 22015
rect 35440 21972 35492 21981
rect 38292 22015 38344 22024
rect 33324 21904 33376 21956
rect 35624 21904 35676 21956
rect 38292 21981 38301 22015
rect 38301 21981 38335 22015
rect 38335 21981 38344 22015
rect 38292 21972 38344 21981
rect 43168 22049 43177 22083
rect 43177 22049 43211 22083
rect 43211 22049 43220 22083
rect 43168 22040 43220 22049
rect 39212 22015 39264 22024
rect 39212 21981 39221 22015
rect 39221 21981 39255 22015
rect 39255 21981 39264 22015
rect 39212 21972 39264 21981
rect 39488 22015 39540 22024
rect 39488 21981 39497 22015
rect 39497 21981 39531 22015
rect 39531 21981 39540 22015
rect 39488 21972 39540 21981
rect 40316 21972 40368 22024
rect 41880 21972 41932 22024
rect 42432 22015 42484 22024
rect 42432 21981 42450 22015
rect 42450 21981 42484 22015
rect 42432 21972 42484 21981
rect 42708 22015 42760 22024
rect 42708 21981 42717 22015
rect 42717 21981 42751 22015
rect 42751 21981 42760 22015
rect 42708 21972 42760 21981
rect 43076 21972 43128 22024
rect 41696 21904 41748 21956
rect 43352 21904 43404 21956
rect 34152 21879 34204 21888
rect 34152 21845 34161 21879
rect 34161 21845 34195 21879
rect 34195 21845 34204 21879
rect 34152 21836 34204 21845
rect 35532 21836 35584 21888
rect 40960 21836 41012 21888
rect 46848 22083 46900 22092
rect 46848 22049 46857 22083
rect 46857 22049 46891 22083
rect 46891 22049 46900 22083
rect 46848 22040 46900 22049
rect 48320 22083 48372 22092
rect 48320 22049 48329 22083
rect 48329 22049 48363 22083
rect 48363 22049 48372 22083
rect 48320 22040 48372 22049
rect 47860 21904 47912 21956
rect 43628 21879 43680 21888
rect 43628 21845 43637 21879
rect 43637 21845 43671 21879
rect 43671 21845 43680 21879
rect 43628 21836 43680 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 11888 21632 11940 21684
rect 14280 21564 14332 21616
rect 16948 21564 17000 21616
rect 3424 21496 3476 21548
rect 13084 21496 13136 21548
rect 16580 21496 16632 21548
rect 17224 21539 17276 21548
rect 17224 21505 17233 21539
rect 17233 21505 17267 21539
rect 17267 21505 17276 21539
rect 17224 21496 17276 21505
rect 17776 21496 17828 21548
rect 17960 21564 18012 21616
rect 21272 21564 21324 21616
rect 16396 21428 16448 21480
rect 16856 21471 16908 21480
rect 16856 21437 16865 21471
rect 16865 21437 16899 21471
rect 16899 21437 16908 21471
rect 16856 21428 16908 21437
rect 17040 21471 17092 21480
rect 17040 21437 17049 21471
rect 17049 21437 17083 21471
rect 17083 21437 17092 21471
rect 17040 21428 17092 21437
rect 17500 21428 17552 21480
rect 17592 21428 17644 21480
rect 22376 21632 22428 21684
rect 23112 21632 23164 21684
rect 24952 21632 25004 21684
rect 26240 21632 26292 21684
rect 29736 21632 29788 21684
rect 30288 21632 30340 21684
rect 18144 21471 18196 21480
rect 18144 21437 18153 21471
rect 18153 21437 18187 21471
rect 18187 21437 18196 21471
rect 18144 21428 18196 21437
rect 23664 21539 23716 21548
rect 23664 21505 23673 21539
rect 23673 21505 23707 21539
rect 23707 21505 23716 21539
rect 24308 21539 24360 21548
rect 23664 21496 23716 21505
rect 24308 21505 24317 21539
rect 24317 21505 24351 21539
rect 24351 21505 24360 21539
rect 24308 21496 24360 21505
rect 25044 21496 25096 21548
rect 26424 21496 26476 21548
rect 26516 21428 26568 21480
rect 26700 21564 26752 21616
rect 27068 21564 27120 21616
rect 27252 21564 27304 21616
rect 27344 21496 27396 21548
rect 28632 21564 28684 21616
rect 30932 21564 30984 21616
rect 32496 21564 32548 21616
rect 29828 21539 29880 21548
rect 29828 21505 29862 21539
rect 29862 21505 29880 21539
rect 29828 21496 29880 21505
rect 33140 21632 33192 21684
rect 33324 21675 33376 21684
rect 33324 21641 33333 21675
rect 33333 21641 33367 21675
rect 33367 21641 33376 21675
rect 33324 21632 33376 21641
rect 35256 21632 35308 21684
rect 38292 21632 38344 21684
rect 42800 21632 42852 21684
rect 43352 21632 43404 21684
rect 47860 21675 47912 21684
rect 47860 21641 47869 21675
rect 47869 21641 47903 21675
rect 47903 21641 47912 21675
rect 47860 21632 47912 21641
rect 33784 21539 33836 21548
rect 27712 21428 27764 21480
rect 17868 21292 17920 21344
rect 20444 21292 20496 21344
rect 26332 21360 26384 21412
rect 28908 21403 28960 21412
rect 24676 21292 24728 21344
rect 27528 21292 27580 21344
rect 28908 21369 28917 21403
rect 28917 21369 28951 21403
rect 28951 21369 28960 21403
rect 28908 21360 28960 21369
rect 30656 21360 30708 21412
rect 33784 21505 33793 21539
rect 33793 21505 33827 21539
rect 33827 21505 33836 21539
rect 33784 21496 33836 21505
rect 34152 21564 34204 21616
rect 35532 21539 35584 21548
rect 35532 21505 35541 21539
rect 35541 21505 35575 21539
rect 35575 21505 35584 21539
rect 35532 21496 35584 21505
rect 36820 21496 36872 21548
rect 36912 21496 36964 21548
rect 37924 21539 37976 21548
rect 37924 21505 37933 21539
rect 37933 21505 37967 21539
rect 37967 21505 37976 21539
rect 37924 21496 37976 21505
rect 43628 21496 43680 21548
rect 44640 21496 44692 21548
rect 46388 21539 46440 21548
rect 46388 21505 46397 21539
rect 46397 21505 46431 21539
rect 46431 21505 46440 21539
rect 46388 21496 46440 21505
rect 47584 21496 47636 21548
rect 47768 21539 47820 21548
rect 47768 21505 47777 21539
rect 47777 21505 47811 21539
rect 47811 21505 47820 21539
rect 47768 21496 47820 21505
rect 33876 21428 33928 21480
rect 35624 21471 35676 21480
rect 35624 21437 35633 21471
rect 35633 21437 35667 21471
rect 35667 21437 35676 21471
rect 35624 21428 35676 21437
rect 42892 21471 42944 21480
rect 42892 21437 42901 21471
rect 42901 21437 42935 21471
rect 42935 21437 42944 21471
rect 42892 21428 42944 21437
rect 43076 21428 43128 21480
rect 30748 21292 30800 21344
rect 31024 21292 31076 21344
rect 39212 21360 39264 21412
rect 43996 21360 44048 21412
rect 44456 21360 44508 21412
rect 35992 21292 36044 21344
rect 37556 21292 37608 21344
rect 42800 21335 42852 21344
rect 42800 21301 42809 21335
rect 42809 21301 42843 21335
rect 42843 21301 42852 21335
rect 42800 21292 42852 21301
rect 43260 21292 43312 21344
rect 46664 21292 46716 21344
rect 47032 21335 47084 21344
rect 47032 21301 47041 21335
rect 47041 21301 47075 21335
rect 47075 21301 47084 21335
rect 47032 21292 47084 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 14464 21088 14516 21140
rect 13820 20952 13872 21004
rect 14924 21088 14976 21140
rect 17040 21020 17092 21072
rect 2044 20884 2096 20936
rect 14556 20884 14608 20936
rect 17868 20952 17920 21004
rect 20076 21088 20128 21140
rect 20444 21088 20496 21140
rect 23112 21020 23164 21072
rect 24308 21088 24360 21140
rect 23480 21020 23532 21072
rect 26148 21088 26200 21140
rect 26240 21088 26292 21140
rect 27528 21088 27580 21140
rect 29920 21088 29972 21140
rect 35532 21088 35584 21140
rect 35624 21088 35676 21140
rect 36912 21131 36964 21140
rect 36912 21097 36921 21131
rect 36921 21097 36955 21131
rect 36955 21097 36964 21131
rect 36912 21088 36964 21097
rect 30472 21020 30524 21072
rect 16396 20884 16448 20936
rect 16764 20927 16816 20936
rect 16764 20893 16773 20927
rect 16773 20893 16807 20927
rect 16807 20893 16816 20927
rect 16764 20884 16816 20893
rect 16948 20884 17000 20936
rect 16580 20816 16632 20868
rect 17592 20884 17644 20936
rect 19432 20884 19484 20936
rect 20444 20884 20496 20936
rect 32680 20952 32732 21004
rect 42708 20952 42760 21004
rect 47032 21020 47084 21072
rect 46664 20995 46716 21004
rect 46664 20961 46673 20995
rect 46673 20961 46707 20995
rect 46707 20961 46716 20995
rect 46664 20952 46716 20961
rect 48228 20995 48280 21004
rect 48228 20961 48237 20995
rect 48237 20961 48271 20995
rect 48271 20961 48280 20995
rect 48228 20952 48280 20961
rect 22376 20884 22428 20936
rect 17776 20816 17828 20868
rect 18144 20816 18196 20868
rect 22008 20816 22060 20868
rect 23296 20884 23348 20936
rect 17408 20748 17460 20800
rect 17500 20748 17552 20800
rect 18052 20748 18104 20800
rect 19340 20748 19392 20800
rect 19984 20748 20036 20800
rect 22928 20748 22980 20800
rect 25228 20884 25280 20936
rect 26332 20884 26384 20936
rect 27068 20927 27120 20936
rect 27068 20893 27077 20927
rect 27077 20893 27111 20927
rect 27111 20893 27120 20927
rect 27068 20884 27120 20893
rect 27344 20884 27396 20936
rect 26700 20748 26752 20800
rect 27252 20748 27304 20800
rect 28080 20884 28132 20936
rect 29920 20884 29972 20936
rect 30196 20927 30248 20936
rect 30196 20893 30205 20927
rect 30205 20893 30239 20927
rect 30239 20893 30248 20927
rect 30196 20884 30248 20893
rect 30380 20884 30432 20936
rect 30656 20927 30708 20936
rect 30656 20893 30665 20927
rect 30665 20893 30699 20927
rect 30699 20893 30708 20927
rect 30656 20884 30708 20893
rect 35348 20927 35400 20936
rect 35348 20893 35357 20927
rect 35357 20893 35391 20927
rect 35391 20893 35400 20927
rect 35348 20884 35400 20893
rect 36544 20927 36596 20936
rect 36544 20893 36553 20927
rect 36553 20893 36587 20927
rect 36587 20893 36596 20927
rect 36544 20884 36596 20893
rect 37372 20884 37424 20936
rect 43720 20816 43772 20868
rect 27620 20748 27672 20800
rect 28632 20748 28684 20800
rect 34888 20791 34940 20800
rect 34888 20757 34897 20791
rect 34897 20757 34931 20791
rect 34931 20757 34940 20791
rect 34888 20748 34940 20757
rect 44456 20748 44508 20800
rect 47308 20748 47360 20800
rect 47768 20748 47820 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 14648 20544 14700 20596
rect 16304 20544 16356 20596
rect 21180 20544 21232 20596
rect 30104 20544 30156 20596
rect 40592 20544 40644 20596
rect 43720 20587 43772 20596
rect 16948 20476 17000 20528
rect 2044 20451 2096 20460
rect 2044 20417 2053 20451
rect 2053 20417 2087 20451
rect 2087 20417 2096 20451
rect 2044 20408 2096 20417
rect 12532 20451 12584 20460
rect 12532 20417 12541 20451
rect 12541 20417 12575 20451
rect 12575 20417 12584 20451
rect 12532 20408 12584 20417
rect 12716 20451 12768 20460
rect 12716 20417 12725 20451
rect 12725 20417 12759 20451
rect 12759 20417 12768 20451
rect 12716 20408 12768 20417
rect 14648 20408 14700 20460
rect 15108 20451 15160 20460
rect 15108 20417 15117 20451
rect 15117 20417 15151 20451
rect 15151 20417 15160 20451
rect 15108 20408 15160 20417
rect 15292 20451 15344 20460
rect 15292 20417 15301 20451
rect 15301 20417 15335 20451
rect 15335 20417 15344 20451
rect 15292 20408 15344 20417
rect 2412 20340 2464 20392
rect 2780 20383 2832 20392
rect 2780 20349 2789 20383
rect 2789 20349 2823 20383
rect 2823 20349 2832 20383
rect 12808 20383 12860 20392
rect 2780 20340 2832 20349
rect 12808 20349 12817 20383
rect 12817 20349 12851 20383
rect 12851 20349 12860 20383
rect 12808 20340 12860 20349
rect 16672 20408 16724 20460
rect 17040 20451 17092 20460
rect 17040 20417 17049 20451
rect 17049 20417 17083 20451
rect 17083 20417 17092 20451
rect 17040 20408 17092 20417
rect 17500 20476 17552 20528
rect 17684 20476 17736 20528
rect 17132 20383 17184 20392
rect 17132 20349 17142 20383
rect 17142 20349 17176 20383
rect 17176 20349 17184 20383
rect 17132 20340 17184 20349
rect 17408 20408 17460 20460
rect 18144 20451 18196 20460
rect 18144 20417 18153 20451
rect 18153 20417 18187 20451
rect 18187 20417 18196 20451
rect 20720 20476 20772 20528
rect 34796 20519 34848 20528
rect 34796 20485 34805 20519
rect 34805 20485 34839 20519
rect 34839 20485 34848 20519
rect 34796 20476 34848 20485
rect 35348 20476 35400 20528
rect 41512 20476 41564 20528
rect 41696 20476 41748 20528
rect 43720 20553 43729 20587
rect 43729 20553 43763 20587
rect 43763 20553 43772 20587
rect 43720 20544 43772 20553
rect 18144 20408 18196 20417
rect 19340 20408 19392 20460
rect 27620 20408 27672 20460
rect 27712 20408 27764 20460
rect 28908 20408 28960 20460
rect 33692 20451 33744 20460
rect 33692 20417 33701 20451
rect 33701 20417 33735 20451
rect 33735 20417 33744 20451
rect 33692 20408 33744 20417
rect 17500 20340 17552 20392
rect 18420 20340 18472 20392
rect 12164 20204 12216 20256
rect 14556 20204 14608 20256
rect 15752 20247 15804 20256
rect 15752 20213 15761 20247
rect 15761 20213 15795 20247
rect 15795 20213 15804 20247
rect 15752 20204 15804 20213
rect 16212 20247 16264 20256
rect 16212 20213 16221 20247
rect 16221 20213 16255 20247
rect 16255 20213 16264 20247
rect 16212 20204 16264 20213
rect 17224 20272 17276 20324
rect 20260 20272 20312 20324
rect 17960 20204 18012 20256
rect 20352 20204 20404 20256
rect 29920 20272 29972 20324
rect 22376 20204 22428 20256
rect 33784 20204 33836 20256
rect 33876 20204 33928 20256
rect 35900 20408 35952 20460
rect 36544 20408 36596 20460
rect 39948 20408 40000 20460
rect 41880 20408 41932 20460
rect 44088 20408 44140 20460
rect 44180 20408 44232 20460
rect 45652 20408 45704 20460
rect 46204 20451 46256 20460
rect 46204 20417 46213 20451
rect 46213 20417 46247 20451
rect 46247 20417 46256 20451
rect 46204 20408 46256 20417
rect 37740 20340 37792 20392
rect 40132 20340 40184 20392
rect 41328 20340 41380 20392
rect 43904 20383 43956 20392
rect 40776 20272 40828 20324
rect 43904 20349 43913 20383
rect 43913 20349 43947 20383
rect 43947 20349 43956 20383
rect 43904 20340 43956 20349
rect 44456 20340 44508 20392
rect 34888 20204 34940 20256
rect 35992 20247 36044 20256
rect 35992 20213 36001 20247
rect 36001 20213 36035 20247
rect 36035 20213 36044 20247
rect 35992 20204 36044 20213
rect 36176 20247 36228 20256
rect 36176 20213 36185 20247
rect 36185 20213 36219 20247
rect 36219 20213 36228 20247
rect 36176 20204 36228 20213
rect 46296 20247 46348 20256
rect 46296 20213 46305 20247
rect 46305 20213 46339 20247
rect 46339 20213 46348 20247
rect 46296 20204 46348 20213
rect 46480 20204 46532 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 2412 20043 2464 20052
rect 2412 20009 2421 20043
rect 2421 20009 2455 20043
rect 2455 20009 2464 20043
rect 2412 20000 2464 20009
rect 12808 20000 12860 20052
rect 15292 20000 15344 20052
rect 17132 20000 17184 20052
rect 17684 20000 17736 20052
rect 19432 20000 19484 20052
rect 28908 20000 28960 20052
rect 33140 20000 33192 20052
rect 20444 19932 20496 19984
rect 35348 20000 35400 20052
rect 35900 20000 35952 20052
rect 44088 20043 44140 20052
rect 33784 19975 33836 19984
rect 33784 19941 33793 19975
rect 33793 19941 33827 19975
rect 33827 19941 33836 19975
rect 33784 19932 33836 19941
rect 16948 19864 17000 19916
rect 2504 19839 2556 19848
rect 2504 19805 2513 19839
rect 2513 19805 2547 19839
rect 2547 19805 2556 19839
rect 2504 19796 2556 19805
rect 3148 19796 3200 19848
rect 16304 19839 16356 19848
rect 12164 19771 12216 19780
rect 12164 19737 12198 19771
rect 12198 19737 12216 19771
rect 12164 19728 12216 19737
rect 12256 19728 12308 19780
rect 14556 19771 14608 19780
rect 14556 19737 14590 19771
rect 14590 19737 14608 19771
rect 14556 19728 14608 19737
rect 16304 19805 16313 19839
rect 16313 19805 16347 19839
rect 16347 19805 16356 19839
rect 16304 19796 16356 19805
rect 17684 19839 17736 19848
rect 17684 19805 17693 19839
rect 17693 19805 17727 19839
rect 17727 19805 17736 19839
rect 17684 19796 17736 19805
rect 19984 19796 20036 19848
rect 20352 19839 20404 19848
rect 17500 19728 17552 19780
rect 20352 19805 20361 19839
rect 20361 19805 20395 19839
rect 20395 19805 20404 19839
rect 20352 19796 20404 19805
rect 21456 19796 21508 19848
rect 22008 19839 22060 19848
rect 22008 19805 22017 19839
rect 22017 19805 22051 19839
rect 22051 19805 22060 19839
rect 22008 19796 22060 19805
rect 22100 19796 22152 19848
rect 25228 19796 25280 19848
rect 26332 19864 26384 19916
rect 31668 19907 31720 19916
rect 31668 19873 31677 19907
rect 31677 19873 31711 19907
rect 31711 19873 31720 19907
rect 31668 19864 31720 19873
rect 33600 19907 33652 19916
rect 33600 19873 33609 19907
rect 33609 19873 33643 19907
rect 33643 19873 33652 19907
rect 33600 19864 33652 19873
rect 33692 19864 33744 19916
rect 26056 19728 26108 19780
rect 29184 19839 29236 19848
rect 29184 19805 29193 19839
rect 29193 19805 29227 19839
rect 29227 19805 29236 19839
rect 29920 19839 29972 19848
rect 29184 19796 29236 19805
rect 29920 19805 29929 19839
rect 29929 19805 29963 19839
rect 29963 19805 29972 19839
rect 29920 19796 29972 19805
rect 30196 19839 30248 19848
rect 30196 19805 30205 19839
rect 30205 19805 30239 19839
rect 30239 19805 30248 19839
rect 30196 19796 30248 19805
rect 30380 19839 30432 19848
rect 30380 19805 30389 19839
rect 30389 19805 30423 19839
rect 30423 19805 30432 19839
rect 30380 19796 30432 19805
rect 33876 19839 33928 19848
rect 33876 19805 33885 19839
rect 33885 19805 33919 19839
rect 33919 19805 33928 19839
rect 33876 19796 33928 19805
rect 35440 19796 35492 19848
rect 39212 19839 39264 19848
rect 39212 19805 39221 19839
rect 39221 19805 39255 19839
rect 39255 19805 39264 19839
rect 39212 19796 39264 19805
rect 40132 19796 40184 19848
rect 44088 20009 44097 20043
rect 44097 20009 44131 20043
rect 44131 20009 44140 20043
rect 44088 20000 44140 20009
rect 41788 19864 41840 19916
rect 40500 19796 40552 19848
rect 40776 19796 40828 19848
rect 41328 19839 41380 19848
rect 41328 19805 41337 19839
rect 41337 19805 41371 19839
rect 41371 19805 41380 19839
rect 41328 19796 41380 19805
rect 32312 19728 32364 19780
rect 13452 19660 13504 19712
rect 15108 19660 15160 19712
rect 22192 19660 22244 19712
rect 25688 19660 25740 19712
rect 27344 19660 27396 19712
rect 28724 19703 28776 19712
rect 28724 19669 28733 19703
rect 28733 19669 28767 19703
rect 28767 19669 28776 19703
rect 28724 19660 28776 19669
rect 32864 19660 32916 19712
rect 33784 19728 33836 19780
rect 39948 19728 40000 19780
rect 33140 19660 33192 19712
rect 40132 19660 40184 19712
rect 41696 19796 41748 19848
rect 43996 19864 44048 19916
rect 46296 19932 46348 19984
rect 46480 19907 46532 19916
rect 46480 19873 46489 19907
rect 46489 19873 46523 19907
rect 46523 19873 46532 19907
rect 46480 19864 46532 19873
rect 48228 19907 48280 19916
rect 48228 19873 48237 19907
rect 48237 19873 48271 19907
rect 48271 19873 48280 19907
rect 48228 19864 48280 19873
rect 44364 19839 44416 19848
rect 44364 19805 44373 19839
rect 44373 19805 44407 19839
rect 44407 19805 44416 19839
rect 44364 19796 44416 19805
rect 44272 19728 44324 19780
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 12532 19456 12584 19508
rect 14648 19499 14700 19508
rect 14648 19465 14657 19499
rect 14657 19465 14691 19499
rect 14691 19465 14700 19499
rect 14648 19456 14700 19465
rect 15752 19456 15804 19508
rect 17684 19456 17736 19508
rect 25228 19499 25280 19508
rect 25228 19465 25237 19499
rect 25237 19465 25271 19499
rect 25271 19465 25280 19499
rect 25228 19456 25280 19465
rect 13360 19388 13412 19440
rect 14464 19388 14516 19440
rect 15292 19388 15344 19440
rect 13452 19363 13504 19372
rect 13452 19329 13461 19363
rect 13461 19329 13495 19363
rect 13495 19329 13504 19363
rect 13452 19320 13504 19329
rect 16672 19388 16724 19440
rect 13544 19252 13596 19304
rect 13820 19252 13872 19304
rect 14924 19252 14976 19304
rect 16948 19320 17000 19372
rect 17224 19363 17276 19372
rect 17224 19329 17233 19363
rect 17233 19329 17267 19363
rect 17267 19329 17276 19363
rect 17224 19320 17276 19329
rect 17592 19388 17644 19440
rect 17408 19320 17460 19372
rect 20076 19388 20128 19440
rect 20628 19431 20680 19440
rect 20628 19397 20637 19431
rect 20637 19397 20671 19431
rect 20671 19397 20680 19431
rect 20628 19388 20680 19397
rect 21180 19388 21232 19440
rect 30380 19456 30432 19508
rect 32312 19499 32364 19508
rect 28724 19431 28776 19440
rect 19984 19320 20036 19372
rect 22192 19363 22244 19372
rect 15108 19184 15160 19236
rect 16488 19252 16540 19304
rect 19248 19295 19300 19304
rect 19248 19261 19257 19295
rect 19257 19261 19291 19295
rect 19291 19261 19300 19295
rect 19248 19252 19300 19261
rect 22192 19329 22201 19363
rect 22201 19329 22235 19363
rect 22235 19329 22244 19363
rect 22192 19320 22244 19329
rect 22376 19363 22428 19372
rect 22376 19329 22385 19363
rect 22385 19329 22419 19363
rect 22419 19329 22428 19363
rect 22376 19320 22428 19329
rect 25228 19320 25280 19372
rect 27344 19363 27396 19372
rect 27344 19329 27353 19363
rect 27353 19329 27387 19363
rect 27387 19329 27396 19363
rect 27344 19320 27396 19329
rect 27436 19320 27488 19372
rect 28724 19397 28758 19431
rect 28758 19397 28776 19431
rect 28724 19388 28776 19397
rect 32312 19465 32321 19499
rect 32321 19465 32355 19499
rect 32355 19465 32364 19499
rect 32312 19456 32364 19465
rect 32404 19456 32456 19508
rect 33324 19456 33376 19508
rect 33416 19388 33468 19440
rect 28540 19320 28592 19372
rect 30656 19363 30708 19372
rect 30656 19329 30665 19363
rect 30665 19329 30699 19363
rect 30699 19329 30708 19363
rect 30656 19320 30708 19329
rect 30840 19363 30892 19372
rect 30840 19329 30849 19363
rect 30849 19329 30883 19363
rect 30883 19329 30892 19363
rect 30840 19320 30892 19329
rect 31300 19320 31352 19372
rect 31852 19320 31904 19372
rect 32404 19320 32456 19372
rect 32864 19363 32916 19372
rect 32864 19329 32872 19363
rect 32872 19329 32906 19363
rect 32906 19329 32916 19363
rect 32864 19320 32916 19329
rect 33140 19320 33192 19372
rect 34704 19456 34756 19508
rect 40224 19456 40276 19508
rect 43904 19456 43956 19508
rect 33876 19388 33928 19440
rect 23020 19252 23072 19304
rect 12624 19116 12676 19168
rect 20628 19184 20680 19236
rect 22836 19184 22888 19236
rect 19708 19159 19760 19168
rect 19708 19125 19717 19159
rect 19717 19125 19751 19159
rect 19751 19125 19760 19159
rect 19708 19116 19760 19125
rect 22008 19159 22060 19168
rect 22008 19125 22017 19159
rect 22017 19125 22051 19159
rect 22051 19125 22060 19159
rect 22008 19116 22060 19125
rect 24768 19159 24820 19168
rect 24768 19125 24777 19159
rect 24777 19125 24811 19159
rect 24811 19125 24820 19159
rect 24768 19116 24820 19125
rect 31576 19252 31628 19304
rect 33784 19320 33836 19372
rect 34428 19363 34480 19372
rect 34428 19329 34437 19363
rect 34437 19329 34471 19363
rect 34471 19329 34480 19363
rect 34428 19320 34480 19329
rect 40408 19388 40460 19440
rect 43996 19388 44048 19440
rect 39948 19363 40000 19372
rect 37740 19295 37792 19304
rect 37740 19261 37749 19295
rect 37749 19261 37783 19295
rect 37783 19261 37792 19295
rect 37740 19252 37792 19261
rect 39948 19329 39957 19363
rect 39957 19329 39991 19363
rect 39991 19329 40000 19363
rect 39948 19320 40000 19329
rect 40592 19320 40644 19372
rect 40960 19363 41012 19372
rect 40960 19329 40969 19363
rect 40969 19329 41003 19363
rect 41003 19329 41012 19363
rect 40960 19320 41012 19329
rect 41788 19363 41840 19372
rect 41788 19329 41797 19363
rect 41797 19329 41831 19363
rect 41831 19329 41840 19363
rect 41788 19320 41840 19329
rect 43444 19363 43496 19372
rect 43444 19329 43453 19363
rect 43453 19329 43487 19363
rect 43487 19329 43496 19363
rect 43444 19320 43496 19329
rect 44272 19363 44324 19372
rect 44272 19329 44281 19363
rect 44281 19329 44315 19363
rect 44315 19329 44324 19363
rect 44272 19320 44324 19329
rect 44364 19363 44416 19372
rect 44364 19329 44373 19363
rect 44373 19329 44407 19363
rect 44407 19329 44416 19363
rect 44364 19320 44416 19329
rect 44640 19320 44692 19372
rect 47216 19363 47268 19372
rect 40224 19295 40276 19304
rect 40224 19261 40233 19295
rect 40233 19261 40267 19295
rect 40267 19261 40276 19295
rect 40224 19252 40276 19261
rect 40776 19252 40828 19304
rect 44548 19252 44600 19304
rect 47216 19329 47225 19363
rect 47225 19329 47259 19363
rect 47259 19329 47268 19363
rect 47216 19320 47268 19329
rect 47584 19320 47636 19372
rect 39948 19184 40000 19236
rect 29184 19116 29236 19168
rect 30472 19159 30524 19168
rect 30472 19125 30481 19159
rect 30481 19125 30515 19159
rect 30515 19125 30524 19159
rect 30472 19116 30524 19125
rect 33692 19116 33744 19168
rect 34796 19116 34848 19168
rect 40868 19116 40920 19168
rect 41236 19116 41288 19168
rect 41604 19159 41656 19168
rect 41604 19125 41613 19159
rect 41613 19125 41647 19159
rect 41647 19125 41656 19159
rect 41604 19116 41656 19125
rect 44180 19116 44232 19168
rect 47124 19159 47176 19168
rect 47124 19125 47133 19159
rect 47133 19125 47167 19159
rect 47167 19125 47176 19159
rect 47124 19116 47176 19125
rect 47768 19159 47820 19168
rect 47768 19125 47777 19159
rect 47777 19125 47811 19159
rect 47811 19125 47820 19159
rect 47768 19116 47820 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 19248 18912 19300 18964
rect 25044 18912 25096 18964
rect 25228 18955 25280 18964
rect 25228 18921 25237 18955
rect 25237 18921 25271 18955
rect 25271 18921 25280 18955
rect 25228 18912 25280 18921
rect 31576 18955 31628 18964
rect 23020 18844 23072 18896
rect 28632 18887 28684 18896
rect 28632 18853 28641 18887
rect 28641 18853 28675 18887
rect 28675 18853 28684 18887
rect 28632 18844 28684 18853
rect 31576 18921 31585 18955
rect 31585 18921 31619 18955
rect 31619 18921 31628 18955
rect 31576 18912 31628 18921
rect 39212 18912 39264 18964
rect 39948 18912 40000 18964
rect 40776 18955 40828 18964
rect 40776 18921 40785 18955
rect 40785 18921 40819 18955
rect 40819 18921 40828 18955
rect 40776 18912 40828 18921
rect 33508 18844 33560 18896
rect 15108 18776 15160 18828
rect 2044 18751 2096 18760
rect 2044 18717 2053 18751
rect 2053 18717 2087 18751
rect 2087 18717 2096 18751
rect 2044 18708 2096 18717
rect 15292 18708 15344 18760
rect 16764 18776 16816 18828
rect 22836 18819 22888 18828
rect 16948 18708 17000 18760
rect 22836 18785 22845 18819
rect 22845 18785 22879 18819
rect 22879 18785 22888 18819
rect 22836 18776 22888 18785
rect 28540 18776 28592 18828
rect 19340 18708 19392 18760
rect 19708 18751 19760 18760
rect 19708 18717 19742 18751
rect 19742 18717 19760 18751
rect 19708 18708 19760 18717
rect 22008 18708 22060 18760
rect 23940 18708 23992 18760
rect 17408 18640 17460 18692
rect 24768 18708 24820 18760
rect 25228 18708 25280 18760
rect 25596 18708 25648 18760
rect 28448 18751 28500 18760
rect 28448 18717 28457 18751
rect 28457 18717 28491 18751
rect 28491 18717 28500 18751
rect 28448 18708 28500 18717
rect 29184 18708 29236 18760
rect 29828 18708 29880 18760
rect 34796 18776 34848 18828
rect 31668 18708 31720 18760
rect 35440 18708 35492 18760
rect 40316 18844 40368 18896
rect 41788 18912 41840 18964
rect 42892 18844 42944 18896
rect 44548 18844 44600 18896
rect 45468 18844 45520 18896
rect 40224 18776 40276 18828
rect 36452 18708 36504 18760
rect 37740 18708 37792 18760
rect 24860 18683 24912 18692
rect 16856 18615 16908 18624
rect 16856 18581 16865 18615
rect 16865 18581 16899 18615
rect 16899 18581 16908 18615
rect 16856 18572 16908 18581
rect 20536 18572 20588 18624
rect 21456 18615 21508 18624
rect 21456 18581 21465 18615
rect 21465 18581 21499 18615
rect 21499 18581 21508 18615
rect 21456 18572 21508 18581
rect 23756 18572 23808 18624
rect 24860 18649 24869 18683
rect 24869 18649 24903 18683
rect 24903 18649 24912 18683
rect 24860 18640 24912 18649
rect 25136 18572 25188 18624
rect 30472 18683 30524 18692
rect 30472 18649 30506 18683
rect 30506 18649 30524 18683
rect 30472 18640 30524 18649
rect 31760 18640 31812 18692
rect 33048 18640 33100 18692
rect 40040 18708 40092 18760
rect 41236 18751 41288 18760
rect 41236 18717 41245 18751
rect 41245 18717 41279 18751
rect 41279 18717 41288 18751
rect 41236 18708 41288 18717
rect 41420 18751 41472 18760
rect 41420 18717 41429 18751
rect 41429 18717 41463 18751
rect 41463 18717 41472 18751
rect 41420 18708 41472 18717
rect 40224 18640 40276 18692
rect 40592 18683 40644 18692
rect 40592 18649 40601 18683
rect 40601 18649 40635 18683
rect 40635 18649 40644 18683
rect 40592 18640 40644 18649
rect 41880 18640 41932 18692
rect 42892 18708 42944 18760
rect 44272 18776 44324 18828
rect 44364 18776 44416 18828
rect 47768 18844 47820 18896
rect 44640 18708 44692 18760
rect 45376 18751 45428 18760
rect 45376 18717 45385 18751
rect 45385 18717 45419 18751
rect 45419 18717 45428 18751
rect 45376 18708 45428 18717
rect 47124 18776 47176 18828
rect 48228 18819 48280 18828
rect 48228 18785 48237 18819
rect 48237 18785 48271 18819
rect 48271 18785 48280 18819
rect 48228 18776 48280 18785
rect 44548 18683 44600 18692
rect 44548 18649 44557 18683
rect 44557 18649 44591 18683
rect 44591 18649 44600 18683
rect 44548 18640 44600 18649
rect 45560 18683 45612 18692
rect 45560 18649 45569 18683
rect 45569 18649 45603 18683
rect 45603 18649 45612 18683
rect 45560 18640 45612 18649
rect 45652 18640 45704 18692
rect 46480 18640 46532 18692
rect 27160 18572 27212 18624
rect 36544 18615 36596 18624
rect 36544 18581 36553 18615
rect 36553 18581 36587 18615
rect 36587 18581 36596 18615
rect 36544 18572 36596 18581
rect 43444 18572 43496 18624
rect 43904 18572 43956 18624
rect 45192 18615 45244 18624
rect 45192 18581 45201 18615
rect 45201 18581 45235 18615
rect 45235 18581 45244 18615
rect 45192 18572 45244 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 19984 18411 20036 18420
rect 19984 18377 19993 18411
rect 19993 18377 20027 18411
rect 20027 18377 20036 18411
rect 19984 18368 20036 18377
rect 23940 18411 23992 18420
rect 23940 18377 23949 18411
rect 23949 18377 23983 18411
rect 23983 18377 23992 18411
rect 23940 18368 23992 18377
rect 25044 18368 25096 18420
rect 21456 18300 21508 18352
rect 23572 18343 23624 18352
rect 23572 18309 23581 18343
rect 23581 18309 23615 18343
rect 23615 18309 23624 18343
rect 23572 18300 23624 18309
rect 23664 18300 23716 18352
rect 2044 18275 2096 18284
rect 2044 18241 2053 18275
rect 2053 18241 2087 18275
rect 2087 18241 2096 18275
rect 2044 18232 2096 18241
rect 13360 18232 13412 18284
rect 13544 18275 13596 18284
rect 13544 18241 13553 18275
rect 13553 18241 13587 18275
rect 13587 18241 13596 18275
rect 13544 18232 13596 18241
rect 13728 18275 13780 18284
rect 13728 18241 13737 18275
rect 13737 18241 13771 18275
rect 13771 18241 13780 18275
rect 13728 18232 13780 18241
rect 16120 18275 16172 18284
rect 16120 18241 16129 18275
rect 16129 18241 16163 18275
rect 16163 18241 16172 18275
rect 16120 18232 16172 18241
rect 16304 18275 16356 18284
rect 16304 18241 16313 18275
rect 16313 18241 16347 18275
rect 16347 18241 16356 18275
rect 16304 18232 16356 18241
rect 17132 18232 17184 18284
rect 18328 18275 18380 18284
rect 2228 18207 2280 18216
rect 2228 18173 2237 18207
rect 2237 18173 2271 18207
rect 2271 18173 2280 18207
rect 2228 18164 2280 18173
rect 2780 18207 2832 18216
rect 2780 18173 2789 18207
rect 2789 18173 2823 18207
rect 2823 18173 2832 18207
rect 2780 18164 2832 18173
rect 12532 18164 12584 18216
rect 12624 18207 12676 18216
rect 12624 18173 12633 18207
rect 12633 18173 12667 18207
rect 12667 18173 12676 18207
rect 12624 18164 12676 18173
rect 14740 18164 14792 18216
rect 18328 18241 18337 18275
rect 18337 18241 18371 18275
rect 18371 18241 18380 18275
rect 18328 18232 18380 18241
rect 20168 18275 20220 18284
rect 20168 18241 20177 18275
rect 20177 18241 20211 18275
rect 20211 18241 20220 18275
rect 20168 18232 20220 18241
rect 20536 18232 20588 18284
rect 24032 18232 24084 18284
rect 25136 18300 25188 18352
rect 28448 18368 28500 18420
rect 30656 18368 30708 18420
rect 29736 18300 29788 18352
rect 24768 18232 24820 18284
rect 27160 18275 27212 18284
rect 27160 18241 27169 18275
rect 27169 18241 27203 18275
rect 27203 18241 27212 18275
rect 27160 18232 27212 18241
rect 27252 18232 27304 18284
rect 27528 18232 27580 18284
rect 27712 18232 27764 18284
rect 29828 18232 29880 18284
rect 30564 18232 30616 18284
rect 30748 18275 30800 18284
rect 30748 18241 30757 18275
rect 30757 18241 30791 18275
rect 30791 18241 30800 18275
rect 30748 18232 30800 18241
rect 33784 18275 33836 18284
rect 33784 18241 33793 18275
rect 33793 18241 33827 18275
rect 33827 18241 33836 18275
rect 33784 18232 33836 18241
rect 34796 18368 34848 18420
rect 34428 18300 34480 18352
rect 36544 18343 36596 18352
rect 36544 18309 36553 18343
rect 36553 18309 36587 18343
rect 36587 18309 36596 18343
rect 36544 18300 36596 18309
rect 40408 18411 40460 18420
rect 36360 18275 36412 18284
rect 21272 18164 21324 18216
rect 21640 18096 21692 18148
rect 24860 18096 24912 18148
rect 12716 18028 12768 18080
rect 16580 18028 16632 18080
rect 18328 18028 18380 18080
rect 23848 18028 23900 18080
rect 23940 18028 23992 18080
rect 33968 18071 34020 18080
rect 33968 18037 33977 18071
rect 33977 18037 34011 18071
rect 34011 18037 34020 18071
rect 36360 18241 36369 18275
rect 36369 18241 36403 18275
rect 36403 18241 36412 18275
rect 36360 18232 36412 18241
rect 34704 18096 34756 18148
rect 35348 18139 35400 18148
rect 35348 18105 35357 18139
rect 35357 18105 35391 18139
rect 35391 18105 35400 18139
rect 35348 18096 35400 18105
rect 36176 18096 36228 18148
rect 40408 18377 40417 18411
rect 40417 18377 40451 18411
rect 40451 18377 40460 18411
rect 40408 18368 40460 18377
rect 44364 18368 44416 18420
rect 45468 18368 45520 18420
rect 37740 18300 37792 18352
rect 40040 18343 40092 18352
rect 40040 18309 40049 18343
rect 40049 18309 40083 18343
rect 40083 18309 40092 18343
rect 40040 18300 40092 18309
rect 40224 18343 40276 18352
rect 40224 18309 40233 18343
rect 40233 18309 40267 18343
rect 40267 18309 40276 18343
rect 40224 18300 40276 18309
rect 41604 18300 41656 18352
rect 44272 18300 44324 18352
rect 45192 18300 45244 18352
rect 41144 18275 41196 18284
rect 41144 18241 41153 18275
rect 41153 18241 41187 18275
rect 41187 18241 41196 18275
rect 41144 18232 41196 18241
rect 43904 18275 43956 18284
rect 43904 18241 43913 18275
rect 43913 18241 43947 18275
rect 43947 18241 43956 18275
rect 43904 18232 43956 18241
rect 45468 18232 45520 18284
rect 33968 18028 34020 18037
rect 36084 18028 36136 18080
rect 40684 18028 40736 18080
rect 41328 18071 41380 18080
rect 41328 18037 41337 18071
rect 41337 18037 41371 18071
rect 41371 18037 41380 18071
rect 41328 18028 41380 18037
rect 43904 18028 43956 18080
rect 44640 18028 44692 18080
rect 48320 18028 48372 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 2228 17824 2280 17876
rect 12624 17824 12676 17876
rect 13728 17824 13780 17876
rect 15936 17824 15988 17876
rect 16120 17824 16172 17876
rect 16304 17824 16356 17876
rect 17132 17867 17184 17876
rect 17132 17833 17141 17867
rect 17141 17833 17175 17867
rect 17175 17833 17184 17867
rect 17132 17824 17184 17833
rect 19248 17824 19300 17876
rect 21088 17824 21140 17876
rect 23664 17824 23716 17876
rect 28908 17824 28960 17876
rect 2596 17620 2648 17672
rect 6736 17620 6788 17672
rect 12072 17620 12124 17672
rect 12256 17663 12308 17672
rect 12256 17629 12265 17663
rect 12265 17629 12299 17663
rect 12299 17629 12308 17663
rect 12256 17620 12308 17629
rect 12900 17620 12952 17672
rect 14464 17663 14516 17672
rect 14464 17629 14473 17663
rect 14473 17629 14507 17663
rect 14507 17629 14516 17663
rect 14464 17620 14516 17629
rect 14740 17663 14792 17672
rect 14740 17629 14749 17663
rect 14749 17629 14783 17663
rect 14783 17629 14792 17663
rect 14740 17620 14792 17629
rect 12532 17595 12584 17604
rect 12532 17561 12566 17595
rect 12566 17561 12584 17595
rect 12532 17552 12584 17561
rect 11980 17484 12032 17536
rect 12072 17484 12124 17536
rect 13268 17484 13320 17536
rect 15108 17620 15160 17672
rect 16856 17688 16908 17740
rect 19340 17688 19392 17740
rect 16672 17663 16724 17672
rect 15200 17552 15252 17604
rect 16672 17629 16681 17663
rect 16681 17629 16715 17663
rect 16715 17629 16724 17663
rect 16672 17620 16724 17629
rect 19432 17663 19484 17672
rect 19432 17629 19441 17663
rect 19441 17629 19475 17663
rect 19475 17629 19484 17663
rect 19432 17620 19484 17629
rect 20260 17620 20312 17672
rect 23204 17688 23256 17740
rect 29460 17688 29512 17740
rect 33784 17824 33836 17876
rect 35348 17824 35400 17876
rect 36360 17824 36412 17876
rect 40040 17867 40092 17876
rect 40040 17833 40049 17867
rect 40049 17833 40083 17867
rect 40083 17833 40092 17867
rect 40040 17824 40092 17833
rect 44548 17824 44600 17876
rect 45376 17867 45428 17876
rect 45376 17833 45385 17867
rect 45385 17833 45419 17867
rect 45419 17833 45428 17867
rect 45376 17824 45428 17833
rect 36452 17756 36504 17808
rect 44364 17756 44416 17808
rect 37740 17688 37792 17740
rect 44456 17688 44508 17740
rect 46848 17731 46900 17740
rect 46848 17697 46857 17731
rect 46857 17697 46891 17731
rect 46891 17697 46900 17731
rect 46848 17688 46900 17697
rect 48320 17731 48372 17740
rect 48320 17697 48329 17731
rect 48329 17697 48363 17731
rect 48363 17697 48372 17731
rect 48320 17688 48372 17697
rect 20444 17620 20496 17672
rect 23756 17663 23808 17672
rect 18512 17552 18564 17604
rect 23756 17629 23765 17663
rect 23765 17629 23799 17663
rect 23799 17629 23808 17663
rect 23756 17620 23808 17629
rect 23940 17663 23992 17672
rect 23940 17629 23949 17663
rect 23949 17629 23983 17663
rect 23983 17629 23992 17663
rect 23940 17620 23992 17629
rect 29920 17663 29972 17672
rect 29920 17629 29929 17663
rect 29929 17629 29963 17663
rect 29963 17629 29972 17663
rect 30196 17663 30248 17672
rect 29920 17620 29972 17629
rect 30196 17629 30205 17663
rect 30205 17629 30239 17663
rect 30239 17629 30248 17663
rect 30196 17620 30248 17629
rect 31116 17663 31168 17672
rect 16948 17484 17000 17536
rect 19432 17484 19484 17536
rect 21732 17527 21784 17536
rect 21732 17493 21741 17527
rect 21741 17493 21775 17527
rect 21775 17493 21784 17527
rect 21732 17484 21784 17493
rect 23480 17552 23532 17604
rect 30288 17552 30340 17604
rect 29000 17484 29052 17536
rect 29184 17527 29236 17536
rect 29184 17493 29193 17527
rect 29193 17493 29227 17527
rect 29227 17493 29236 17527
rect 29184 17484 29236 17493
rect 30104 17484 30156 17536
rect 31116 17629 31125 17663
rect 31125 17629 31159 17663
rect 31159 17629 31168 17663
rect 31116 17620 31168 17629
rect 31300 17663 31352 17672
rect 31300 17629 31309 17663
rect 31309 17629 31343 17663
rect 31343 17629 31352 17663
rect 31300 17620 31352 17629
rect 31576 17620 31628 17672
rect 33784 17620 33836 17672
rect 34796 17552 34848 17604
rect 36360 17620 36412 17672
rect 40316 17620 40368 17672
rect 41328 17663 41380 17672
rect 40960 17595 41012 17604
rect 40960 17561 40969 17595
rect 40969 17561 41003 17595
rect 41003 17561 41012 17595
rect 40960 17552 41012 17561
rect 41328 17629 41337 17663
rect 41337 17629 41371 17663
rect 41371 17629 41380 17663
rect 41328 17620 41380 17629
rect 43720 17663 43772 17672
rect 43720 17629 43729 17663
rect 43729 17629 43763 17663
rect 43763 17629 43772 17663
rect 43720 17620 43772 17629
rect 41604 17552 41656 17604
rect 40132 17484 40184 17536
rect 41144 17527 41196 17536
rect 41144 17493 41153 17527
rect 41153 17493 41187 17527
rect 41187 17493 41196 17527
rect 41144 17484 41196 17493
rect 41512 17527 41564 17536
rect 41512 17493 41521 17527
rect 41521 17493 41555 17527
rect 41555 17493 41564 17527
rect 41512 17484 41564 17493
rect 43352 17484 43404 17536
rect 44640 17620 44692 17672
rect 45468 17663 45520 17672
rect 45468 17629 45477 17663
rect 45477 17629 45511 17663
rect 45511 17629 45520 17663
rect 45468 17620 45520 17629
rect 44272 17552 44324 17604
rect 47860 17552 47912 17604
rect 44548 17484 44600 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 1952 17280 2004 17332
rect 13268 17323 13320 17332
rect 12256 17212 12308 17264
rect 11980 17144 12032 17196
rect 13268 17289 13277 17323
rect 13277 17289 13311 17323
rect 13311 17289 13320 17323
rect 13268 17280 13320 17289
rect 15108 17323 15160 17332
rect 15108 17289 15117 17323
rect 15117 17289 15151 17323
rect 15151 17289 15160 17323
rect 15108 17280 15160 17289
rect 16948 17323 17000 17332
rect 16948 17289 16957 17323
rect 16957 17289 16991 17323
rect 16991 17289 17000 17323
rect 16948 17280 17000 17289
rect 17776 17280 17828 17332
rect 18052 17280 18104 17332
rect 18512 17323 18564 17332
rect 18512 17289 18521 17323
rect 18521 17289 18555 17323
rect 18555 17289 18564 17323
rect 18512 17280 18564 17289
rect 20260 17280 20312 17332
rect 21272 17280 21324 17332
rect 22100 17280 22152 17332
rect 30104 17323 30156 17332
rect 30104 17289 30113 17323
rect 30113 17289 30147 17323
rect 30147 17289 30156 17323
rect 30104 17280 30156 17289
rect 32496 17280 32548 17332
rect 33048 17280 33100 17332
rect 13728 17212 13780 17264
rect 15936 17255 15988 17264
rect 15936 17221 15945 17255
rect 15945 17221 15979 17255
rect 15979 17221 15988 17255
rect 15936 17212 15988 17221
rect 16304 17212 16356 17264
rect 2044 17119 2096 17128
rect 2044 17085 2053 17119
rect 2053 17085 2087 17119
rect 2087 17085 2096 17119
rect 2044 17076 2096 17085
rect 2780 17076 2832 17128
rect 2872 17119 2924 17128
rect 2872 17085 2881 17119
rect 2881 17085 2915 17119
rect 2915 17085 2924 17119
rect 15016 17144 15068 17196
rect 17132 17212 17184 17264
rect 16672 17144 16724 17196
rect 19432 17212 19484 17264
rect 20168 17212 20220 17264
rect 18052 17187 18104 17196
rect 18052 17153 18061 17187
rect 18061 17153 18095 17187
rect 18095 17153 18104 17187
rect 18052 17144 18104 17153
rect 18328 17187 18380 17196
rect 18328 17153 18337 17187
rect 18337 17153 18371 17187
rect 18371 17153 18380 17187
rect 18328 17144 18380 17153
rect 22008 17212 22060 17264
rect 29184 17212 29236 17264
rect 32772 17255 32824 17264
rect 32772 17221 32781 17255
rect 32781 17221 32815 17255
rect 32815 17221 32824 17255
rect 32772 17212 32824 17221
rect 34704 17212 34756 17264
rect 35440 17280 35492 17332
rect 44272 17323 44324 17332
rect 44272 17289 44281 17323
rect 44281 17289 44315 17323
rect 44315 17289 44324 17323
rect 44272 17280 44324 17289
rect 47860 17323 47912 17332
rect 47860 17289 47869 17323
rect 47869 17289 47903 17323
rect 47903 17289 47912 17323
rect 47860 17280 47912 17289
rect 36452 17212 36504 17264
rect 21272 17187 21324 17196
rect 21272 17153 21281 17187
rect 21281 17153 21315 17187
rect 21315 17153 21324 17187
rect 21272 17144 21324 17153
rect 21548 17144 21600 17196
rect 21732 17144 21784 17196
rect 23480 17144 23532 17196
rect 28540 17144 28592 17196
rect 33968 17144 34020 17196
rect 35348 17144 35400 17196
rect 40408 17144 40460 17196
rect 40960 17144 41012 17196
rect 41420 17144 41472 17196
rect 42984 17144 43036 17196
rect 44456 17187 44508 17196
rect 44456 17153 44465 17187
rect 44465 17153 44499 17187
rect 44499 17153 44508 17187
rect 44456 17144 44508 17153
rect 44548 17187 44600 17196
rect 44548 17153 44557 17187
rect 44557 17153 44591 17187
rect 44591 17153 44600 17187
rect 44548 17144 44600 17153
rect 47216 17144 47268 17196
rect 47676 17144 47728 17196
rect 2872 17076 2924 17085
rect 23020 17076 23072 17128
rect 16856 17008 16908 17060
rect 18144 17008 18196 17060
rect 20536 17008 20588 17060
rect 23112 17008 23164 17060
rect 23940 17076 23992 17128
rect 43444 17076 43496 17128
rect 43720 17076 43772 17128
rect 45284 17076 45336 17128
rect 41788 17008 41840 17060
rect 16304 16983 16356 16992
rect 16304 16949 16313 16983
rect 16313 16949 16347 16983
rect 16347 16949 16356 16983
rect 16304 16940 16356 16949
rect 17316 16983 17368 16992
rect 17316 16949 17325 16983
rect 17325 16949 17359 16983
rect 17359 16949 17368 16983
rect 17316 16940 17368 16949
rect 20996 16940 21048 16992
rect 23204 16983 23256 16992
rect 23204 16949 23213 16983
rect 23213 16949 23247 16983
rect 23247 16949 23256 16983
rect 23204 16940 23256 16949
rect 24032 16940 24084 16992
rect 40132 16940 40184 16992
rect 41420 16940 41472 16992
rect 43352 16940 43404 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 2044 16736 2096 16788
rect 17316 16736 17368 16788
rect 20628 16736 20680 16788
rect 18052 16668 18104 16720
rect 13728 16600 13780 16652
rect 2780 16532 2832 16584
rect 2964 16575 3016 16584
rect 2964 16541 2973 16575
rect 2973 16541 3007 16575
rect 3007 16541 3016 16575
rect 16028 16600 16080 16652
rect 16304 16600 16356 16652
rect 16580 16600 16632 16652
rect 2964 16532 3016 16541
rect 15016 16532 15068 16584
rect 15936 16532 15988 16584
rect 15844 16507 15896 16516
rect 15844 16473 15853 16507
rect 15853 16473 15887 16507
rect 15887 16473 15896 16507
rect 15844 16464 15896 16473
rect 20260 16464 20312 16516
rect 15200 16396 15252 16448
rect 20076 16396 20128 16448
rect 20444 16396 20496 16448
rect 23020 16736 23072 16788
rect 23388 16736 23440 16788
rect 31116 16736 31168 16788
rect 37556 16736 37608 16788
rect 21640 16575 21692 16584
rect 21640 16541 21649 16575
rect 21649 16541 21683 16575
rect 21683 16541 21692 16575
rect 21640 16532 21692 16541
rect 23480 16575 23532 16584
rect 21548 16507 21600 16516
rect 21548 16473 21557 16507
rect 21557 16473 21591 16507
rect 21591 16473 21600 16507
rect 21548 16464 21600 16473
rect 23480 16541 23489 16575
rect 23489 16541 23523 16575
rect 23523 16541 23532 16575
rect 23480 16532 23532 16541
rect 24860 16600 24912 16652
rect 25228 16575 25280 16584
rect 25228 16541 25237 16575
rect 25237 16541 25271 16575
rect 25271 16541 25280 16575
rect 25228 16532 25280 16541
rect 25596 16575 25648 16584
rect 25596 16541 25605 16575
rect 25605 16541 25639 16575
rect 25639 16541 25648 16575
rect 25596 16532 25648 16541
rect 29460 16532 29512 16584
rect 23296 16507 23348 16516
rect 23296 16473 23305 16507
rect 23305 16473 23339 16507
rect 23339 16473 23348 16507
rect 23296 16464 23348 16473
rect 30748 16532 30800 16584
rect 36084 16575 36136 16584
rect 36084 16541 36093 16575
rect 36093 16541 36127 16575
rect 36127 16541 36136 16575
rect 36084 16532 36136 16541
rect 37280 16600 37332 16652
rect 40224 16736 40276 16788
rect 43444 16779 43496 16788
rect 43444 16745 43453 16779
rect 43453 16745 43487 16779
rect 43487 16745 43496 16779
rect 43444 16736 43496 16745
rect 45468 16736 45520 16788
rect 40040 16600 40092 16652
rect 41512 16600 41564 16652
rect 40132 16532 40184 16584
rect 41788 16532 41840 16584
rect 42340 16600 42392 16652
rect 46112 16643 46164 16652
rect 25228 16396 25280 16448
rect 30564 16464 30616 16516
rect 31760 16464 31812 16516
rect 27804 16396 27856 16448
rect 34152 16396 34204 16448
rect 36176 16396 36228 16448
rect 36452 16396 36504 16448
rect 39948 16396 40000 16448
rect 40684 16464 40736 16516
rect 42248 16575 42300 16584
rect 42248 16541 42257 16575
rect 42257 16541 42291 16575
rect 42291 16541 42300 16575
rect 46112 16609 46121 16643
rect 46121 16609 46155 16643
rect 46155 16609 46164 16643
rect 46112 16600 46164 16609
rect 42248 16532 42300 16541
rect 43076 16575 43128 16584
rect 43076 16541 43085 16575
rect 43085 16541 43119 16575
rect 43119 16541 43128 16575
rect 43076 16532 43128 16541
rect 43260 16575 43312 16584
rect 43260 16541 43269 16575
rect 43269 16541 43303 16575
rect 43303 16541 43312 16575
rect 45192 16575 45244 16584
rect 43260 16532 43312 16541
rect 45192 16541 45201 16575
rect 45201 16541 45235 16575
rect 45235 16541 45244 16575
rect 45192 16532 45244 16541
rect 45468 16532 45520 16584
rect 46664 16464 46716 16516
rect 42800 16396 42852 16448
rect 47400 16396 47452 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 16304 16192 16356 16244
rect 20260 16235 20312 16244
rect 15200 16124 15252 16176
rect 14648 16099 14700 16108
rect 14648 16065 14657 16099
rect 14657 16065 14691 16099
rect 14691 16065 14700 16099
rect 14648 16056 14700 16065
rect 14832 16099 14884 16108
rect 14832 16065 14841 16099
rect 14841 16065 14875 16099
rect 14875 16065 14884 16099
rect 14832 16056 14884 16065
rect 16028 16056 16080 16108
rect 20260 16201 20269 16235
rect 20269 16201 20303 16235
rect 20303 16201 20312 16235
rect 20260 16192 20312 16201
rect 20536 16192 20588 16244
rect 20444 16099 20496 16108
rect 15844 16031 15896 16040
rect 15844 15997 15853 16031
rect 15853 15997 15887 16031
rect 15887 15997 15896 16031
rect 15844 15988 15896 15997
rect 20444 16065 20453 16099
rect 20453 16065 20487 16099
rect 20487 16065 20496 16099
rect 20444 16056 20496 16065
rect 21456 16056 21508 16108
rect 22836 16056 22888 16108
rect 23388 16056 23440 16108
rect 23480 16099 23532 16108
rect 23480 16065 23489 16099
rect 23489 16065 23523 16099
rect 23523 16065 23532 16099
rect 23480 16056 23532 16065
rect 23112 16031 23164 16040
rect 23112 15997 23121 16031
rect 23121 15997 23155 16031
rect 23155 15997 23164 16031
rect 24032 16031 24084 16040
rect 23112 15988 23164 15997
rect 24032 15997 24041 16031
rect 24041 15997 24075 16031
rect 24075 15997 24084 16031
rect 24032 15988 24084 15997
rect 23204 15920 23256 15972
rect 23296 15920 23348 15972
rect 26516 16192 26568 16244
rect 28632 16192 28684 16244
rect 36084 16192 36136 16244
rect 27712 16124 27764 16176
rect 25228 16099 25280 16108
rect 25228 16065 25237 16099
rect 25237 16065 25271 16099
rect 25271 16065 25280 16099
rect 25228 16056 25280 16065
rect 27344 16099 27396 16108
rect 27344 16065 27353 16099
rect 27353 16065 27387 16099
rect 27387 16065 27396 16099
rect 27620 16099 27672 16108
rect 27344 16056 27396 16065
rect 27620 16065 27629 16099
rect 27629 16065 27663 16099
rect 27663 16065 27672 16099
rect 27620 16056 27672 16065
rect 27804 16099 27856 16108
rect 27804 16065 27813 16099
rect 27813 16065 27847 16099
rect 27847 16065 27856 16099
rect 27804 16056 27856 16065
rect 28724 16124 28776 16176
rect 31760 16167 31812 16176
rect 31760 16133 31769 16167
rect 31769 16133 31803 16167
rect 31803 16133 31812 16167
rect 31760 16124 31812 16133
rect 28632 16099 28684 16108
rect 28632 16065 28666 16099
rect 28666 16065 28684 16099
rect 32312 16099 32364 16108
rect 28632 16056 28684 16065
rect 32312 16065 32321 16099
rect 32321 16065 32355 16099
rect 32355 16065 32364 16099
rect 32312 16056 32364 16065
rect 32404 16056 32456 16108
rect 37280 16124 37332 16176
rect 34244 16056 34296 16108
rect 36176 16099 36228 16108
rect 26516 16031 26568 16040
rect 26516 15997 26525 16031
rect 26525 15997 26559 16031
rect 26559 15997 26568 16031
rect 26516 15988 26568 15997
rect 36176 16065 36185 16099
rect 36185 16065 36219 16099
rect 36219 16065 36228 16099
rect 36176 16056 36228 16065
rect 37556 16235 37608 16244
rect 37556 16201 37565 16235
rect 37565 16201 37599 16235
rect 37599 16201 37608 16235
rect 37556 16192 37608 16201
rect 40316 16192 40368 16244
rect 42340 16192 42392 16244
rect 43076 16192 43128 16244
rect 37740 16099 37792 16108
rect 37740 16065 37749 16099
rect 37749 16065 37783 16099
rect 37783 16065 37792 16099
rect 37740 16056 37792 16065
rect 41052 16124 41104 16176
rect 45284 16192 45336 16244
rect 46664 16235 46716 16244
rect 40316 16056 40368 16108
rect 44456 16124 44508 16176
rect 46664 16201 46673 16235
rect 46673 16201 46707 16235
rect 46707 16201 46716 16235
rect 46664 16192 46716 16201
rect 42892 16056 42944 16108
rect 39948 16031 40000 16040
rect 16948 15895 17000 15904
rect 16948 15861 16957 15895
rect 16957 15861 16991 15895
rect 16991 15861 17000 15895
rect 16948 15852 17000 15861
rect 20812 15852 20864 15904
rect 25412 15895 25464 15904
rect 25412 15861 25421 15895
rect 25421 15861 25455 15895
rect 25455 15861 25464 15895
rect 25412 15852 25464 15861
rect 26148 15895 26200 15904
rect 26148 15861 26157 15895
rect 26157 15861 26191 15895
rect 26191 15861 26200 15895
rect 26148 15852 26200 15861
rect 26608 15852 26660 15904
rect 29460 15852 29512 15904
rect 30840 15852 30892 15904
rect 31760 15852 31812 15904
rect 33692 15895 33744 15904
rect 33692 15861 33701 15895
rect 33701 15861 33735 15895
rect 33735 15861 33744 15895
rect 33692 15852 33744 15861
rect 35440 15852 35492 15904
rect 39948 15997 39957 16031
rect 39957 15997 39991 16031
rect 39991 15997 40000 16031
rect 39948 15988 40000 15997
rect 44456 15988 44508 16040
rect 42248 15920 42300 15972
rect 45192 16056 45244 16108
rect 45376 16031 45428 16040
rect 45376 15997 45385 16031
rect 45385 15997 45419 16031
rect 45419 15997 45428 16031
rect 45376 15988 45428 15997
rect 45560 16056 45612 16108
rect 47400 16124 47452 16176
rect 46480 16099 46532 16108
rect 46480 16065 46489 16099
rect 46489 16065 46523 16099
rect 46523 16065 46532 16099
rect 46480 16056 46532 16065
rect 36360 15895 36412 15904
rect 36360 15861 36369 15895
rect 36369 15861 36403 15895
rect 36403 15861 36412 15895
rect 36360 15852 36412 15861
rect 40408 15895 40460 15904
rect 40408 15861 40417 15895
rect 40417 15861 40451 15895
rect 40451 15861 40460 15895
rect 40408 15852 40460 15861
rect 40960 15895 41012 15904
rect 40960 15861 40969 15895
rect 40969 15861 41003 15895
rect 41003 15861 41012 15895
rect 40960 15852 41012 15861
rect 44640 15895 44692 15904
rect 44640 15861 44649 15895
rect 44649 15861 44683 15895
rect 44683 15861 44692 15895
rect 44640 15852 44692 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 14280 15648 14332 15700
rect 14832 15648 14884 15700
rect 21456 15691 21508 15700
rect 21456 15657 21465 15691
rect 21465 15657 21499 15691
rect 21499 15657 21508 15691
rect 21456 15648 21508 15657
rect 23296 15691 23348 15700
rect 23296 15657 23305 15691
rect 23305 15657 23339 15691
rect 23339 15657 23348 15691
rect 23296 15648 23348 15657
rect 22836 15580 22888 15632
rect 27804 15648 27856 15700
rect 28632 15648 28684 15700
rect 28908 15648 28960 15700
rect 30012 15648 30064 15700
rect 32404 15648 32456 15700
rect 34244 15648 34296 15700
rect 36820 15648 36872 15700
rect 43260 15648 43312 15700
rect 44640 15648 44692 15700
rect 45376 15648 45428 15700
rect 6000 15444 6052 15496
rect 13268 15444 13320 15496
rect 14372 15444 14424 15496
rect 14648 15512 14700 15564
rect 16948 15512 17000 15564
rect 19432 15512 19484 15564
rect 20996 15555 21048 15564
rect 20996 15521 21005 15555
rect 21005 15521 21039 15555
rect 21039 15521 21048 15555
rect 20996 15512 21048 15521
rect 15844 15444 15896 15496
rect 18052 15487 18104 15496
rect 18052 15453 18061 15487
rect 18061 15453 18095 15487
rect 18095 15453 18104 15487
rect 18052 15444 18104 15453
rect 18236 15487 18288 15496
rect 18236 15453 18245 15487
rect 18245 15453 18279 15487
rect 18279 15453 18288 15487
rect 18236 15444 18288 15453
rect 20444 15487 20496 15496
rect 20444 15453 20453 15487
rect 20453 15453 20487 15487
rect 20487 15453 20496 15487
rect 20444 15444 20496 15453
rect 20812 15487 20864 15496
rect 20812 15453 20821 15487
rect 20821 15453 20855 15487
rect 20855 15453 20864 15487
rect 20812 15444 20864 15453
rect 21456 15487 21508 15496
rect 21456 15453 21465 15487
rect 21465 15453 21499 15487
rect 21499 15453 21508 15487
rect 21456 15444 21508 15453
rect 16028 15351 16080 15360
rect 16028 15317 16037 15351
rect 16037 15317 16071 15351
rect 16071 15317 16080 15351
rect 16028 15308 16080 15317
rect 17868 15351 17920 15360
rect 17868 15317 17877 15351
rect 17877 15317 17911 15351
rect 17911 15317 17920 15351
rect 17868 15308 17920 15317
rect 20260 15308 20312 15360
rect 23480 15444 23532 15496
rect 25596 15580 25648 15632
rect 25504 15512 25556 15564
rect 29000 15512 29052 15564
rect 30564 15580 30616 15632
rect 33692 15580 33744 15632
rect 30104 15512 30156 15564
rect 25596 15444 25648 15496
rect 28724 15444 28776 15496
rect 26148 15376 26200 15428
rect 30288 15444 30340 15496
rect 30840 15487 30892 15496
rect 30840 15453 30849 15487
rect 30849 15453 30883 15487
rect 30883 15453 30892 15487
rect 30840 15444 30892 15453
rect 31484 15487 31536 15496
rect 31484 15453 31493 15487
rect 31493 15453 31527 15487
rect 31527 15453 31536 15487
rect 31484 15444 31536 15453
rect 31576 15444 31628 15496
rect 31760 15487 31812 15496
rect 31760 15453 31769 15487
rect 31769 15453 31803 15487
rect 31803 15453 31812 15487
rect 35440 15512 35492 15564
rect 31760 15444 31812 15453
rect 30472 15376 30524 15428
rect 34152 15487 34204 15496
rect 33048 15376 33100 15428
rect 34152 15453 34161 15487
rect 34161 15453 34195 15487
rect 34195 15453 34204 15487
rect 34152 15444 34204 15453
rect 36176 15580 36228 15632
rect 40408 15580 40460 15632
rect 36360 15555 36412 15564
rect 36360 15521 36369 15555
rect 36369 15521 36403 15555
rect 36403 15521 36412 15555
rect 36360 15512 36412 15521
rect 36452 15555 36504 15564
rect 36452 15521 36461 15555
rect 36461 15521 36495 15555
rect 36495 15521 36504 15555
rect 36452 15512 36504 15521
rect 37556 15555 37608 15564
rect 37556 15521 37565 15555
rect 37565 15521 37599 15555
rect 37599 15521 37608 15555
rect 37556 15512 37608 15521
rect 42984 15512 43036 15564
rect 45560 15512 45612 15564
rect 38476 15487 38528 15496
rect 38476 15453 38485 15487
rect 38485 15453 38519 15487
rect 38519 15453 38528 15487
rect 38476 15444 38528 15453
rect 39856 15444 39908 15496
rect 40040 15487 40092 15496
rect 40040 15453 40049 15487
rect 40049 15453 40083 15487
rect 40083 15453 40092 15487
rect 40040 15444 40092 15453
rect 40132 15444 40184 15496
rect 42248 15444 42300 15496
rect 43260 15487 43312 15496
rect 43260 15453 43269 15487
rect 43269 15453 43303 15487
rect 43303 15453 43312 15487
rect 43260 15444 43312 15453
rect 43352 15487 43404 15496
rect 43352 15453 43361 15487
rect 43361 15453 43395 15487
rect 43395 15453 43404 15487
rect 43352 15444 43404 15453
rect 42340 15419 42392 15428
rect 42340 15385 42349 15419
rect 42349 15385 42383 15419
rect 42383 15385 42392 15419
rect 42340 15376 42392 15385
rect 44180 15419 44232 15428
rect 44180 15385 44207 15419
rect 44207 15385 44232 15419
rect 44180 15376 44232 15385
rect 44456 15444 44508 15496
rect 45284 15487 45336 15496
rect 45284 15453 45293 15487
rect 45293 15453 45327 15487
rect 45327 15453 45336 15487
rect 45284 15444 45336 15453
rect 48320 15444 48372 15496
rect 45008 15376 45060 15428
rect 45468 15419 45520 15428
rect 45468 15385 45477 15419
rect 45477 15385 45511 15419
rect 45511 15385 45520 15419
rect 45468 15376 45520 15385
rect 33324 15308 33376 15360
rect 36176 15351 36228 15360
rect 36176 15317 36185 15351
rect 36185 15317 36219 15351
rect 36219 15317 36228 15351
rect 36176 15308 36228 15317
rect 36820 15351 36872 15360
rect 36820 15317 36829 15351
rect 36829 15317 36863 15351
rect 36863 15317 36872 15351
rect 36820 15308 36872 15317
rect 40316 15308 40368 15360
rect 43536 15351 43588 15360
rect 43536 15317 43545 15351
rect 43545 15317 43579 15351
rect 43579 15317 43588 15351
rect 43536 15308 43588 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 14280 15147 14332 15156
rect 14280 15113 14289 15147
rect 14289 15113 14323 15147
rect 14323 15113 14332 15147
rect 14280 15104 14332 15113
rect 20444 15104 20496 15156
rect 21456 15104 21508 15156
rect 30472 15104 30524 15156
rect 31484 15104 31536 15156
rect 37740 15104 37792 15156
rect 3424 15036 3476 15088
rect 17868 15036 17920 15088
rect 25412 15036 25464 15088
rect 30656 15036 30708 15088
rect 6000 15011 6052 15020
rect 6000 14977 6009 15011
rect 6009 14977 6043 15011
rect 6043 14977 6052 15011
rect 6000 14968 6052 14977
rect 13268 14968 13320 15020
rect 14372 15011 14424 15020
rect 14372 14977 14381 15011
rect 14381 14977 14415 15011
rect 14415 14977 14424 15011
rect 14372 14968 14424 14977
rect 17500 15011 17552 15020
rect 17500 14977 17509 15011
rect 17509 14977 17543 15011
rect 17543 14977 17552 15011
rect 17500 14968 17552 14977
rect 19432 14968 19484 15020
rect 20168 14968 20220 15020
rect 20812 14968 20864 15020
rect 25780 14968 25832 15020
rect 26516 14968 26568 15020
rect 27436 14968 27488 15020
rect 28724 15011 28776 15020
rect 28724 14977 28733 15011
rect 28733 14977 28767 15011
rect 28767 14977 28776 15011
rect 28724 14968 28776 14977
rect 30472 14968 30524 15020
rect 30564 15011 30616 15020
rect 30564 14977 30573 15011
rect 30573 14977 30607 15011
rect 30607 14977 30616 15011
rect 43260 15036 43312 15088
rect 30564 14968 30616 14977
rect 30840 14968 30892 15020
rect 32312 15011 32364 15020
rect 32312 14977 32321 15011
rect 32321 14977 32355 15011
rect 32355 14977 32364 15011
rect 32312 14968 32364 14977
rect 32588 15011 32640 15020
rect 32588 14977 32622 15011
rect 32622 14977 32640 15011
rect 32588 14968 32640 14977
rect 36176 14968 36228 15020
rect 36360 14968 36412 15020
rect 36820 15011 36872 15020
rect 36820 14977 36829 15011
rect 36829 14977 36863 15011
rect 36863 14977 36872 15011
rect 36820 14968 36872 14977
rect 36912 14968 36964 15020
rect 5080 14900 5132 14952
rect 22652 14900 22704 14952
rect 26608 14900 26660 14952
rect 37556 14943 37608 14952
rect 25596 14832 25648 14884
rect 33968 14832 34020 14884
rect 35440 14832 35492 14884
rect 37556 14909 37565 14943
rect 37565 14909 37599 14943
rect 37599 14909 37608 14943
rect 37556 14900 37608 14909
rect 40408 14943 40460 14952
rect 40408 14909 40417 14943
rect 40417 14909 40451 14943
rect 40451 14909 40460 14943
rect 40408 14900 40460 14909
rect 42892 15011 42944 15020
rect 42892 14977 42901 15011
rect 42901 14977 42935 15011
rect 42935 14977 42944 15011
rect 42892 14968 42944 14977
rect 43536 14968 43588 15020
rect 45008 15011 45060 15020
rect 45008 14977 45017 15011
rect 45017 14977 45051 15011
rect 45051 14977 45060 15011
rect 45008 14968 45060 14977
rect 47492 14968 47544 15020
rect 40960 14900 41012 14952
rect 41144 14875 41196 14884
rect 3424 14764 3476 14816
rect 18788 14764 18840 14816
rect 20996 14764 21048 14816
rect 26240 14764 26292 14816
rect 33876 14764 33928 14816
rect 41144 14841 41153 14875
rect 41153 14841 41187 14875
rect 41187 14841 41196 14875
rect 41144 14832 41196 14841
rect 43352 14900 43404 14952
rect 44272 14943 44324 14952
rect 44272 14909 44281 14943
rect 44281 14909 44315 14943
rect 44315 14909 44324 14943
rect 44272 14900 44324 14909
rect 44364 14943 44416 14952
rect 44364 14909 44373 14943
rect 44373 14909 44407 14943
rect 44407 14909 44416 14943
rect 44364 14900 44416 14909
rect 40868 14764 40920 14816
rect 43720 14807 43772 14816
rect 43720 14773 43729 14807
rect 43729 14773 43763 14807
rect 43763 14773 43772 14807
rect 43720 14764 43772 14773
rect 45468 14832 45520 14884
rect 44364 14764 44416 14816
rect 48136 14764 48188 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 5080 14603 5132 14612
rect 5080 14569 5089 14603
rect 5089 14569 5123 14603
rect 5123 14569 5132 14603
rect 5080 14560 5132 14569
rect 18052 14560 18104 14612
rect 20168 14603 20220 14612
rect 20168 14569 20177 14603
rect 20177 14569 20211 14603
rect 20211 14569 20220 14603
rect 20168 14560 20220 14569
rect 21088 14560 21140 14612
rect 30472 14560 30524 14612
rect 32588 14603 32640 14612
rect 32588 14569 32597 14603
rect 32597 14569 32631 14603
rect 32631 14569 32640 14603
rect 32588 14560 32640 14569
rect 3424 14467 3476 14476
rect 3424 14433 3433 14467
rect 3433 14433 3467 14467
rect 3467 14433 3476 14467
rect 3424 14424 3476 14433
rect 14372 14424 14424 14476
rect 14924 14424 14976 14476
rect 1584 14399 1636 14408
rect 1584 14365 1593 14399
rect 1593 14365 1627 14399
rect 1627 14365 1636 14399
rect 1584 14356 1636 14365
rect 5816 14356 5868 14408
rect 16028 14424 16080 14476
rect 20444 14492 20496 14544
rect 30012 14492 30064 14544
rect 25688 14424 25740 14476
rect 2412 14288 2464 14340
rect 13452 14220 13504 14272
rect 17500 14356 17552 14408
rect 18328 14399 18380 14408
rect 18328 14365 18337 14399
rect 18337 14365 18371 14399
rect 18371 14365 18380 14399
rect 18328 14356 18380 14365
rect 18512 14356 18564 14408
rect 18788 14399 18840 14408
rect 18788 14365 18797 14399
rect 18797 14365 18831 14399
rect 18831 14365 18840 14399
rect 19984 14399 20036 14408
rect 18788 14356 18840 14365
rect 19984 14365 19993 14399
rect 19993 14365 20027 14399
rect 20027 14365 20036 14399
rect 19984 14356 20036 14365
rect 21088 14399 21140 14408
rect 21088 14365 21097 14399
rect 21097 14365 21131 14399
rect 21131 14365 21140 14399
rect 21088 14356 21140 14365
rect 21364 14399 21416 14408
rect 21364 14365 21373 14399
rect 21373 14365 21407 14399
rect 21407 14365 21416 14399
rect 21364 14356 21416 14365
rect 26240 14356 26292 14408
rect 28724 14356 28776 14408
rect 20076 14288 20128 14340
rect 30104 14356 30156 14408
rect 30288 14356 30340 14408
rect 33600 14560 33652 14612
rect 35440 14603 35492 14612
rect 34152 14492 34204 14544
rect 33876 14424 33928 14476
rect 33324 14399 33376 14408
rect 20352 14220 20404 14272
rect 20904 14263 20956 14272
rect 20904 14229 20913 14263
rect 20913 14229 20947 14263
rect 20947 14229 20956 14263
rect 20904 14220 20956 14229
rect 25504 14263 25556 14272
rect 25504 14229 25513 14263
rect 25513 14229 25547 14263
rect 25547 14229 25556 14263
rect 25504 14220 25556 14229
rect 30380 14288 30432 14340
rect 29920 14220 29972 14272
rect 33324 14365 33333 14399
rect 33333 14365 33367 14399
rect 33367 14365 33376 14399
rect 33324 14356 33376 14365
rect 33416 14356 33468 14408
rect 33968 14399 34020 14408
rect 33968 14365 33977 14399
rect 33977 14365 34011 14399
rect 34011 14365 34020 14399
rect 33968 14356 34020 14365
rect 34980 14399 35032 14408
rect 34980 14365 34989 14399
rect 34989 14365 35023 14399
rect 35023 14365 35032 14399
rect 34980 14356 35032 14365
rect 35440 14569 35449 14603
rect 35449 14569 35483 14603
rect 35483 14569 35492 14603
rect 35440 14560 35492 14569
rect 40960 14560 41012 14612
rect 44364 14560 44416 14612
rect 36360 14492 36412 14544
rect 36636 14467 36688 14476
rect 36636 14433 36645 14467
rect 36645 14433 36679 14467
rect 36679 14433 36688 14467
rect 36636 14424 36688 14433
rect 46848 14467 46900 14476
rect 46848 14433 46857 14467
rect 46857 14433 46891 14467
rect 46891 14433 46900 14467
rect 46848 14424 46900 14433
rect 48136 14467 48188 14476
rect 48136 14433 48145 14467
rect 48145 14433 48179 14467
rect 48179 14433 48188 14467
rect 48136 14424 48188 14433
rect 48320 14467 48372 14476
rect 48320 14433 48329 14467
rect 48329 14433 48363 14467
rect 48363 14433 48372 14467
rect 48320 14424 48372 14433
rect 36452 14356 36504 14408
rect 40224 14399 40276 14408
rect 40224 14365 40233 14399
rect 40233 14365 40267 14399
rect 40267 14365 40276 14399
rect 40224 14356 40276 14365
rect 46112 14356 46164 14408
rect 40500 14331 40552 14340
rect 40500 14297 40534 14331
rect 40534 14297 40552 14331
rect 40500 14288 40552 14297
rect 43720 14288 43772 14340
rect 33048 14220 33100 14272
rect 37648 14220 37700 14272
rect 40684 14220 40736 14272
rect 44272 14220 44324 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 2412 14059 2464 14068
rect 2412 14025 2421 14059
rect 2421 14025 2455 14059
rect 2455 14025 2464 14059
rect 2412 14016 2464 14025
rect 14372 14016 14424 14068
rect 19432 14016 19484 14068
rect 20076 14016 20128 14068
rect 21180 14016 21232 14068
rect 25780 14059 25832 14068
rect 2504 13923 2556 13932
rect 2504 13889 2513 13923
rect 2513 13889 2547 13923
rect 2547 13889 2556 13923
rect 2504 13880 2556 13889
rect 5172 13880 5224 13932
rect 12256 13880 12308 13932
rect 16212 13948 16264 14000
rect 13452 13923 13504 13932
rect 13452 13889 13486 13923
rect 13486 13889 13504 13923
rect 13452 13880 13504 13889
rect 19892 13948 19944 14000
rect 19984 13880 20036 13932
rect 19340 13812 19392 13864
rect 20628 13948 20680 14000
rect 22652 13948 22704 14000
rect 20904 13880 20956 13932
rect 23388 13923 23440 13932
rect 23388 13889 23397 13923
rect 23397 13889 23431 13923
rect 23431 13889 23440 13923
rect 23388 13880 23440 13889
rect 25780 14025 25789 14059
rect 25789 14025 25823 14059
rect 25823 14025 25832 14059
rect 25780 14016 25832 14025
rect 34980 14016 35032 14068
rect 40500 14059 40552 14068
rect 40500 14025 40509 14059
rect 40509 14025 40543 14059
rect 40543 14025 40552 14059
rect 40500 14016 40552 14025
rect 25504 13948 25556 14000
rect 34152 13991 34204 14000
rect 23664 13855 23716 13864
rect 23664 13821 23673 13855
rect 23673 13821 23707 13855
rect 23707 13821 23716 13855
rect 23664 13812 23716 13821
rect 25688 13880 25740 13932
rect 26240 13923 26292 13932
rect 26240 13889 26249 13923
rect 26249 13889 26283 13923
rect 26283 13889 26292 13923
rect 26240 13880 26292 13889
rect 34152 13957 34161 13991
rect 34161 13957 34195 13991
rect 34195 13957 34204 13991
rect 34152 13948 34204 13957
rect 36176 13948 36228 14000
rect 40868 13991 40920 14000
rect 40868 13957 40877 13991
rect 40877 13957 40911 13991
rect 40911 13957 40920 13991
rect 40868 13948 40920 13957
rect 30012 13923 30064 13932
rect 30012 13889 30021 13923
rect 30021 13889 30055 13923
rect 30055 13889 30064 13923
rect 30012 13880 30064 13889
rect 30196 13923 30248 13932
rect 30196 13889 30205 13923
rect 30205 13889 30239 13923
rect 30239 13889 30248 13923
rect 30196 13880 30248 13889
rect 33048 13923 33100 13932
rect 33048 13889 33057 13923
rect 33057 13889 33091 13923
rect 33091 13889 33100 13923
rect 33048 13880 33100 13889
rect 33416 13880 33468 13932
rect 33784 13923 33836 13932
rect 33784 13889 33793 13923
rect 33793 13889 33827 13923
rect 33827 13889 33836 13923
rect 33784 13880 33836 13889
rect 40684 13923 40736 13932
rect 40684 13889 40693 13923
rect 40693 13889 40727 13923
rect 40727 13889 40736 13923
rect 40684 13880 40736 13889
rect 40960 13880 41012 13932
rect 42984 13880 43036 13932
rect 26700 13812 26752 13864
rect 30564 13812 30616 13864
rect 48320 13812 48372 13864
rect 34980 13744 35032 13796
rect 35808 13744 35860 13796
rect 21640 13676 21692 13728
rect 23204 13719 23256 13728
rect 23204 13685 23213 13719
rect 23213 13685 23247 13719
rect 23247 13685 23256 13719
rect 23204 13676 23256 13685
rect 30380 13719 30432 13728
rect 30380 13685 30389 13719
rect 30389 13685 30423 13719
rect 30423 13685 30432 13719
rect 30380 13676 30432 13685
rect 36360 13719 36412 13728
rect 36360 13685 36369 13719
rect 36369 13685 36403 13719
rect 36403 13685 36412 13719
rect 36360 13676 36412 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 21088 13472 21140 13524
rect 26608 13472 26660 13524
rect 27344 13515 27396 13524
rect 27344 13481 27353 13515
rect 27353 13481 27387 13515
rect 27387 13481 27396 13515
rect 27344 13472 27396 13481
rect 30012 13472 30064 13524
rect 33416 13472 33468 13524
rect 36912 13472 36964 13524
rect 19984 13404 20036 13456
rect 30472 13404 30524 13456
rect 30748 13404 30800 13456
rect 31024 13404 31076 13456
rect 33324 13404 33376 13456
rect 37188 13404 37240 13456
rect 18328 13336 18380 13388
rect 22652 13379 22704 13388
rect 22652 13345 22661 13379
rect 22661 13345 22695 13379
rect 22695 13345 22704 13379
rect 22652 13336 22704 13345
rect 16212 13311 16264 13320
rect 16212 13277 16221 13311
rect 16221 13277 16255 13311
rect 16255 13277 16264 13311
rect 16212 13268 16264 13277
rect 18512 13311 18564 13320
rect 18512 13277 18521 13311
rect 18521 13277 18555 13311
rect 18555 13277 18564 13311
rect 18512 13268 18564 13277
rect 19892 13311 19944 13320
rect 17040 13200 17092 13252
rect 18328 13200 18380 13252
rect 19892 13277 19901 13311
rect 19901 13277 19935 13311
rect 19935 13277 19944 13311
rect 19892 13268 19944 13277
rect 20076 13268 20128 13320
rect 20260 13268 20312 13320
rect 21180 13311 21232 13320
rect 21180 13277 21189 13311
rect 21189 13277 21223 13311
rect 21223 13277 21232 13311
rect 21180 13268 21232 13277
rect 21640 13311 21692 13320
rect 21640 13277 21649 13311
rect 21649 13277 21683 13311
rect 21683 13277 21692 13311
rect 21640 13268 21692 13277
rect 23204 13268 23256 13320
rect 26056 13311 26108 13320
rect 26056 13277 26065 13311
rect 26065 13277 26099 13311
rect 26099 13277 26108 13311
rect 26056 13268 26108 13277
rect 27620 13336 27672 13388
rect 28724 13336 28776 13388
rect 30012 13336 30064 13388
rect 33140 13336 33192 13388
rect 36452 13336 36504 13388
rect 37648 13379 37700 13388
rect 37648 13345 37657 13379
rect 37657 13345 37691 13379
rect 37691 13345 37700 13379
rect 37648 13336 37700 13345
rect 38476 13336 38528 13388
rect 46848 13379 46900 13388
rect 46848 13345 46857 13379
rect 46857 13345 46891 13379
rect 46891 13345 46900 13379
rect 46848 13336 46900 13345
rect 48320 13379 48372 13388
rect 48320 13345 48329 13379
rect 48329 13345 48363 13379
rect 48363 13345 48372 13379
rect 48320 13336 48372 13345
rect 26608 13268 26660 13320
rect 28356 13311 28408 13320
rect 22100 13200 22152 13252
rect 23756 13200 23808 13252
rect 25872 13200 25924 13252
rect 28356 13277 28365 13311
rect 28365 13277 28399 13311
rect 28399 13277 28408 13311
rect 28356 13268 28408 13277
rect 28632 13311 28684 13320
rect 28632 13277 28641 13311
rect 28641 13277 28675 13311
rect 28675 13277 28684 13311
rect 29920 13311 29972 13320
rect 28632 13268 28684 13277
rect 29920 13277 29929 13311
rect 29929 13277 29963 13311
rect 29963 13277 29972 13311
rect 29920 13268 29972 13277
rect 28540 13200 28592 13252
rect 29644 13200 29696 13252
rect 30472 13268 30524 13320
rect 33416 13268 33468 13320
rect 35808 13268 35860 13320
rect 36728 13268 36780 13320
rect 37832 13311 37884 13320
rect 37832 13277 37841 13311
rect 37841 13277 37875 13311
rect 37875 13277 37884 13311
rect 37832 13268 37884 13277
rect 30656 13200 30708 13252
rect 36176 13200 36228 13252
rect 47860 13200 47912 13252
rect 18052 13175 18104 13184
rect 18052 13141 18061 13175
rect 18061 13141 18095 13175
rect 18095 13141 18104 13175
rect 18052 13132 18104 13141
rect 24032 13175 24084 13184
rect 24032 13141 24041 13175
rect 24041 13141 24075 13175
rect 24075 13141 24084 13175
rect 24032 13132 24084 13141
rect 26424 13132 26476 13184
rect 27988 13132 28040 13184
rect 36820 13132 36872 13184
rect 37372 13175 37424 13184
rect 37372 13141 37381 13175
rect 37381 13141 37415 13175
rect 37415 13141 37424 13175
rect 37372 13132 37424 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 17040 12971 17092 12980
rect 17040 12937 17049 12971
rect 17049 12937 17083 12971
rect 17083 12937 17092 12971
rect 17040 12928 17092 12937
rect 21640 12928 21692 12980
rect 23388 12928 23440 12980
rect 25320 12928 25372 12980
rect 26056 12928 26108 12980
rect 26608 12928 26660 12980
rect 33784 12928 33836 12980
rect 36728 12971 36780 12980
rect 18052 12792 18104 12844
rect 4712 12724 4764 12776
rect 21364 12860 21416 12912
rect 20444 12792 20496 12844
rect 20260 12724 20312 12776
rect 21180 12792 21232 12844
rect 23756 12835 23808 12844
rect 23756 12801 23765 12835
rect 23765 12801 23799 12835
rect 23799 12801 23808 12835
rect 23756 12792 23808 12801
rect 24032 12792 24084 12844
rect 26332 12835 26384 12844
rect 28724 12860 28776 12912
rect 30380 12860 30432 12912
rect 33324 12860 33376 12912
rect 36728 12937 36737 12971
rect 36737 12937 36771 12971
rect 36771 12937 36780 12971
rect 36728 12928 36780 12937
rect 37004 12928 37056 12980
rect 42340 12928 42392 12980
rect 47860 12971 47912 12980
rect 47860 12937 47869 12971
rect 47869 12937 47903 12971
rect 47903 12937 47912 12971
rect 47860 12928 47912 12937
rect 37372 12860 37424 12912
rect 26332 12801 26350 12835
rect 26350 12801 26384 12835
rect 26332 12792 26384 12801
rect 27988 12835 28040 12844
rect 27988 12801 28022 12835
rect 28022 12801 28040 12835
rect 27988 12792 28040 12801
rect 29828 12792 29880 12844
rect 30012 12835 30064 12844
rect 30012 12801 30021 12835
rect 30021 12801 30055 12835
rect 30055 12801 30064 12835
rect 30012 12792 30064 12801
rect 33232 12835 33284 12844
rect 33232 12801 33241 12835
rect 33241 12801 33275 12835
rect 33275 12801 33284 12835
rect 33232 12792 33284 12801
rect 23296 12724 23348 12776
rect 18236 12656 18288 12708
rect 34612 12792 34664 12844
rect 34796 12724 34848 12776
rect 35808 12656 35860 12708
rect 36636 12792 36688 12844
rect 40224 12792 40276 12844
rect 46756 12792 46808 12844
rect 47492 12792 47544 12844
rect 47676 12792 47728 12844
rect 36452 12767 36504 12776
rect 36452 12733 36461 12767
rect 36461 12733 36495 12767
rect 36495 12733 36504 12767
rect 36452 12724 36504 12733
rect 37556 12656 37608 12708
rect 17960 12588 18012 12640
rect 29092 12631 29144 12640
rect 29092 12597 29101 12631
rect 29101 12597 29135 12631
rect 29135 12597 29144 12631
rect 29092 12588 29144 12597
rect 31392 12631 31444 12640
rect 31392 12597 31401 12631
rect 31401 12597 31435 12631
rect 31435 12597 31444 12631
rect 31392 12588 31444 12597
rect 35440 12588 35492 12640
rect 36176 12588 36228 12640
rect 36360 12631 36412 12640
rect 36360 12597 36369 12631
rect 36369 12597 36403 12631
rect 36403 12597 36412 12631
rect 36360 12588 36412 12597
rect 37464 12588 37516 12640
rect 46664 12588 46716 12640
rect 47032 12631 47084 12640
rect 47032 12597 47041 12631
rect 47041 12597 47075 12631
rect 47075 12597 47084 12631
rect 47032 12588 47084 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 17500 12384 17552 12436
rect 20536 12384 20588 12436
rect 26332 12384 26384 12436
rect 26608 12384 26660 12436
rect 28356 12384 28408 12436
rect 30196 12427 30248 12436
rect 30196 12393 30205 12427
rect 30205 12393 30239 12427
rect 30239 12393 30248 12427
rect 30196 12384 30248 12393
rect 34704 12384 34756 12436
rect 35900 12384 35952 12436
rect 36360 12384 36412 12436
rect 37832 12384 37884 12436
rect 20260 12359 20312 12368
rect 20260 12325 20269 12359
rect 20269 12325 20303 12359
rect 20303 12325 20312 12359
rect 20260 12316 20312 12325
rect 29092 12316 29144 12368
rect 19984 12291 20036 12300
rect 19984 12257 19993 12291
rect 19993 12257 20027 12291
rect 20027 12257 20036 12291
rect 19984 12248 20036 12257
rect 23296 12248 23348 12300
rect 23848 12248 23900 12300
rect 26608 12291 26660 12300
rect 26608 12257 26617 12291
rect 26617 12257 26651 12291
rect 26651 12257 26660 12291
rect 26608 12248 26660 12257
rect 30564 12248 30616 12300
rect 33784 12248 33836 12300
rect 2596 12180 2648 12232
rect 17960 12180 18012 12232
rect 18328 12180 18380 12232
rect 24032 12180 24084 12232
rect 25872 12180 25924 12232
rect 26424 12180 26476 12232
rect 29092 12223 29144 12232
rect 19984 12112 20036 12164
rect 22928 12112 22980 12164
rect 2228 12044 2280 12096
rect 17040 12044 17092 12096
rect 17316 12087 17368 12096
rect 17316 12053 17325 12087
rect 17325 12053 17359 12087
rect 17359 12053 17368 12087
rect 17316 12044 17368 12053
rect 18236 12087 18288 12096
rect 18236 12053 18245 12087
rect 18245 12053 18279 12087
rect 18279 12053 18288 12087
rect 18236 12044 18288 12053
rect 18972 12044 19024 12096
rect 20812 12044 20864 12096
rect 25596 12087 25648 12096
rect 25596 12053 25605 12087
rect 25605 12053 25639 12087
rect 25639 12053 25648 12087
rect 25596 12044 25648 12053
rect 29092 12189 29101 12223
rect 29101 12189 29135 12223
rect 29135 12189 29144 12223
rect 29092 12180 29144 12189
rect 30288 12180 30340 12232
rect 30104 12112 30156 12164
rect 31392 12180 31444 12232
rect 35992 12248 36044 12300
rect 37004 12248 37056 12300
rect 35348 12180 35400 12232
rect 35440 12180 35492 12232
rect 34704 12112 34756 12164
rect 30288 12044 30340 12096
rect 33508 12044 33560 12096
rect 35532 12044 35584 12096
rect 36360 12223 36412 12232
rect 36360 12189 36369 12223
rect 36369 12189 36403 12223
rect 36403 12189 36412 12223
rect 36360 12180 36412 12189
rect 37464 12223 37516 12232
rect 37464 12189 37473 12223
rect 37473 12189 37507 12223
rect 37507 12189 37516 12223
rect 37464 12180 37516 12189
rect 39304 12248 39356 12300
rect 47032 12316 47084 12368
rect 46664 12291 46716 12300
rect 46664 12257 46673 12291
rect 46673 12257 46707 12291
rect 46707 12257 46716 12291
rect 46664 12248 46716 12257
rect 48228 12291 48280 12300
rect 48228 12257 48237 12291
rect 48237 12257 48271 12291
rect 48271 12257 48280 12291
rect 48228 12248 48280 12257
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 19432 11840 19484 11892
rect 20352 11840 20404 11892
rect 22284 11883 22336 11892
rect 2228 11815 2280 11824
rect 2228 11781 2237 11815
rect 2237 11781 2271 11815
rect 2271 11781 2280 11815
rect 2228 11772 2280 11781
rect 18972 11815 19024 11824
rect 18972 11781 18981 11815
rect 18981 11781 19015 11815
rect 19015 11781 19024 11815
rect 18972 11772 19024 11781
rect 17040 11747 17092 11756
rect 17040 11713 17049 11747
rect 17049 11713 17083 11747
rect 17083 11713 17092 11747
rect 17040 11704 17092 11713
rect 2044 11679 2096 11688
rect 2044 11645 2053 11679
rect 2053 11645 2087 11679
rect 2087 11645 2096 11679
rect 2044 11636 2096 11645
rect 2780 11679 2832 11688
rect 2780 11645 2789 11679
rect 2789 11645 2823 11679
rect 2823 11645 2832 11679
rect 2780 11636 2832 11645
rect 18236 11568 18288 11620
rect 19984 11704 20036 11756
rect 21916 11772 21968 11824
rect 22284 11849 22293 11883
rect 22293 11849 22327 11883
rect 22327 11849 22336 11883
rect 22284 11840 22336 11849
rect 25320 11883 25372 11892
rect 25320 11849 25329 11883
rect 25329 11849 25363 11883
rect 25363 11849 25372 11883
rect 25320 11840 25372 11849
rect 29000 11840 29052 11892
rect 31024 11840 31076 11892
rect 34796 11840 34848 11892
rect 35440 11772 35492 11824
rect 22560 11747 22612 11756
rect 22560 11713 22569 11747
rect 22569 11713 22603 11747
rect 22603 11713 22612 11747
rect 22560 11704 22612 11713
rect 23848 11704 23900 11756
rect 28540 11747 28592 11756
rect 21548 11636 21600 11688
rect 25228 11636 25280 11688
rect 28540 11713 28549 11747
rect 28549 11713 28583 11747
rect 28583 11713 28592 11747
rect 28540 11704 28592 11713
rect 30656 11747 30708 11756
rect 30656 11713 30665 11747
rect 30665 11713 30699 11747
rect 30699 11713 30708 11747
rect 30656 11704 30708 11713
rect 29644 11636 29696 11688
rect 31024 11704 31076 11756
rect 31576 11568 31628 11620
rect 33140 11704 33192 11756
rect 33508 11747 33560 11756
rect 33508 11713 33517 11747
rect 33517 11713 33551 11747
rect 33551 11713 33560 11747
rect 33508 11704 33560 11713
rect 34704 11747 34756 11756
rect 34704 11713 34713 11747
rect 34713 11713 34747 11747
rect 34747 11713 34756 11747
rect 34704 11704 34756 11713
rect 35532 11747 35584 11756
rect 35532 11713 35541 11747
rect 35541 11713 35575 11747
rect 35575 11713 35584 11747
rect 35532 11704 35584 11713
rect 35992 11704 36044 11756
rect 36912 11840 36964 11892
rect 37556 11883 37608 11892
rect 37556 11849 37565 11883
rect 37565 11849 37599 11883
rect 37599 11849 37608 11883
rect 37556 11840 37608 11849
rect 36268 11747 36320 11756
rect 36268 11713 36277 11747
rect 36277 11713 36311 11747
rect 36311 11713 36320 11747
rect 36268 11704 36320 11713
rect 36636 11704 36688 11756
rect 37648 11747 37700 11756
rect 33048 11636 33100 11688
rect 37648 11713 37657 11747
rect 37657 11713 37691 11747
rect 37691 11713 37700 11747
rect 37648 11704 37700 11713
rect 35348 11611 35400 11620
rect 35348 11577 35357 11611
rect 35357 11577 35391 11611
rect 35391 11577 35400 11611
rect 35348 11568 35400 11577
rect 16212 11500 16264 11552
rect 22468 11500 22520 11552
rect 24952 11543 25004 11552
rect 24952 11509 24961 11543
rect 24961 11509 24995 11543
rect 24995 11509 25004 11543
rect 24952 11500 25004 11509
rect 32312 11543 32364 11552
rect 32312 11509 32321 11543
rect 32321 11509 32355 11543
rect 32355 11509 32364 11543
rect 32312 11500 32364 11509
rect 33416 11500 33468 11552
rect 34612 11500 34664 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 2044 11339 2096 11348
rect 2044 11305 2053 11339
rect 2053 11305 2087 11339
rect 2087 11305 2096 11339
rect 2044 11296 2096 11305
rect 17316 11339 17368 11348
rect 17316 11305 17325 11339
rect 17325 11305 17359 11339
rect 17359 11305 17368 11339
rect 17316 11296 17368 11305
rect 22928 11339 22980 11348
rect 22928 11305 22937 11339
rect 22937 11305 22971 11339
rect 22971 11305 22980 11339
rect 22928 11296 22980 11305
rect 26516 11339 26568 11348
rect 18144 11271 18196 11280
rect 18144 11237 18153 11271
rect 18153 11237 18187 11271
rect 18187 11237 18196 11271
rect 26516 11305 26525 11339
rect 26525 11305 26559 11339
rect 26559 11305 26568 11339
rect 26516 11296 26568 11305
rect 33048 11339 33100 11348
rect 33048 11305 33057 11339
rect 33057 11305 33091 11339
rect 33091 11305 33100 11339
rect 33048 11296 33100 11305
rect 34612 11296 34664 11348
rect 35532 11296 35584 11348
rect 18144 11228 18196 11237
rect 22468 11203 22520 11212
rect 22468 11169 22477 11203
rect 22477 11169 22511 11203
rect 22511 11169 22520 11203
rect 22468 11160 22520 11169
rect 25136 11203 25188 11212
rect 25136 11169 25145 11203
rect 25145 11169 25179 11203
rect 25179 11169 25188 11203
rect 25136 11160 25188 11169
rect 26608 11160 26660 11212
rect 17316 11092 17368 11144
rect 17960 11135 18012 11144
rect 17960 11101 17969 11135
rect 17969 11101 18003 11135
rect 18003 11101 18012 11135
rect 17960 11092 18012 11101
rect 18236 11135 18288 11144
rect 18236 11101 18245 11135
rect 18245 11101 18279 11135
rect 18279 11101 18288 11135
rect 18236 11092 18288 11101
rect 19984 11092 20036 11144
rect 22376 11092 22428 11144
rect 23388 11092 23440 11144
rect 24952 11135 25004 11144
rect 24952 11101 24961 11135
rect 24961 11101 24995 11135
rect 24995 11101 25004 11135
rect 24952 11092 25004 11101
rect 26700 11135 26752 11144
rect 26700 11101 26709 11135
rect 26709 11101 26743 11135
rect 26743 11101 26752 11135
rect 26700 11092 26752 11101
rect 16212 11067 16264 11076
rect 16212 11033 16246 11067
rect 16246 11033 16264 11067
rect 16212 11024 16264 11033
rect 16304 11024 16356 11076
rect 23664 11024 23716 11076
rect 28632 11092 28684 11144
rect 29644 11160 29696 11212
rect 29000 11135 29052 11144
rect 29000 11101 29009 11135
rect 29009 11101 29043 11135
rect 29043 11101 29052 11135
rect 29000 11092 29052 11101
rect 29092 11092 29144 11144
rect 29828 11092 29880 11144
rect 31668 11135 31720 11144
rect 31668 11101 31677 11135
rect 31677 11101 31711 11135
rect 31711 11101 31720 11135
rect 31668 11092 31720 11101
rect 32312 11092 32364 11144
rect 36268 11296 36320 11348
rect 34704 11160 34756 11212
rect 28264 11024 28316 11076
rect 29552 11024 29604 11076
rect 37648 11228 37700 11280
rect 37464 11024 37516 11076
rect 17776 10999 17828 11008
rect 17776 10965 17785 10999
rect 17785 10965 17819 10999
rect 17819 10965 17828 10999
rect 17776 10956 17828 10965
rect 19432 10956 19484 11008
rect 24676 10956 24728 11008
rect 25044 10999 25096 11008
rect 25044 10965 25053 10999
rect 25053 10965 25087 10999
rect 25087 10965 25096 10999
rect 25044 10956 25096 10965
rect 29736 10956 29788 11008
rect 31116 10999 31168 11008
rect 31116 10965 31125 10999
rect 31125 10965 31159 10999
rect 31159 10965 31168 10999
rect 31116 10956 31168 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 17776 10684 17828 10736
rect 4620 10616 4672 10668
rect 17316 10659 17368 10668
rect 17316 10625 17325 10659
rect 17325 10625 17359 10659
rect 17359 10625 17368 10659
rect 17316 10616 17368 10625
rect 19340 10752 19392 10804
rect 22560 10752 22612 10804
rect 19432 10727 19484 10736
rect 19432 10693 19466 10727
rect 19466 10693 19484 10727
rect 19432 10684 19484 10693
rect 21548 10684 21600 10736
rect 22284 10727 22336 10736
rect 20720 10616 20772 10668
rect 21456 10659 21508 10668
rect 21456 10625 21465 10659
rect 21465 10625 21499 10659
rect 21499 10625 21508 10659
rect 21456 10616 21508 10625
rect 21824 10616 21876 10668
rect 22284 10693 22293 10727
rect 22293 10693 22327 10727
rect 22327 10693 22336 10727
rect 22284 10684 22336 10693
rect 22192 10616 22244 10668
rect 22744 10616 22796 10668
rect 23388 10659 23440 10668
rect 23388 10625 23397 10659
rect 23397 10625 23431 10659
rect 23431 10625 23440 10659
rect 23388 10616 23440 10625
rect 24032 10659 24084 10668
rect 24032 10625 24041 10659
rect 24041 10625 24075 10659
rect 24075 10625 24084 10659
rect 24032 10616 24084 10625
rect 25044 10752 25096 10804
rect 29552 10795 29604 10804
rect 29552 10761 29561 10795
rect 29561 10761 29595 10795
rect 29595 10761 29604 10795
rect 29552 10752 29604 10761
rect 34704 10752 34756 10804
rect 24860 10616 24912 10668
rect 28264 10659 28316 10668
rect 28264 10625 28282 10659
rect 28282 10625 28316 10659
rect 28264 10616 28316 10625
rect 29092 10616 29144 10668
rect 29736 10659 29788 10668
rect 29736 10625 29745 10659
rect 29745 10625 29779 10659
rect 29779 10625 29788 10659
rect 29736 10616 29788 10625
rect 31116 10616 31168 10668
rect 31668 10616 31720 10668
rect 33416 10659 33468 10668
rect 33416 10625 33450 10659
rect 33450 10625 33468 10659
rect 33416 10616 33468 10625
rect 31576 10548 31628 10600
rect 22468 10480 22520 10532
rect 2320 10455 2372 10464
rect 2320 10421 2329 10455
rect 2329 10421 2363 10455
rect 2363 10421 2372 10455
rect 2320 10412 2372 10421
rect 3240 10412 3292 10464
rect 18880 10412 18932 10464
rect 20720 10412 20772 10464
rect 22192 10412 22244 10464
rect 23204 10455 23256 10464
rect 23204 10421 23213 10455
rect 23213 10421 23247 10455
rect 23247 10421 23256 10455
rect 23204 10412 23256 10421
rect 23848 10412 23900 10464
rect 25228 10412 25280 10464
rect 26884 10412 26936 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 17960 10208 18012 10260
rect 19984 10208 20036 10260
rect 20720 10208 20772 10260
rect 21824 10251 21876 10260
rect 21824 10217 21833 10251
rect 21833 10217 21867 10251
rect 21867 10217 21876 10251
rect 21824 10208 21876 10217
rect 2320 10140 2372 10192
rect 23848 10183 23900 10192
rect 1584 10115 1636 10124
rect 1584 10081 1593 10115
rect 1593 10081 1627 10115
rect 1627 10081 1636 10115
rect 1584 10072 1636 10081
rect 3240 10115 3292 10124
rect 3240 10081 3249 10115
rect 3249 10081 3283 10115
rect 3283 10081 3292 10115
rect 3240 10072 3292 10081
rect 18420 10047 18472 10056
rect 18420 10013 18429 10047
rect 18429 10013 18463 10047
rect 18463 10013 18472 10047
rect 18420 10004 18472 10013
rect 18512 10004 18564 10056
rect 20536 10115 20588 10124
rect 20536 10081 20545 10115
rect 20545 10081 20579 10115
rect 20579 10081 20588 10115
rect 20536 10072 20588 10081
rect 23204 10072 23256 10124
rect 23848 10149 23857 10183
rect 23857 10149 23891 10183
rect 23891 10149 23900 10183
rect 23848 10140 23900 10149
rect 24860 10183 24912 10192
rect 24860 10149 24869 10183
rect 24869 10149 24903 10183
rect 24903 10149 24912 10183
rect 24860 10140 24912 10149
rect 25136 10072 25188 10124
rect 26700 10208 26752 10260
rect 26240 10072 26292 10124
rect 18880 10047 18932 10056
rect 18880 10013 18889 10047
rect 18889 10013 18923 10047
rect 18923 10013 18932 10047
rect 18880 10004 18932 10013
rect 20720 10004 20772 10056
rect 22744 10004 22796 10056
rect 24032 10004 24084 10056
rect 24676 10047 24728 10056
rect 24676 10013 24685 10047
rect 24685 10013 24719 10047
rect 24719 10013 24728 10047
rect 24676 10004 24728 10013
rect 25320 10004 25372 10056
rect 25596 10004 25648 10056
rect 26884 10047 26936 10056
rect 26884 10013 26893 10047
rect 26893 10013 26927 10047
rect 26927 10013 26936 10047
rect 26884 10004 26936 10013
rect 20812 9936 20864 9988
rect 21456 9979 21508 9988
rect 21456 9945 21465 9979
rect 21465 9945 21499 9979
rect 21499 9945 21508 9979
rect 21456 9936 21508 9945
rect 22284 9936 22336 9988
rect 23204 9936 23256 9988
rect 21272 9868 21324 9920
rect 23296 9868 23348 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 18420 9664 18472 9716
rect 20720 9596 20772 9648
rect 21272 9639 21324 9648
rect 21272 9605 21281 9639
rect 21281 9605 21315 9639
rect 21315 9605 21324 9639
rect 21272 9596 21324 9605
rect 22376 9664 22428 9716
rect 24032 9664 24084 9716
rect 25320 9664 25372 9716
rect 22192 9571 22244 9580
rect 22192 9537 22201 9571
rect 22201 9537 22235 9571
rect 22235 9537 22244 9571
rect 22192 9528 22244 9537
rect 22744 9528 22796 9580
rect 23204 9571 23256 9580
rect 23204 9537 23213 9571
rect 23213 9537 23247 9571
rect 23247 9537 23256 9571
rect 23204 9528 23256 9537
rect 23296 9528 23348 9580
rect 2044 9503 2096 9512
rect 2044 9469 2053 9503
rect 2053 9469 2087 9503
rect 2087 9469 2096 9503
rect 2044 9460 2096 9469
rect 2872 9460 2924 9512
rect 2964 9503 3016 9512
rect 2964 9469 2973 9503
rect 2973 9469 3007 9503
rect 3007 9469 3016 9503
rect 2964 9460 3016 9469
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 2044 9120 2096 9172
rect 2872 9163 2924 9172
rect 2872 9129 2881 9163
rect 2881 9129 2915 9163
rect 2915 9129 2924 9163
rect 2872 9120 2924 9129
rect 39580 9120 39632 9172
rect 2780 8916 2832 8968
rect 4988 8916 5040 8968
rect 48228 8891 48280 8900
rect 48228 8857 48237 8891
rect 48237 8857 48271 8891
rect 48271 8857 48280 8891
rect 48228 8848 48280 8857
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 48228 8440 48280 8492
rect 28540 8372 28592 8424
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 3424 7871 3476 7880
rect 3424 7837 3433 7871
rect 3433 7837 3467 7871
rect 3467 7837 3476 7871
rect 3424 7828 3476 7837
rect 1584 7803 1636 7812
rect 1584 7769 1593 7803
rect 1593 7769 1627 7803
rect 1627 7769 1636 7803
rect 1584 7760 1636 7769
rect 2872 7760 2924 7812
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 2872 7531 2924 7540
rect 2872 7497 2881 7531
rect 2881 7497 2915 7531
rect 2915 7497 2924 7531
rect 2872 7488 2924 7497
rect 3424 7420 3476 7472
rect 3148 7352 3200 7404
rect 5448 7352 5500 7404
rect 3424 7191 3476 7200
rect 3424 7157 3433 7191
rect 3433 7157 3467 7191
rect 3467 7157 3476 7191
rect 3424 7148 3476 7157
rect 43260 7191 43312 7200
rect 43260 7157 43269 7191
rect 43269 7157 43303 7191
rect 43303 7157 43312 7191
rect 43260 7148 43312 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 1584 6851 1636 6860
rect 1584 6817 1593 6851
rect 1593 6817 1627 6851
rect 1627 6817 1636 6851
rect 1584 6808 1636 6817
rect 3424 6851 3476 6860
rect 3424 6817 3433 6851
rect 3433 6817 3467 6851
rect 3467 6817 3476 6851
rect 3424 6808 3476 6817
rect 32220 6808 32272 6860
rect 43260 6808 43312 6860
rect 46848 6808 46900 6860
rect 46112 6740 46164 6792
rect 47308 6740 47360 6792
rect 47676 6783 47728 6792
rect 47676 6749 47685 6783
rect 47685 6749 47719 6783
rect 47719 6749 47728 6783
rect 47676 6740 47728 6749
rect 47952 6740 48004 6792
rect 2412 6672 2464 6724
rect 32404 6672 32456 6724
rect 43076 6672 43128 6724
rect 46296 6604 46348 6656
rect 47584 6647 47636 6656
rect 47584 6613 47593 6647
rect 47593 6613 47627 6647
rect 47627 6613 47636 6647
rect 47584 6604 47636 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 2412 6443 2464 6452
rect 2412 6409 2421 6443
rect 2421 6409 2455 6443
rect 2455 6409 2464 6443
rect 2412 6400 2464 6409
rect 32404 6443 32456 6452
rect 32404 6409 32413 6443
rect 32413 6409 32447 6443
rect 32447 6409 32456 6443
rect 32404 6400 32456 6409
rect 43076 6443 43128 6452
rect 43076 6409 43085 6443
rect 43085 6409 43119 6443
rect 43119 6409 43128 6443
rect 43076 6400 43128 6409
rect 2504 6307 2556 6316
rect 2504 6273 2513 6307
rect 2513 6273 2547 6307
rect 2547 6273 2556 6307
rect 2504 6264 2556 6273
rect 47308 6332 47360 6384
rect 43076 6264 43128 6316
rect 46388 6307 46440 6316
rect 46388 6273 46397 6307
rect 46397 6273 46431 6307
rect 46431 6273 46440 6307
rect 46388 6264 46440 6273
rect 47216 6307 47268 6316
rect 47216 6273 47225 6307
rect 47225 6273 47259 6307
rect 47259 6273 47268 6307
rect 47768 6307 47820 6316
rect 47216 6264 47268 6273
rect 47768 6273 47777 6307
rect 47777 6273 47811 6307
rect 47811 6273 47820 6307
rect 47768 6264 47820 6273
rect 47308 6196 47360 6248
rect 2964 6060 3016 6112
rect 3424 6060 3476 6112
rect 46940 6060 46992 6112
rect 47032 6060 47084 6112
rect 48136 6060 48188 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 2504 5788 2556 5840
rect 3424 5763 3476 5772
rect 3424 5729 3433 5763
rect 3433 5729 3467 5763
rect 3467 5729 3476 5763
rect 3424 5720 3476 5729
rect 46848 5788 46900 5840
rect 46112 5763 46164 5772
rect 46112 5729 46121 5763
rect 46121 5729 46155 5763
rect 46155 5729 46164 5763
rect 46112 5720 46164 5729
rect 46296 5763 46348 5772
rect 46296 5729 46305 5763
rect 46305 5729 46339 5763
rect 46339 5729 46348 5763
rect 46296 5720 46348 5729
rect 47124 5763 47176 5772
rect 47124 5729 47133 5763
rect 47133 5729 47167 5763
rect 47167 5729 47176 5763
rect 47124 5720 47176 5729
rect 17592 5652 17644 5704
rect 45652 5695 45704 5704
rect 45652 5661 45661 5695
rect 45661 5661 45695 5695
rect 45695 5661 45704 5695
rect 45652 5652 45704 5661
rect 1584 5627 1636 5636
rect 1584 5593 1593 5627
rect 1593 5593 1627 5627
rect 1627 5593 1636 5627
rect 1584 5584 1636 5593
rect 45560 5559 45612 5568
rect 45560 5525 45569 5559
rect 45569 5525 45603 5559
rect 45603 5525 45612 5559
rect 45560 5516 45612 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 47032 5287 47084 5296
rect 47032 5253 47041 5287
rect 47041 5253 47075 5287
rect 47075 5253 47084 5287
rect 47032 5244 47084 5253
rect 4620 5219 4672 5228
rect 4620 5185 4629 5219
rect 4629 5185 4663 5219
rect 4663 5185 4672 5219
rect 4620 5176 4672 5185
rect 12532 5176 12584 5228
rect 2780 5151 2832 5160
rect 2780 5117 2789 5151
rect 2789 5117 2823 5151
rect 2823 5117 2832 5151
rect 2780 5108 2832 5117
rect 3056 5108 3108 5160
rect 47216 5151 47268 5160
rect 2504 5040 2556 5092
rect 47216 5117 47225 5151
rect 47225 5117 47259 5151
rect 47259 5117 47268 5151
rect 47216 5108 47268 5117
rect 48412 5040 48464 5092
rect 4804 4972 4856 5024
rect 44732 5015 44784 5024
rect 44732 4981 44741 5015
rect 44741 4981 44775 5015
rect 44775 4981 44784 5015
rect 44732 4972 44784 4981
rect 48320 4972 48372 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 2504 4811 2556 4820
rect 2504 4777 2513 4811
rect 2513 4777 2547 4811
rect 2547 4777 2556 4811
rect 2504 4768 2556 4777
rect 3056 4811 3108 4820
rect 3056 4777 3065 4811
rect 3065 4777 3099 4811
rect 3099 4777 3108 4811
rect 3056 4768 3108 4777
rect 18236 4632 18288 4684
rect 1308 4564 1360 4616
rect 3240 4564 3292 4616
rect 4068 4564 4120 4616
rect 4712 4564 4764 4616
rect 5448 4607 5500 4616
rect 5448 4573 5457 4607
rect 5457 4573 5491 4607
rect 5491 4573 5500 4607
rect 5448 4564 5500 4573
rect 24860 4564 24912 4616
rect 39028 4607 39080 4616
rect 39028 4573 39037 4607
rect 39037 4573 39071 4607
rect 39071 4573 39080 4607
rect 39028 4564 39080 4573
rect 43076 4607 43128 4616
rect 43076 4573 43085 4607
rect 43085 4573 43119 4607
rect 43119 4573 43128 4607
rect 43076 4564 43128 4573
rect 44364 4564 44416 4616
rect 44548 4607 44600 4616
rect 44548 4573 44557 4607
rect 44557 4573 44591 4607
rect 44591 4573 44600 4607
rect 44548 4564 44600 4573
rect 47768 4700 47820 4752
rect 46848 4675 46900 4684
rect 46848 4641 46857 4675
rect 46857 4641 46891 4675
rect 46891 4641 46900 4675
rect 46848 4632 46900 4641
rect 48136 4675 48188 4684
rect 48136 4641 48145 4675
rect 48145 4641 48179 4675
rect 48179 4641 48188 4675
rect 48136 4632 48188 4641
rect 48320 4675 48372 4684
rect 48320 4641 48329 4675
rect 48329 4641 48363 4675
rect 48363 4641 48372 4675
rect 48320 4632 48372 4641
rect 46756 4564 46808 4616
rect 4988 4496 5040 4548
rect 19432 4496 19484 4548
rect 3516 4428 3568 4480
rect 5356 4471 5408 4480
rect 5356 4437 5365 4471
rect 5365 4437 5399 4471
rect 5399 4437 5408 4471
rect 5356 4428 5408 4437
rect 45100 4428 45152 4480
rect 45376 4428 45428 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 2780 4156 2832 4208
rect 4068 4131 4120 4140
rect 4068 4097 4077 4131
rect 4077 4097 4111 4131
rect 4111 4097 4120 4131
rect 5816 4131 5868 4140
rect 4068 4088 4120 4097
rect 5816 4097 5825 4131
rect 5825 4097 5859 4131
rect 5859 4097 5868 4131
rect 5816 4088 5868 4097
rect 7564 4131 7616 4140
rect 7564 4097 7573 4131
rect 7573 4097 7607 4131
rect 7607 4097 7616 4131
rect 7564 4088 7616 4097
rect 12532 4131 12584 4140
rect 12532 4097 12541 4131
rect 12541 4097 12575 4131
rect 12575 4097 12584 4131
rect 12532 4088 12584 4097
rect 13176 4131 13228 4140
rect 13176 4097 13185 4131
rect 13185 4097 13219 4131
rect 13219 4097 13228 4131
rect 13176 4088 13228 4097
rect 27160 4131 27212 4140
rect 7196 3952 7248 4004
rect 24860 4020 24912 4072
rect 27160 4097 27169 4131
rect 27169 4097 27203 4131
rect 27203 4097 27212 4131
rect 27160 4088 27212 4097
rect 38384 4131 38436 4140
rect 38384 4097 38393 4131
rect 38393 4097 38427 4131
rect 38427 4097 38436 4131
rect 38384 4088 38436 4097
rect 39028 4131 39080 4140
rect 39028 4097 39037 4131
rect 39037 4097 39071 4131
rect 39071 4097 39080 4131
rect 39028 4088 39080 4097
rect 41972 4088 42024 4140
rect 20168 3952 20220 4004
rect 38200 4020 38252 4072
rect 40500 4063 40552 4072
rect 40500 4029 40509 4063
rect 40509 4029 40543 4063
rect 40543 4029 40552 4063
rect 40500 4020 40552 4029
rect 44180 4020 44232 4072
rect 38108 3952 38160 4004
rect 38384 3952 38436 4004
rect 44088 3952 44140 4004
rect 3700 3884 3752 3936
rect 4620 3884 4672 3936
rect 4988 3927 5040 3936
rect 4988 3893 4997 3927
rect 4997 3893 5031 3927
rect 5031 3893 5040 3927
rect 4988 3884 5040 3893
rect 6092 3884 6144 3936
rect 6828 3884 6880 3936
rect 7656 3927 7708 3936
rect 7656 3893 7665 3927
rect 7665 3893 7699 3927
rect 7699 3893 7708 3927
rect 7656 3884 7708 3893
rect 10692 3884 10744 3936
rect 12532 3884 12584 3936
rect 13360 3884 13412 3936
rect 20076 3927 20128 3936
rect 20076 3893 20085 3927
rect 20085 3893 20119 3927
rect 20119 3893 20128 3927
rect 20076 3884 20128 3893
rect 24768 3884 24820 3936
rect 25964 3884 26016 3936
rect 27344 3884 27396 3936
rect 38936 3884 38988 3936
rect 40776 3884 40828 3936
rect 46756 4131 46808 4140
rect 46756 4097 46765 4131
rect 46765 4097 46799 4131
rect 46799 4097 46808 4131
rect 46756 4088 46808 4097
rect 47216 4088 47268 4140
rect 45744 4063 45796 4072
rect 45744 4029 45753 4063
rect 45753 4029 45787 4063
rect 45787 4029 45796 4063
rect 45744 4020 45796 4029
rect 47860 4020 47912 4072
rect 47584 3952 47636 4004
rect 47952 3884 48004 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 7196 3680 7248 3732
rect 12808 3680 12860 3732
rect 4804 3612 4856 3664
rect 4896 3612 4948 3664
rect 13176 3612 13228 3664
rect 17592 3612 17644 3664
rect 27160 3680 27212 3732
rect 43076 3680 43128 3732
rect 44088 3680 44140 3732
rect 47308 3680 47360 3732
rect 30288 3612 30340 3664
rect 38200 3655 38252 3664
rect 4712 3544 4764 3596
rect 6092 3587 6144 3596
rect 6092 3553 6101 3587
rect 6101 3553 6135 3587
rect 6135 3553 6144 3587
rect 6092 3544 6144 3553
rect 6460 3587 6512 3596
rect 6460 3553 6469 3587
rect 6469 3553 6503 3587
rect 6503 3553 6512 3587
rect 6460 3544 6512 3553
rect 10692 3587 10744 3596
rect 10692 3553 10701 3587
rect 10701 3553 10735 3587
rect 10735 3553 10744 3587
rect 10692 3544 10744 3553
rect 10968 3587 11020 3596
rect 10968 3553 10977 3587
rect 10977 3553 11011 3587
rect 11011 3553 11020 3587
rect 10968 3544 11020 3553
rect 25964 3587 26016 3596
rect 25964 3553 25973 3587
rect 25973 3553 26007 3587
rect 26007 3553 26016 3587
rect 25964 3544 26016 3553
rect 26424 3587 26476 3596
rect 26424 3553 26433 3587
rect 26433 3553 26467 3587
rect 26467 3553 26476 3587
rect 26424 3544 26476 3553
rect 1584 3519 1636 3528
rect 1584 3485 1593 3519
rect 1593 3485 1627 3519
rect 1627 3485 1636 3519
rect 1584 3476 1636 3485
rect 4160 3519 4212 3528
rect 4160 3485 4169 3519
rect 4169 3485 4203 3519
rect 4203 3485 4212 3519
rect 4160 3476 4212 3485
rect 4896 3476 4948 3528
rect 7472 3476 7524 3528
rect 10508 3519 10560 3528
rect 10508 3485 10517 3519
rect 10517 3485 10551 3519
rect 10551 3485 10560 3519
rect 10508 3476 10560 3485
rect 13176 3519 13228 3528
rect 13176 3485 13185 3519
rect 13185 3485 13219 3519
rect 13219 3485 13228 3519
rect 13176 3476 13228 3485
rect 16856 3476 16908 3528
rect 17592 3519 17644 3528
rect 17592 3485 17601 3519
rect 17601 3485 17635 3519
rect 17635 3485 17644 3519
rect 17592 3476 17644 3485
rect 19340 3476 19392 3528
rect 19432 3519 19484 3528
rect 19432 3485 19441 3519
rect 19441 3485 19475 3519
rect 19475 3485 19484 3519
rect 19432 3476 19484 3485
rect 19984 3476 20036 3528
rect 27160 3476 27212 3528
rect 33324 3408 33376 3460
rect 38200 3621 38209 3655
rect 38209 3621 38243 3655
rect 38243 3621 38252 3655
rect 38200 3612 38252 3621
rect 34060 3544 34112 3596
rect 45284 3612 45336 3664
rect 40776 3587 40828 3596
rect 40776 3553 40785 3587
rect 40785 3553 40819 3587
rect 40819 3553 40828 3587
rect 40776 3544 40828 3553
rect 41236 3587 41288 3596
rect 41236 3553 41245 3587
rect 41245 3553 41279 3587
rect 41279 3553 41288 3587
rect 41236 3544 41288 3553
rect 44548 3544 44600 3596
rect 45376 3587 45428 3596
rect 45376 3553 45385 3587
rect 45385 3553 45419 3587
rect 45419 3553 45428 3587
rect 45376 3544 45428 3553
rect 38108 3519 38160 3528
rect 38108 3485 38117 3519
rect 38117 3485 38151 3519
rect 38151 3485 38160 3519
rect 38108 3476 38160 3485
rect 38752 3519 38804 3528
rect 38752 3485 38761 3519
rect 38761 3485 38795 3519
rect 38795 3485 38804 3519
rect 38752 3476 38804 3485
rect 40592 3519 40644 3528
rect 40592 3485 40601 3519
rect 40601 3485 40635 3519
rect 40635 3485 40644 3519
rect 40592 3476 40644 3485
rect 41972 3476 42024 3528
rect 48320 3519 48372 3528
rect 4344 3340 4396 3392
rect 17040 3340 17092 3392
rect 19432 3340 19484 3392
rect 42800 3340 42852 3392
rect 43812 3408 43864 3460
rect 48320 3485 48329 3519
rect 48329 3485 48363 3519
rect 48363 3485 48372 3519
rect 48320 3476 48372 3485
rect 45652 3408 45704 3460
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 47860 3179 47912 3188
rect 47860 3145 47869 3179
rect 47869 3145 47903 3179
rect 47903 3145 47912 3179
rect 47860 3136 47912 3145
rect 3516 3111 3568 3120
rect 3516 3077 3525 3111
rect 3525 3077 3559 3111
rect 3559 3077 3568 3111
rect 3516 3068 3568 3077
rect 4344 3111 4396 3120
rect 4344 3077 4353 3111
rect 4353 3077 4387 3111
rect 4387 3077 4396 3111
rect 4344 3068 4396 3077
rect 7656 3111 7708 3120
rect 7656 3077 7665 3111
rect 7665 3077 7699 3111
rect 7699 3077 7708 3111
rect 7656 3068 7708 3077
rect 13360 3111 13412 3120
rect 13360 3077 13369 3111
rect 13369 3077 13403 3111
rect 13403 3077 13412 3111
rect 13360 3068 13412 3077
rect 17040 3111 17092 3120
rect 17040 3077 17049 3111
rect 17049 3077 17083 3111
rect 17083 3077 17092 3111
rect 17040 3068 17092 3077
rect 19432 3068 19484 3120
rect 27344 3111 27396 3120
rect 27344 3077 27353 3111
rect 27353 3077 27387 3111
rect 27387 3077 27396 3111
rect 27344 3068 27396 3077
rect 38936 3111 38988 3120
rect 38936 3077 38945 3111
rect 38945 3077 38979 3111
rect 38979 3077 38988 3111
rect 38936 3068 38988 3077
rect 42800 3111 42852 3120
rect 42800 3077 42809 3111
rect 42809 3077 42843 3111
rect 42843 3077 42852 3111
rect 42800 3068 42852 3077
rect 45100 3111 45152 3120
rect 45100 3077 45109 3111
rect 45109 3077 45143 3111
rect 45143 3077 45152 3111
rect 45100 3068 45152 3077
rect 3700 3043 3752 3052
rect 3700 3009 3709 3043
rect 3709 3009 3743 3043
rect 3743 3009 3752 3043
rect 7472 3043 7524 3052
rect 3700 3000 3752 3009
rect 7472 3009 7481 3043
rect 7481 3009 7515 3043
rect 7515 3009 7524 3043
rect 7472 3000 7524 3009
rect 10508 3043 10560 3052
rect 10508 3009 10517 3043
rect 10517 3009 10551 3043
rect 10551 3009 10560 3043
rect 10508 3000 10560 3009
rect 11612 3000 11664 3052
rect 13176 3043 13228 3052
rect 13176 3009 13185 3043
rect 13185 3009 13219 3043
rect 13219 3009 13228 3043
rect 13176 3000 13228 3009
rect 16856 3043 16908 3052
rect 16856 3009 16865 3043
rect 16865 3009 16899 3043
rect 16899 3009 16908 3043
rect 16856 3000 16908 3009
rect 24768 3043 24820 3052
rect 24768 3009 24777 3043
rect 24777 3009 24811 3043
rect 24811 3009 24820 3043
rect 24768 3000 24820 3009
rect 27160 3043 27212 3052
rect 27160 3009 27169 3043
rect 27169 3009 27203 3043
rect 27203 3009 27212 3043
rect 27160 3000 27212 3009
rect 38752 3043 38804 3052
rect 38752 3009 38761 3043
rect 38761 3009 38795 3043
rect 38795 3009 38804 3043
rect 38752 3000 38804 3009
rect 40592 3000 40644 3052
rect 44364 3000 44416 3052
rect 46296 3000 46348 3052
rect 3240 2975 3292 2984
rect 3240 2941 3249 2975
rect 3249 2941 3283 2975
rect 3283 2941 3292 2975
rect 3240 2932 3292 2941
rect 4988 2932 5040 2984
rect 5172 2975 5224 2984
rect 5172 2941 5181 2975
rect 5181 2941 5215 2975
rect 5215 2941 5224 2975
rect 5172 2932 5224 2941
rect 7748 2932 7800 2984
rect 13544 2932 13596 2984
rect 17408 2975 17460 2984
rect 17408 2941 17417 2975
rect 17417 2941 17451 2975
rect 17451 2941 17460 2975
rect 17408 2932 17460 2941
rect 20076 2932 20128 2984
rect 20628 2975 20680 2984
rect 20628 2941 20637 2975
rect 20637 2941 20671 2975
rect 20671 2941 20680 2975
rect 20628 2932 20680 2941
rect 24952 2975 25004 2984
rect 24952 2941 24961 2975
rect 24961 2941 24995 2975
rect 24995 2941 25004 2975
rect 24952 2932 25004 2941
rect 25780 2975 25832 2984
rect 25780 2941 25789 2975
rect 25789 2941 25823 2975
rect 25823 2941 25832 2975
rect 25780 2932 25832 2941
rect 27712 2975 27764 2984
rect 27712 2941 27721 2975
rect 27721 2941 27755 2975
rect 27755 2941 27764 2975
rect 27712 2932 27764 2941
rect 39304 2975 39356 2984
rect 39304 2941 39313 2975
rect 39313 2941 39347 2975
rect 39347 2941 39356 2975
rect 39304 2932 39356 2941
rect 46756 2975 46808 2984
rect 23572 2864 23624 2916
rect 6644 2839 6696 2848
rect 6644 2805 6653 2839
rect 6653 2805 6687 2839
rect 6687 2805 6696 2839
rect 6644 2796 6696 2805
rect 12440 2839 12492 2848
rect 12440 2805 12449 2839
rect 12449 2805 12483 2839
rect 12483 2805 12492 2839
rect 12440 2796 12492 2805
rect 41880 2796 41932 2848
rect 46756 2941 46765 2975
rect 46765 2941 46799 2975
rect 46799 2941 46808 2975
rect 46756 2932 46808 2941
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 12624 2592 12676 2644
rect 24952 2592 25004 2644
rect 29644 2592 29696 2644
rect 1584 2499 1636 2508
rect 1584 2465 1593 2499
rect 1593 2465 1627 2499
rect 1627 2465 1636 2499
rect 1584 2456 1636 2465
rect 2964 2456 3016 2508
rect 4068 2499 4120 2508
rect 4068 2465 4077 2499
rect 4077 2465 4111 2499
rect 4111 2465 4120 2499
rect 4068 2456 4120 2465
rect 4528 2499 4580 2508
rect 4528 2465 4537 2499
rect 4537 2465 4571 2499
rect 4571 2465 4580 2499
rect 4528 2456 4580 2465
rect 6644 2499 6696 2508
rect 6644 2465 6653 2499
rect 6653 2465 6687 2499
rect 6687 2465 6696 2499
rect 6644 2456 6696 2465
rect 6828 2499 6880 2508
rect 6828 2465 6837 2499
rect 6837 2465 6871 2499
rect 6871 2465 6880 2499
rect 6828 2456 6880 2465
rect 7104 2499 7156 2508
rect 7104 2465 7113 2499
rect 7113 2465 7147 2499
rect 7147 2465 7156 2499
rect 7104 2456 7156 2465
rect 12440 2456 12492 2508
rect 12900 2499 12952 2508
rect 12900 2465 12909 2499
rect 12909 2465 12943 2499
rect 12943 2465 12952 2499
rect 12900 2456 12952 2465
rect 19340 2456 19392 2508
rect 19616 2456 19668 2508
rect 48964 2524 49016 2576
rect 44732 2456 44784 2508
rect 47676 2456 47728 2508
rect 14188 2388 14240 2440
rect 38384 2388 38436 2440
rect 4620 2320 4672 2372
rect 12532 2320 12584 2372
rect 20168 2320 20220 2372
rect 29000 2320 29052 2372
rect 38660 2320 38712 2372
rect 45560 2320 45612 2372
rect 46940 2320 46992 2372
rect 5356 2252 5408 2304
rect 30656 2252 30708 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 44180 2048 44232 2100
rect 46848 2048 46900 2100
rect 2872 1640 2924 1692
rect 5540 1640 5592 1692
<< metal2 >>
rect 47044 49830 47256 49858
rect 47044 49800 47072 49830
rect -10 49200 102 49800
rect 1278 49200 1390 49800
rect 1922 49200 2034 49800
rect 2566 49200 2678 49800
rect 3854 49200 3966 49800
rect 4498 49200 4610 49800
rect 5786 49200 5898 49800
rect 6430 49200 6542 49800
rect 7718 49200 7830 49800
rect 8362 49200 8474 49800
rect 9006 49200 9118 49800
rect 10294 49200 10406 49800
rect 10938 49200 11050 49800
rect 12226 49200 12338 49800
rect 12870 49200 12982 49800
rect 14158 49200 14270 49800
rect 14802 49200 14914 49800
rect 15446 49200 15558 49800
rect 16734 49200 16846 49800
rect 17378 49200 17490 49800
rect 18666 49200 18778 49800
rect 19310 49200 19422 49800
rect 20598 49200 20710 49800
rect 21242 49200 21354 49800
rect 21886 49200 21998 49800
rect 23174 49200 23286 49800
rect 23818 49200 23930 49800
rect 25106 49200 25218 49800
rect 25750 49200 25862 49800
rect 27038 49200 27150 49800
rect 27682 49200 27794 49800
rect 28970 49200 29082 49800
rect 29614 49200 29726 49800
rect 30258 49200 30370 49800
rect 31546 49200 31658 49800
rect 32190 49200 32302 49800
rect 33478 49200 33590 49800
rect 34122 49200 34234 49800
rect 35410 49200 35522 49800
rect 36054 49200 36166 49800
rect 36698 49200 36810 49800
rect 37986 49200 38098 49800
rect 38630 49200 38742 49800
rect 39918 49200 40030 49800
rect 40562 49200 40674 49800
rect 41850 49200 41962 49800
rect 42494 49200 42606 49800
rect 43138 49200 43250 49800
rect 44426 49200 44538 49800
rect 45070 49200 45182 49800
rect 46358 49200 46470 49800
rect 47002 49200 47114 49800
rect 47228 49314 47256 49830
rect 47228 49286 47348 49314
rect 1320 46918 1348 49200
rect 1308 46912 1360 46918
rect 1308 46854 1360 46860
rect 1964 46714 1992 49200
rect 2320 46980 2372 46986
rect 2320 46922 2372 46928
rect 1952 46708 2004 46714
rect 1952 46650 2004 46656
rect 2332 44878 2360 46922
rect 2608 46510 2636 49200
rect 2870 48376 2926 48385
rect 2870 48311 2926 48320
rect 2778 47696 2834 47705
rect 2778 47631 2834 47640
rect 2596 46504 2648 46510
rect 2596 46446 2648 46452
rect 2792 46034 2820 47631
rect 2780 46028 2832 46034
rect 2780 45970 2832 45976
rect 2884 45422 2912 48311
rect 4540 47546 4568 49200
rect 4540 47518 4660 47546
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4528 47048 4580 47054
rect 4528 46990 4580 46996
rect 3516 46912 3568 46918
rect 3516 46854 3568 46860
rect 3528 46646 3556 46854
rect 3516 46640 3568 46646
rect 3516 46582 3568 46588
rect 4540 46578 4568 46990
rect 4632 46646 4660 47518
rect 4804 47184 4856 47190
rect 4804 47126 4856 47132
rect 4712 46980 4764 46986
rect 4712 46922 4764 46928
rect 4620 46640 4672 46646
rect 4620 46582 4672 46588
rect 4528 46572 4580 46578
rect 4528 46514 4580 46520
rect 4068 46436 4120 46442
rect 4068 46378 4120 46384
rect 4080 46345 4108 46378
rect 4066 46336 4122 46345
rect 4066 46271 4122 46280
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4620 46028 4672 46034
rect 4620 45970 4672 45976
rect 3146 45656 3202 45665
rect 3146 45591 3202 45600
rect 2872 45416 2924 45422
rect 2872 45358 2924 45364
rect 2044 44872 2096 44878
rect 2044 44814 2096 44820
rect 2320 44872 2372 44878
rect 2320 44814 2372 44820
rect 2056 44402 2084 44814
rect 2044 44396 2096 44402
rect 2044 44338 2096 44344
rect 3160 44334 3188 45591
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 3240 44804 3292 44810
rect 3240 44746 3292 44752
rect 3252 44470 3280 44746
rect 4632 44538 4660 45970
rect 4620 44532 4672 44538
rect 4620 44474 4672 44480
rect 3240 44464 3292 44470
rect 3240 44406 3292 44412
rect 3056 44328 3108 44334
rect 3056 44270 3108 44276
rect 3148 44328 3200 44334
rect 3148 44270 3200 44276
rect 2044 43784 2096 43790
rect 2044 43726 2096 43732
rect 2056 43314 2084 43726
rect 2778 43616 2834 43625
rect 2778 43551 2834 43560
rect 2044 43308 2096 43314
rect 2044 43250 2096 43256
rect 2792 43246 2820 43551
rect 2228 43240 2280 43246
rect 2228 43182 2280 43188
rect 2780 43240 2832 43246
rect 2780 43182 2832 43188
rect 2240 42906 2268 43182
rect 2228 42900 2280 42906
rect 2228 42842 2280 42848
rect 3068 42770 3096 44270
rect 3056 42764 3108 42770
rect 3056 42706 3108 42712
rect 2504 42696 2556 42702
rect 2504 42638 2556 42644
rect 1676 38956 1728 38962
rect 1676 38898 1728 38904
rect 1688 38865 1716 38898
rect 1674 38856 1730 38865
rect 1674 38791 1730 38800
rect 1860 38820 1912 38826
rect 1860 38762 1912 38768
rect 1676 37188 1728 37194
rect 1676 37130 1728 37136
rect 1688 36825 1716 37130
rect 1674 36816 1730 36825
rect 1674 36751 1730 36760
rect 1584 34604 1636 34610
rect 1584 34546 1636 34552
rect 1596 34105 1624 34546
rect 1582 34096 1638 34105
rect 1582 34031 1638 34040
rect 1584 32428 1636 32434
rect 1584 32370 1636 32376
rect 1596 32065 1624 32370
rect 1582 32056 1638 32065
rect 1582 31991 1638 32000
rect 204 29776 256 29782
rect 204 29718 256 29724
rect 216 16574 244 29718
rect 1872 27334 1900 38762
rect 1952 34740 2004 34746
rect 1952 34682 2004 34688
rect 1860 27328 1912 27334
rect 1860 27270 1912 27276
rect 1584 25288 1636 25294
rect 1582 25256 1584 25265
rect 1636 25256 1638 25265
rect 1582 25191 1638 25200
rect 1584 21956 1636 21962
rect 1584 21898 1636 21904
rect 1596 21865 1624 21898
rect 1582 21856 1638 21865
rect 1582 21791 1638 21800
rect 1964 17338 1992 34682
rect 2044 20936 2096 20942
rect 2044 20878 2096 20884
rect 2056 20466 2084 20878
rect 2044 20460 2096 20466
rect 2044 20402 2096 20408
rect 2412 20392 2464 20398
rect 2412 20334 2464 20340
rect 2424 20058 2452 20334
rect 2412 20052 2464 20058
rect 2412 19994 2464 20000
rect 2516 19854 2544 42638
rect 3054 41576 3110 41585
rect 3054 41511 3056 41520
rect 3108 41511 3110 41520
rect 3056 41482 3108 41488
rect 3252 41414 3280 44406
rect 4620 44260 4672 44266
rect 4620 44202 4672 44208
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 3516 43852 3568 43858
rect 3516 43794 3568 43800
rect 3528 43314 3556 43794
rect 3516 43308 3568 43314
rect 3516 43250 3568 43256
rect 3528 42838 3556 43250
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 3516 42832 3568 42838
rect 3516 42774 3568 42780
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 3068 41386 3280 41414
rect 2688 37324 2740 37330
rect 2688 37266 2740 37272
rect 2700 33114 2728 37266
rect 2688 33108 2740 33114
rect 2688 33050 2740 33056
rect 3068 26234 3096 41386
rect 3238 40896 3294 40905
rect 3238 40831 3294 40840
rect 3252 40118 3280 40831
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 3240 40112 3292 40118
rect 3240 40054 3292 40060
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4068 36712 4120 36718
rect 4068 36654 4120 36660
rect 4080 36378 4108 36654
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4068 36372 4120 36378
rect 4068 36314 4120 36320
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4344 35080 4396 35086
rect 4344 35022 4396 35028
rect 4356 34746 4384 35022
rect 4344 34740 4396 34746
rect 4344 34682 4396 34688
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4160 33992 4212 33998
rect 4160 33934 4212 33940
rect 4172 33658 4200 33934
rect 4160 33652 4212 33658
rect 4160 33594 4212 33600
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 3792 32904 3844 32910
rect 3792 32846 3844 32852
rect 3804 32434 3832 32846
rect 4066 32736 4122 32745
rect 4066 32671 4122 32680
rect 3792 32428 3844 32434
rect 3792 32370 3844 32376
rect 4080 32366 4108 32671
rect 3976 32360 4028 32366
rect 3976 32302 4028 32308
rect 4068 32360 4120 32366
rect 4068 32302 4120 32308
rect 3988 32026 4016 32302
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 3976 32020 4028 32026
rect 3976 31962 4028 31968
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 2976 26206 3096 26234
rect 2596 24812 2648 24818
rect 2596 24754 2648 24760
rect 2608 22642 2636 24754
rect 2596 22636 2648 22642
rect 2596 22578 2648 22584
rect 2778 20496 2834 20505
rect 2778 20431 2834 20440
rect 2792 20398 2820 20431
rect 2780 20392 2832 20398
rect 2780 20334 2832 20340
rect 2504 19848 2556 19854
rect 2504 19790 2556 19796
rect 2044 18760 2096 18766
rect 2044 18702 2096 18708
rect 2056 18290 2084 18702
rect 2778 18456 2834 18465
rect 2778 18391 2834 18400
rect 2044 18284 2096 18290
rect 2044 18226 2096 18232
rect 2792 18222 2820 18391
rect 2228 18216 2280 18222
rect 2228 18158 2280 18164
rect 2780 18216 2832 18222
rect 2780 18158 2832 18164
rect 2240 17882 2268 18158
rect 2228 17876 2280 17882
rect 2228 17818 2280 17824
rect 2596 17672 2648 17678
rect 2596 17614 2648 17620
rect 1952 17332 2004 17338
rect 1952 17274 2004 17280
rect 2044 17128 2096 17134
rect 2044 17070 2096 17076
rect 2056 16794 2084 17070
rect 2044 16788 2096 16794
rect 2044 16730 2096 16736
rect 216 16546 704 16574
rect 676 800 704 16546
rect 1584 14408 1636 14414
rect 1582 14376 1584 14385
rect 1636 14376 1638 14385
rect 1582 14311 1638 14320
rect 2412 14340 2464 14346
rect 2412 14282 2464 14288
rect 2424 14074 2452 14282
rect 2412 14068 2464 14074
rect 2412 14010 2464 14016
rect 2504 13932 2556 13938
rect 2504 13874 2556 13880
rect 2228 12096 2280 12102
rect 2228 12038 2280 12044
rect 2240 11830 2268 12038
rect 2228 11824 2280 11830
rect 2228 11766 2280 11772
rect 2044 11688 2096 11694
rect 2044 11630 2096 11636
rect 2056 11354 2084 11630
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 2320 10464 2372 10470
rect 2320 10406 2372 10412
rect 1582 10296 1638 10305
rect 1582 10231 1638 10240
rect 1596 10130 1624 10231
rect 2332 10198 2360 10406
rect 2320 10192 2372 10198
rect 2320 10134 2372 10140
rect 1584 10124 1636 10130
rect 1584 10066 1636 10072
rect 2044 9512 2096 9518
rect 2044 9454 2096 9460
rect 2056 9178 2084 9454
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 1584 7812 1636 7818
rect 1584 7754 1636 7760
rect 1596 7585 1624 7754
rect 1582 7576 1638 7585
rect 1582 7511 1638 7520
rect 1582 6896 1638 6905
rect 1582 6831 1584 6840
rect 1636 6831 1638 6840
rect 1584 6802 1636 6808
rect 2412 6724 2464 6730
rect 2412 6666 2464 6672
rect 2424 6458 2452 6666
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 2516 6322 2544 13874
rect 2608 12238 2636 17614
rect 2780 17128 2832 17134
rect 2872 17128 2924 17134
rect 2780 17070 2832 17076
rect 2870 17096 2872 17105
rect 2924 17096 2926 17105
rect 2792 16590 2820 17070
rect 2870 17031 2926 17040
rect 2976 16590 3004 26206
rect 3424 25696 3476 25702
rect 3424 25638 3476 25644
rect 3436 25362 3464 25638
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 3424 25356 3476 25362
rect 3424 25298 3476 25304
rect 3240 25220 3292 25226
rect 3240 25162 3292 25168
rect 3252 24750 3280 25162
rect 3240 24744 3292 24750
rect 3240 24686 3292 24692
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 3332 24132 3384 24138
rect 3332 24074 3384 24080
rect 3344 23905 3372 24074
rect 3330 23896 3386 23905
rect 3330 23831 3386 23840
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 3240 22432 3292 22438
rect 3240 22374 3292 22380
rect 3252 22098 3280 22374
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 3240 22092 3292 22098
rect 3240 22034 3292 22040
rect 3424 22024 3476 22030
rect 3424 21966 3476 21972
rect 3436 21554 3464 21966
rect 3424 21548 3476 21554
rect 3424 21490 3476 21496
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 3148 19848 3200 19854
rect 3148 19790 3200 19796
rect 2780 16584 2832 16590
rect 2780 16526 2832 16532
rect 2964 16584 3016 16590
rect 2964 16526 3016 16532
rect 2976 12434 3004 16526
rect 2976 12406 3096 12434
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2608 11098 2636 12174
rect 2780 11688 2832 11694
rect 2778 11656 2780 11665
rect 2832 11656 2834 11665
rect 2778 11591 2834 11600
rect 2608 11070 2820 11098
rect 2792 8974 2820 11070
rect 2962 9616 3018 9625
rect 2962 9551 3018 9560
rect 2976 9518 3004 9551
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 2884 9178 2912 9454
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 2872 7812 2924 7818
rect 2872 7754 2924 7760
rect 2884 7546 2912 7754
rect 2872 7540 2924 7546
rect 2872 7482 2924 7488
rect 3068 6914 3096 12406
rect 3160 7410 3188 19790
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 3424 15088 3476 15094
rect 3422 15056 3424 15065
rect 3476 15056 3478 15065
rect 3422 14991 3478 15000
rect 3424 14816 3476 14822
rect 3424 14758 3476 14764
rect 3436 14482 3464 14758
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 3424 14476 3476 14482
rect 3424 14418 3476 14424
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4632 10674 4660 44202
rect 4724 12782 4752 46922
rect 4816 45966 4844 47126
rect 4988 47116 5040 47122
rect 4988 47058 5040 47064
rect 4896 46368 4948 46374
rect 4896 46310 4948 46316
rect 4804 45960 4856 45966
rect 4804 45902 4856 45908
rect 4908 45422 4936 46310
rect 4896 45416 4948 45422
rect 4896 45358 4948 45364
rect 5000 45082 5028 47058
rect 5828 46594 5856 49200
rect 7196 47252 7248 47258
rect 7196 47194 7248 47200
rect 6000 47116 6052 47122
rect 6000 47058 6052 47064
rect 5736 46566 5856 46594
rect 6012 46578 6040 47058
rect 7208 46714 7236 47194
rect 8300 47184 8352 47190
rect 8300 47126 8352 47132
rect 7196 46708 7248 46714
rect 7196 46650 7248 46656
rect 6000 46572 6052 46578
rect 5080 46096 5132 46102
rect 5080 46038 5132 46044
rect 4988 45076 5040 45082
rect 4988 45018 5040 45024
rect 4988 44396 5040 44402
rect 4988 44338 5040 44344
rect 5000 43790 5028 44338
rect 5092 44266 5120 46038
rect 5540 45892 5592 45898
rect 5540 45834 5592 45840
rect 5552 45490 5580 45834
rect 5540 45484 5592 45490
rect 5540 45426 5592 45432
rect 5356 45416 5408 45422
rect 5356 45358 5408 45364
rect 5172 44396 5224 44402
rect 5172 44338 5224 44344
rect 5080 44260 5132 44266
rect 5080 44202 5132 44208
rect 4988 43784 5040 43790
rect 4988 43726 5040 43732
rect 5000 42702 5028 43726
rect 5184 43382 5212 44338
rect 5264 43852 5316 43858
rect 5264 43794 5316 43800
rect 5172 43376 5224 43382
rect 5172 43318 5224 43324
rect 4988 42696 5040 42702
rect 4988 42638 5040 42644
rect 5184 41414 5212 43318
rect 5276 42770 5304 43794
rect 5264 42764 5316 42770
rect 5264 42706 5316 42712
rect 5092 41386 5212 41414
rect 4804 38344 4856 38350
rect 4804 38286 4856 38292
rect 4816 37874 4844 38286
rect 4804 37868 4856 37874
rect 4804 37810 4856 37816
rect 4816 37754 4844 37810
rect 4816 37726 5028 37754
rect 4804 37664 4856 37670
rect 4804 37606 4856 37612
rect 4816 37330 4844 37606
rect 4804 37324 4856 37330
rect 4804 37266 4856 37272
rect 4896 37256 4948 37262
rect 4896 37198 4948 37204
rect 4908 36378 4936 37198
rect 4896 36372 4948 36378
rect 4896 36314 4948 36320
rect 4896 36236 4948 36242
rect 4896 36178 4948 36184
rect 4804 34604 4856 34610
rect 4804 34546 4856 34552
rect 4816 33522 4844 34546
rect 4804 33516 4856 33522
rect 4804 33458 4856 33464
rect 4908 26234 4936 36178
rect 5000 36174 5028 37726
rect 4988 36168 5040 36174
rect 4988 36110 5040 36116
rect 5000 34610 5028 36110
rect 4988 34604 5040 34610
rect 4988 34546 5040 34552
rect 4988 34468 5040 34474
rect 4988 34410 5040 34416
rect 5000 33522 5028 34410
rect 4988 33516 5040 33522
rect 4988 33458 5040 33464
rect 5000 33046 5028 33458
rect 4988 33040 5040 33046
rect 4988 32982 5040 32988
rect 4816 26206 4936 26234
rect 5092 26234 5120 41386
rect 5172 35692 5224 35698
rect 5172 35634 5224 35640
rect 5184 34542 5212 35634
rect 5172 34536 5224 34542
rect 5172 34478 5224 34484
rect 5172 34400 5224 34406
rect 5172 34342 5224 34348
rect 5184 34066 5212 34342
rect 5172 34060 5224 34066
rect 5172 34002 5224 34008
rect 5276 33946 5304 42706
rect 5368 36242 5396 45358
rect 5448 45280 5500 45286
rect 5448 45222 5500 45228
rect 5460 45082 5488 45222
rect 5448 45076 5500 45082
rect 5448 45018 5500 45024
rect 5460 36666 5488 45018
rect 5552 44878 5580 45426
rect 5540 44872 5592 44878
rect 5540 44814 5592 44820
rect 5552 44470 5580 44814
rect 5540 44464 5592 44470
rect 5540 44406 5592 44412
rect 5736 43858 5764 46566
rect 6000 46514 6052 46520
rect 5816 46504 5868 46510
rect 5816 46446 5868 46452
rect 5828 46170 5856 46446
rect 5816 46164 5868 46170
rect 5816 46106 5868 46112
rect 6368 45960 6420 45966
rect 6368 45902 6420 45908
rect 7012 45960 7064 45966
rect 7012 45902 7064 45908
rect 6380 45422 6408 45902
rect 6920 45824 6972 45830
rect 6920 45766 6972 45772
rect 6932 45558 6960 45766
rect 7024 45558 7052 45902
rect 6920 45552 6972 45558
rect 6920 45494 6972 45500
rect 7012 45552 7064 45558
rect 7012 45494 7064 45500
rect 6736 45484 6788 45490
rect 6736 45426 6788 45432
rect 6368 45416 6420 45422
rect 6368 45358 6420 45364
rect 6748 45286 6776 45426
rect 7380 45416 7432 45422
rect 7380 45358 7432 45364
rect 6736 45280 6788 45286
rect 6736 45222 6788 45228
rect 5816 44328 5868 44334
rect 5816 44270 5868 44276
rect 5724 43852 5776 43858
rect 5724 43794 5776 43800
rect 5632 42628 5684 42634
rect 5632 42570 5684 42576
rect 5460 36638 5580 36666
rect 5448 36576 5500 36582
rect 5448 36518 5500 36524
rect 5460 36378 5488 36518
rect 5448 36372 5500 36378
rect 5448 36314 5500 36320
rect 5552 36258 5580 36638
rect 5356 36236 5408 36242
rect 5356 36178 5408 36184
rect 5460 36230 5580 36258
rect 5460 35894 5488 36230
rect 5184 33918 5304 33946
rect 5368 35866 5488 35894
rect 5184 29850 5212 33918
rect 5264 33856 5316 33862
rect 5264 33798 5316 33804
rect 5276 33318 5304 33798
rect 5264 33312 5316 33318
rect 5264 33254 5316 33260
rect 5172 29844 5224 29850
rect 5172 29786 5224 29792
rect 5368 26234 5396 35866
rect 5448 35488 5500 35494
rect 5448 35430 5500 35436
rect 5460 35290 5488 35430
rect 5448 35284 5500 35290
rect 5448 35226 5500 35232
rect 5448 32836 5500 32842
rect 5448 32778 5500 32784
rect 5460 32570 5488 32778
rect 5448 32564 5500 32570
rect 5448 32506 5500 32512
rect 5460 31822 5488 32506
rect 5448 31816 5500 31822
rect 5448 31758 5500 31764
rect 5644 29170 5672 42570
rect 5828 41414 5856 44270
rect 5908 43716 5960 43722
rect 5908 43658 5960 43664
rect 5920 43450 5948 43658
rect 5908 43444 5960 43450
rect 5908 43386 5960 43392
rect 6748 43382 6776 45222
rect 7392 45014 7420 45358
rect 7380 45008 7432 45014
rect 7380 44950 7432 44956
rect 6828 44940 6880 44946
rect 6828 44882 6880 44888
rect 6840 44538 6868 44882
rect 6828 44532 6880 44538
rect 6828 44474 6880 44480
rect 6736 43376 6788 43382
rect 6736 43318 6788 43324
rect 6000 43308 6052 43314
rect 6000 43250 6052 43256
rect 6012 42634 6040 43250
rect 6000 42628 6052 42634
rect 6000 42570 6052 42576
rect 6840 41414 6868 44474
rect 7288 44192 7340 44198
rect 7288 44134 7340 44140
rect 7300 43858 7328 44134
rect 7288 43852 7340 43858
rect 7288 43794 7340 43800
rect 7288 42016 7340 42022
rect 7288 41958 7340 41964
rect 7300 41682 7328 41958
rect 7288 41676 7340 41682
rect 7288 41618 7340 41624
rect 7104 41540 7156 41546
rect 7104 41482 7156 41488
rect 5736 41386 5856 41414
rect 6748 41386 6868 41414
rect 5736 35894 5764 41386
rect 6092 41132 6144 41138
rect 6092 41074 6144 41080
rect 5816 37868 5868 37874
rect 5816 37810 5868 37816
rect 5828 37398 5856 37810
rect 5816 37392 5868 37398
rect 5816 37334 5868 37340
rect 6000 36780 6052 36786
rect 6000 36722 6052 36728
rect 6012 36378 6040 36722
rect 6000 36372 6052 36378
rect 6000 36314 6052 36320
rect 5736 35866 5856 35894
rect 5724 35012 5776 35018
rect 5724 34954 5776 34960
rect 5736 34746 5764 34954
rect 5724 34740 5776 34746
rect 5724 34682 5776 34688
rect 5632 29164 5684 29170
rect 5632 29106 5684 29112
rect 5540 28620 5592 28626
rect 5540 28562 5592 28568
rect 5092 26206 5212 26234
rect 4816 22094 4844 26206
rect 4816 22066 4936 22094
rect 4712 12776 4764 12782
rect 4712 12718 4764 12724
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 3240 10464 3292 10470
rect 3240 10406 3292 10412
rect 3252 10130 3280 10406
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 3240 10124 3292 10130
rect 3240 10066 3292 10072
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3424 7880 3476 7886
rect 3424 7822 3476 7828
rect 3436 7478 3464 7822
rect 3424 7472 3476 7478
rect 3424 7414 3476 7420
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3424 7200 3476 7206
rect 3424 7142 3476 7148
rect 3068 6886 3280 6914
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 2516 5846 2544 6258
rect 2964 6112 3016 6118
rect 2964 6054 3016 6060
rect 2504 5840 2556 5846
rect 2504 5782 2556 5788
rect 1584 5636 1636 5642
rect 1584 5578 1636 5584
rect 1596 5545 1624 5578
rect 1582 5536 1638 5545
rect 1582 5471 1638 5480
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 2504 5092 2556 5098
rect 2504 5034 2556 5040
rect 2516 4826 2544 5034
rect 2792 4865 2820 5102
rect 2778 4856 2834 4865
rect 2504 4820 2556 4826
rect 2778 4791 2834 4800
rect 2504 4762 2556 4768
rect 1308 4616 1360 4622
rect 1308 4558 1360 4564
rect 1320 800 1348 4558
rect 2780 4208 2832 4214
rect 2780 4150 2832 4156
rect 1584 3528 1636 3534
rect 1582 3496 1584 3505
rect 1636 3496 1638 3505
rect 1582 3431 1638 3440
rect 1582 2816 1638 2825
rect 1582 2751 1638 2760
rect 1596 2514 1624 2751
rect 1584 2508 1636 2514
rect 1584 2450 1636 2456
rect -10 200 102 800
rect 634 200 746 800
rect 1278 200 1390 800
rect 2566 200 2678 800
rect 2792 785 2820 4150
rect 2976 2514 3004 6054
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 3068 4826 3096 5102
rect 3056 4820 3108 4826
rect 3056 4762 3108 4768
rect 3252 4622 3280 6886
rect 3436 6866 3464 7142
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3436 5778 3464 6054
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 3424 5772 3476 5778
rect 3424 5714 3476 5720
rect 4632 5234 4660 10610
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 3516 4480 3568 4486
rect 3516 4422 3568 4428
rect 3528 3126 3556 4422
rect 4080 4146 4108 4558
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 3700 3936 3752 3942
rect 3700 3878 3752 3884
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 3516 3120 3568 3126
rect 3516 3062 3568 3068
rect 3712 3058 3740 3878
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 3240 2984 3292 2990
rect 4172 2938 4200 3470
rect 4344 3392 4396 3398
rect 4344 3334 4396 3340
rect 4356 3126 4384 3334
rect 4344 3120 4396 3126
rect 4344 3062 4396 3068
rect 3240 2926 3292 2932
rect 2964 2508 3016 2514
rect 2964 2450 3016 2456
rect 2872 1692 2924 1698
rect 2872 1634 2924 1640
rect 2884 1465 2912 1634
rect 2870 1456 2926 1465
rect 2870 1391 2926 1400
rect 3252 800 3280 2926
rect 4080 2910 4200 2938
rect 4080 2514 4108 2910
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 4528 2508 4580 2514
rect 4528 2450 4580 2456
rect 4540 800 4568 2450
rect 4632 2378 4660 3878
rect 4724 3602 4752 4558
rect 4816 3670 4844 4966
rect 4908 3670 4936 22066
rect 5080 14952 5132 14958
rect 5080 14894 5132 14900
rect 5092 14618 5120 14894
rect 5080 14612 5132 14618
rect 5080 14554 5132 14560
rect 5184 13938 5212 26206
rect 5276 26206 5396 26234
rect 5276 24818 5304 26206
rect 5264 24812 5316 24818
rect 5264 24754 5316 24760
rect 5172 13932 5224 13938
rect 5172 13874 5224 13880
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 5000 4554 5028 8910
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5460 4622 5488 7346
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 4988 4548 5040 4554
rect 4988 4490 5040 4496
rect 5356 4480 5408 4486
rect 5356 4422 5408 4428
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 4804 3664 4856 3670
rect 4804 3606 4856 3612
rect 4896 3664 4948 3670
rect 4896 3606 4948 3612
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4908 3534 4936 3606
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 5000 2990 5028 3878
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 4620 2372 4672 2378
rect 4620 2314 4672 2320
rect 5184 800 5212 2926
rect 5368 2310 5396 4422
rect 5356 2304 5408 2310
rect 5356 2246 5408 2252
rect 5552 1698 5580 28562
rect 5828 14414 5856 35866
rect 5908 34604 5960 34610
rect 5908 34546 5960 34552
rect 5920 33658 5948 34546
rect 5908 33652 5960 33658
rect 5908 33594 5960 33600
rect 6000 32904 6052 32910
rect 6000 32846 6052 32852
rect 6012 32570 6040 32846
rect 6000 32564 6052 32570
rect 6000 32506 6052 32512
rect 6104 31278 6132 41074
rect 6552 38208 6604 38214
rect 6552 38150 6604 38156
rect 6564 37874 6592 38150
rect 6552 37868 6604 37874
rect 6552 37810 6604 37816
rect 6184 36168 6236 36174
rect 6184 36110 6236 36116
rect 6196 35834 6224 36110
rect 6184 35828 6236 35834
rect 6184 35770 6236 35776
rect 6748 31890 6776 41386
rect 7116 41274 7144 41482
rect 7104 41268 7156 41274
rect 7104 41210 7156 41216
rect 7392 41138 7420 44950
rect 7380 41132 7432 41138
rect 7380 41074 7432 41080
rect 8208 40112 8260 40118
rect 8208 40054 8260 40060
rect 8116 37868 8168 37874
rect 8116 37810 8168 37816
rect 7932 37664 7984 37670
rect 7932 37606 7984 37612
rect 7944 37466 7972 37606
rect 7932 37460 7984 37466
rect 7932 37402 7984 37408
rect 7104 37256 7156 37262
rect 7104 37198 7156 37204
rect 7116 36106 7144 37198
rect 8128 36174 8156 37810
rect 8116 36168 8168 36174
rect 8116 36110 8168 36116
rect 7104 36100 7156 36106
rect 7104 36042 7156 36048
rect 8128 35894 8156 36110
rect 8036 35866 8156 35894
rect 7104 34944 7156 34950
rect 7104 34886 7156 34892
rect 7012 34400 7064 34406
rect 7012 34342 7064 34348
rect 7024 33998 7052 34342
rect 7012 33992 7064 33998
rect 7012 33934 7064 33940
rect 6828 33856 6880 33862
rect 6828 33798 6880 33804
rect 6840 32910 6868 33798
rect 6828 32904 6880 32910
rect 6828 32846 6880 32852
rect 6920 32428 6972 32434
rect 6920 32370 6972 32376
rect 6736 31884 6788 31890
rect 6736 31826 6788 31832
rect 6552 31680 6604 31686
rect 6552 31622 6604 31628
rect 6564 31346 6592 31622
rect 6932 31414 6960 32370
rect 7012 31884 7064 31890
rect 7012 31826 7064 31832
rect 6920 31408 6972 31414
rect 6920 31350 6972 31356
rect 6552 31340 6604 31346
rect 6552 31282 6604 31288
rect 6092 31272 6144 31278
rect 6092 31214 6144 31220
rect 6460 31272 6512 31278
rect 6460 31214 6512 31220
rect 6092 27396 6144 27402
rect 6092 27338 6144 27344
rect 6104 27130 6132 27338
rect 6092 27124 6144 27130
rect 6092 27066 6144 27072
rect 6472 26234 6500 31214
rect 6564 30190 6592 31282
rect 6932 30802 6960 31350
rect 6920 30796 6972 30802
rect 6920 30738 6972 30744
rect 6552 30184 6604 30190
rect 6552 30126 6604 30132
rect 6736 30048 6788 30054
rect 6736 29990 6788 29996
rect 6748 29714 6776 29990
rect 6828 29844 6880 29850
rect 6828 29786 6880 29792
rect 6736 29708 6788 29714
rect 6736 29650 6788 29656
rect 6840 29170 6868 29786
rect 6920 29572 6972 29578
rect 6920 29514 6972 29520
rect 6932 29306 6960 29514
rect 6920 29300 6972 29306
rect 6920 29242 6972 29248
rect 6828 29164 6880 29170
rect 6828 29106 6880 29112
rect 6840 26234 6868 29106
rect 6920 29028 6972 29034
rect 6920 28970 6972 28976
rect 6932 28626 6960 28970
rect 6920 28620 6972 28626
rect 6920 28562 6972 28568
rect 7024 28014 7052 31826
rect 7116 31822 7144 34886
rect 8036 34746 8064 35866
rect 8116 35488 8168 35494
rect 8116 35430 8168 35436
rect 8128 35086 8156 35430
rect 8116 35080 8168 35086
rect 8116 35022 8168 35028
rect 7748 34740 7800 34746
rect 7748 34682 7800 34688
rect 8024 34740 8076 34746
rect 8024 34682 8076 34688
rect 7760 34610 7788 34682
rect 7748 34604 7800 34610
rect 7748 34546 7800 34552
rect 7288 34536 7340 34542
rect 7288 34478 7340 34484
rect 7300 33998 7328 34478
rect 7288 33992 7340 33998
rect 7288 33934 7340 33940
rect 7760 33930 7788 34546
rect 8036 33998 8064 34682
rect 8128 34542 8156 35022
rect 8116 34536 8168 34542
rect 8116 34478 8168 34484
rect 8024 33992 8076 33998
rect 8024 33934 8076 33940
rect 7748 33924 7800 33930
rect 7748 33866 7800 33872
rect 7380 33856 7432 33862
rect 7380 33798 7432 33804
rect 7392 33522 7420 33798
rect 7760 33590 7788 33866
rect 7748 33584 7800 33590
rect 7748 33526 7800 33532
rect 7196 33516 7248 33522
rect 7196 33458 7248 33464
rect 7380 33516 7432 33522
rect 7380 33458 7432 33464
rect 7208 33046 7236 33458
rect 7196 33040 7248 33046
rect 7196 32982 7248 32988
rect 7104 31816 7156 31822
rect 7104 31758 7156 31764
rect 8024 31408 8076 31414
rect 8024 31350 8076 31356
rect 7104 30728 7156 30734
rect 7104 30670 7156 30676
rect 7116 28626 7144 30670
rect 7104 28620 7156 28626
rect 7104 28562 7156 28568
rect 8036 28558 8064 31350
rect 8220 31278 8248 40054
rect 8312 35222 8340 47126
rect 9048 47054 9076 49200
rect 9036 47048 9088 47054
rect 9036 46990 9088 46996
rect 10508 46368 10560 46374
rect 10508 46310 10560 46316
rect 10520 46034 10548 46310
rect 10980 46034 11008 49200
rect 12440 47048 12492 47054
rect 12440 46990 12492 46996
rect 12452 46646 12480 46990
rect 12440 46640 12492 46646
rect 12440 46582 12492 46588
rect 12912 46594 12940 49200
rect 14200 47122 14228 49200
rect 14188 47116 14240 47122
rect 14188 47058 14240 47064
rect 13820 46980 13872 46986
rect 13820 46922 13872 46928
rect 12912 46566 13032 46594
rect 13004 46510 13032 46566
rect 12900 46504 12952 46510
rect 12900 46446 12952 46452
rect 12992 46504 13044 46510
rect 12992 46446 13044 46452
rect 12912 46170 12940 46446
rect 12992 46368 13044 46374
rect 12992 46310 13044 46316
rect 12900 46164 12952 46170
rect 12900 46106 12952 46112
rect 10508 46028 10560 46034
rect 10508 45970 10560 45976
rect 10968 46028 11020 46034
rect 10968 45970 11020 45976
rect 10692 45892 10744 45898
rect 10692 45834 10744 45840
rect 10704 45626 10732 45834
rect 10692 45620 10744 45626
rect 10692 45562 10744 45568
rect 12532 45416 12584 45422
rect 12532 45358 12584 45364
rect 12544 45286 12572 45358
rect 12532 45280 12584 45286
rect 12532 45222 12584 45228
rect 13004 40118 13032 46310
rect 13832 46170 13860 46922
rect 14844 46510 14872 49200
rect 14372 46504 14424 46510
rect 14372 46446 14424 46452
rect 14556 46504 14608 46510
rect 14556 46446 14608 46452
rect 14832 46504 14884 46510
rect 14832 46446 14884 46452
rect 13820 46164 13872 46170
rect 13820 46106 13872 46112
rect 13268 45960 13320 45966
rect 13268 45902 13320 45908
rect 13280 44470 13308 45902
rect 14384 45490 14412 46446
rect 14568 46170 14596 46446
rect 14556 46164 14608 46170
rect 14556 46106 14608 46112
rect 15488 46034 15516 49200
rect 17420 48226 17448 49200
rect 17420 48198 17540 48226
rect 17408 47184 17460 47190
rect 17408 47126 17460 47132
rect 16856 46368 16908 46374
rect 16856 46310 16908 46316
rect 16868 46034 16896 46310
rect 15476 46028 15528 46034
rect 15476 45970 15528 45976
rect 16856 46028 16908 46034
rect 16856 45970 16908 45976
rect 16672 45892 16724 45898
rect 16672 45834 16724 45840
rect 16684 45490 16712 45834
rect 14372 45484 14424 45490
rect 14372 45426 14424 45432
rect 15108 45484 15160 45490
rect 15108 45426 15160 45432
rect 16672 45484 16724 45490
rect 16672 45426 16724 45432
rect 15120 45082 15148 45426
rect 15108 45076 15160 45082
rect 15108 45018 15160 45024
rect 15120 44538 15148 45018
rect 15108 44532 15160 44538
rect 15108 44474 15160 44480
rect 13268 44464 13320 44470
rect 13268 44406 13320 44412
rect 13084 42628 13136 42634
rect 13084 42570 13136 42576
rect 12992 40112 13044 40118
rect 12992 40054 13044 40060
rect 13096 39914 13124 42570
rect 13084 39908 13136 39914
rect 13084 39850 13136 39856
rect 13096 39438 13124 39850
rect 13084 39432 13136 39438
rect 13084 39374 13136 39380
rect 8484 38344 8536 38350
rect 8484 38286 8536 38292
rect 12900 38344 12952 38350
rect 12900 38286 12952 38292
rect 8496 37874 8524 38286
rect 12808 38276 12860 38282
rect 12808 38218 12860 38224
rect 12820 38010 12848 38218
rect 12808 38004 12860 38010
rect 12808 37946 12860 37952
rect 8484 37868 8536 37874
rect 8484 37810 8536 37816
rect 8484 37664 8536 37670
rect 8484 37606 8536 37612
rect 8496 36786 8524 37606
rect 9128 37120 9180 37126
rect 9128 37062 9180 37068
rect 9140 36854 9168 37062
rect 9128 36848 9180 36854
rect 9128 36790 9180 36796
rect 12912 36786 12940 38286
rect 13176 37120 13228 37126
rect 13176 37062 13228 37068
rect 13188 36854 13216 37062
rect 13176 36848 13228 36854
rect 13176 36790 13228 36796
rect 8484 36780 8536 36786
rect 8484 36722 8536 36728
rect 12900 36780 12952 36786
rect 12900 36722 12952 36728
rect 9220 36576 9272 36582
rect 9220 36518 9272 36524
rect 9232 36378 9260 36518
rect 9220 36372 9272 36378
rect 9220 36314 9272 36320
rect 9220 36168 9272 36174
rect 9220 36110 9272 36116
rect 8300 35216 8352 35222
rect 8300 35158 8352 35164
rect 9232 34474 9260 36110
rect 9588 36100 9640 36106
rect 9588 36042 9640 36048
rect 9600 35698 9628 36042
rect 10048 36032 10100 36038
rect 10048 35974 10100 35980
rect 10060 35766 10088 35974
rect 10048 35760 10100 35766
rect 10048 35702 10100 35708
rect 9588 35692 9640 35698
rect 9588 35634 9640 35640
rect 9680 34740 9732 34746
rect 9680 34682 9732 34688
rect 9220 34468 9272 34474
rect 9220 34410 9272 34416
rect 9232 33522 9260 34410
rect 9404 34400 9456 34406
rect 9404 34342 9456 34348
rect 9416 34066 9444 34342
rect 9404 34060 9456 34066
rect 9404 34002 9456 34008
rect 9692 33998 9720 34682
rect 9772 34536 9824 34542
rect 9772 34478 9824 34484
rect 9680 33992 9732 33998
rect 9680 33934 9732 33940
rect 9784 33658 9812 34478
rect 12440 34400 12492 34406
rect 12440 34342 12492 34348
rect 12452 33998 12480 34342
rect 12072 33992 12124 33998
rect 12072 33934 12124 33940
rect 12440 33992 12492 33998
rect 12440 33934 12492 33940
rect 10324 33856 10376 33862
rect 10324 33798 10376 33804
rect 9772 33652 9824 33658
rect 9772 33594 9824 33600
rect 10336 33522 10364 33798
rect 9220 33516 9272 33522
rect 9220 33458 9272 33464
rect 10324 33516 10376 33522
rect 10324 33458 10376 33464
rect 9232 32910 9260 33458
rect 11704 33312 11756 33318
rect 11704 33254 11756 33260
rect 9404 32972 9456 32978
rect 9404 32914 9456 32920
rect 9220 32904 9272 32910
rect 9220 32846 9272 32852
rect 8944 32360 8996 32366
rect 8944 32302 8996 32308
rect 8956 32026 8984 32302
rect 8944 32020 8996 32026
rect 8944 31962 8996 31968
rect 9416 31958 9444 32914
rect 11716 32910 11744 33254
rect 11704 32904 11756 32910
rect 11704 32846 11756 32852
rect 9772 32768 9824 32774
rect 9772 32710 9824 32716
rect 10324 32768 10376 32774
rect 10324 32710 10376 32716
rect 9404 31952 9456 31958
rect 9404 31894 9456 31900
rect 9220 31816 9272 31822
rect 9220 31758 9272 31764
rect 9232 31414 9260 31758
rect 9220 31408 9272 31414
rect 9220 31350 9272 31356
rect 8208 31272 8260 31278
rect 8208 31214 8260 31220
rect 9232 31226 9260 31350
rect 9232 31198 9352 31226
rect 9220 31136 9272 31142
rect 9220 31078 9272 31084
rect 8392 30592 8444 30598
rect 8392 30534 8444 30540
rect 8404 29238 8432 30534
rect 9232 30258 9260 31078
rect 9324 30734 9352 31198
rect 9312 30728 9364 30734
rect 9312 30670 9364 30676
rect 9416 30580 9444 31894
rect 9784 30802 9812 32710
rect 10336 32570 10364 32710
rect 12084 32570 12112 33934
rect 12256 33856 12308 33862
rect 12256 33798 12308 33804
rect 12348 33856 12400 33862
rect 12348 33798 12400 33804
rect 12268 33590 12296 33798
rect 12256 33584 12308 33590
rect 12256 33526 12308 33532
rect 12164 32768 12216 32774
rect 12164 32710 12216 32716
rect 10324 32564 10376 32570
rect 10324 32506 10376 32512
rect 12072 32564 12124 32570
rect 12072 32506 12124 32512
rect 11060 32428 11112 32434
rect 11060 32370 11112 32376
rect 11072 32026 11100 32370
rect 11888 32360 11940 32366
rect 11888 32302 11940 32308
rect 11060 32020 11112 32026
rect 11060 31962 11112 31968
rect 11900 31822 11928 32302
rect 12176 32298 12204 32710
rect 12164 32292 12216 32298
rect 12164 32234 12216 32240
rect 10600 31816 10652 31822
rect 10600 31758 10652 31764
rect 11888 31816 11940 31822
rect 11888 31758 11940 31764
rect 10324 31136 10376 31142
rect 10324 31078 10376 31084
rect 9772 30796 9824 30802
rect 9772 30738 9824 30744
rect 9324 30552 9444 30580
rect 9220 30252 9272 30258
rect 9220 30194 9272 30200
rect 9324 30054 9352 30552
rect 10336 30326 10364 31078
rect 10324 30320 10376 30326
rect 10324 30262 10376 30268
rect 10612 30122 10640 31758
rect 11704 31340 11756 31346
rect 11704 31282 11756 31288
rect 10784 31136 10836 31142
rect 10784 31078 10836 31084
rect 10796 30734 10824 31078
rect 10784 30728 10836 30734
rect 10784 30670 10836 30676
rect 11716 30394 11744 31282
rect 11704 30388 11756 30394
rect 11704 30330 11756 30336
rect 10600 30116 10652 30122
rect 10600 30058 10652 30064
rect 9312 30048 9364 30054
rect 9312 29990 9364 29996
rect 8392 29232 8444 29238
rect 8392 29174 8444 29180
rect 8116 29096 8168 29102
rect 8116 29038 8168 29044
rect 8128 28762 8156 29038
rect 8116 28756 8168 28762
rect 8116 28698 8168 28704
rect 9324 28558 9352 29990
rect 10612 29646 10640 30058
rect 10600 29640 10652 29646
rect 10600 29582 10652 29588
rect 10232 29504 10284 29510
rect 10232 29446 10284 29452
rect 9496 28960 9548 28966
rect 9496 28902 9548 28908
rect 9508 28626 9536 28902
rect 9496 28620 9548 28626
rect 9496 28562 9548 28568
rect 8024 28552 8076 28558
rect 8024 28494 8076 28500
rect 9312 28552 9364 28558
rect 9312 28494 9364 28500
rect 7196 28076 7248 28082
rect 7196 28018 7248 28024
rect 7012 28008 7064 28014
rect 7012 27950 7064 27956
rect 7208 27606 7236 28018
rect 7196 27600 7248 27606
rect 7196 27542 7248 27548
rect 7932 27532 7984 27538
rect 7932 27474 7984 27480
rect 7944 26994 7972 27474
rect 8036 27402 8064 28494
rect 9128 28416 9180 28422
rect 9128 28358 9180 28364
rect 9140 28082 9168 28358
rect 9128 28076 9180 28082
rect 9128 28018 9180 28024
rect 9220 28076 9272 28082
rect 9220 28018 9272 28024
rect 8208 27940 8260 27946
rect 8208 27882 8260 27888
rect 8024 27396 8076 27402
rect 8024 27338 8076 27344
rect 8036 26994 8064 27338
rect 7932 26988 7984 26994
rect 7932 26930 7984 26936
rect 8024 26988 8076 26994
rect 8024 26930 8076 26936
rect 6472 26206 6592 26234
rect 6460 25832 6512 25838
rect 6460 25774 6512 25780
rect 6472 25498 6500 25774
rect 6460 25492 6512 25498
rect 6460 25434 6512 25440
rect 6564 23730 6592 26206
rect 6748 26206 6868 26234
rect 6644 24132 6696 24138
rect 6644 24074 6696 24080
rect 6656 23866 6684 24074
rect 6644 23860 6696 23866
rect 6644 23802 6696 23808
rect 6552 23724 6604 23730
rect 6552 23666 6604 23672
rect 6748 17678 6776 26206
rect 7944 26042 7972 26930
rect 7932 26036 7984 26042
rect 7932 25978 7984 25984
rect 7104 25900 7156 25906
rect 7104 25842 7156 25848
rect 7116 25498 7144 25842
rect 7104 25492 7156 25498
rect 7104 25434 7156 25440
rect 8036 25362 8064 26930
rect 8024 25356 8076 25362
rect 8024 25298 8076 25304
rect 8036 25226 8064 25298
rect 8024 25220 8076 25226
rect 8024 25162 8076 25168
rect 8036 24818 8064 25162
rect 8024 24812 8076 24818
rect 8024 24754 8076 24760
rect 8220 24206 8248 27882
rect 9036 27872 9088 27878
rect 9036 27814 9088 27820
rect 9048 26994 9076 27814
rect 9232 27606 9260 28018
rect 9220 27600 9272 27606
rect 9220 27542 9272 27548
rect 9324 27062 9352 28494
rect 9956 27532 10008 27538
rect 9956 27474 10008 27480
rect 9312 27056 9364 27062
rect 9312 26998 9364 27004
rect 9036 26988 9088 26994
rect 9036 26930 9088 26936
rect 9324 25430 9352 26998
rect 9968 26586 9996 27474
rect 10244 27470 10272 29446
rect 11900 28490 11928 31758
rect 12360 30802 12388 33798
rect 12348 30796 12400 30802
rect 12348 30738 12400 30744
rect 12452 30666 12480 33934
rect 13176 33516 13228 33522
rect 13176 33458 13228 33464
rect 13188 32434 13216 33458
rect 13176 32428 13228 32434
rect 13176 32370 13228 32376
rect 12532 31204 12584 31210
rect 12532 31146 12584 31152
rect 12440 30660 12492 30666
rect 12440 30602 12492 30608
rect 12164 30592 12216 30598
rect 12544 30546 12572 31146
rect 12900 30660 12952 30666
rect 12900 30602 12952 30608
rect 12164 30534 12216 30540
rect 12176 30190 12204 30534
rect 12452 30518 12572 30546
rect 12164 30184 12216 30190
rect 12164 30126 12216 30132
rect 12176 29714 12204 30126
rect 12452 30122 12480 30518
rect 12912 30394 12940 30602
rect 12900 30388 12952 30394
rect 12900 30330 12952 30336
rect 13084 30252 13136 30258
rect 13084 30194 13136 30200
rect 12440 30116 12492 30122
rect 12440 30058 12492 30064
rect 12452 29714 12480 30058
rect 13096 29782 13124 30194
rect 13084 29776 13136 29782
rect 13084 29718 13136 29724
rect 12164 29708 12216 29714
rect 12164 29650 12216 29656
rect 12440 29708 12492 29714
rect 12440 29650 12492 29656
rect 12624 29504 12676 29510
rect 12624 29446 12676 29452
rect 12164 28688 12216 28694
rect 12164 28630 12216 28636
rect 11888 28484 11940 28490
rect 11888 28426 11940 28432
rect 10600 28008 10652 28014
rect 10600 27950 10652 27956
rect 10612 27606 10640 27950
rect 11796 27872 11848 27878
rect 11796 27814 11848 27820
rect 10600 27600 10652 27606
rect 10600 27542 10652 27548
rect 10232 27464 10284 27470
rect 10232 27406 10284 27412
rect 11808 27402 11836 27814
rect 11796 27396 11848 27402
rect 11796 27338 11848 27344
rect 11808 27130 11836 27338
rect 11796 27124 11848 27130
rect 11796 27066 11848 27072
rect 10140 26784 10192 26790
rect 10140 26726 10192 26732
rect 9956 26580 10008 26586
rect 9956 26522 10008 26528
rect 10152 26450 10180 26726
rect 10140 26444 10192 26450
rect 10140 26386 10192 26392
rect 9588 26376 9640 26382
rect 9588 26318 9640 26324
rect 9312 25424 9364 25430
rect 9312 25366 9364 25372
rect 8576 25220 8628 25226
rect 8576 25162 8628 25168
rect 8588 24274 8616 25162
rect 8852 24812 8904 24818
rect 8852 24754 8904 24760
rect 8576 24268 8628 24274
rect 8576 24210 8628 24216
rect 8208 24200 8260 24206
rect 8208 24142 8260 24148
rect 8864 23866 8892 24754
rect 9324 24750 9352 25366
rect 9600 25362 9628 26318
rect 10152 26234 10180 26386
rect 10152 26206 10272 26234
rect 9588 25356 9640 25362
rect 9588 25298 9640 25304
rect 9600 24954 9628 25298
rect 9588 24948 9640 24954
rect 9588 24890 9640 24896
rect 10244 24818 10272 26206
rect 11612 25220 11664 25226
rect 11612 25162 11664 25168
rect 11624 24954 11652 25162
rect 11612 24948 11664 24954
rect 11612 24890 11664 24896
rect 10232 24812 10284 24818
rect 10232 24754 10284 24760
rect 11796 24812 11848 24818
rect 11796 24754 11848 24760
rect 9312 24744 9364 24750
rect 9312 24686 9364 24692
rect 8852 23860 8904 23866
rect 8852 23802 8904 23808
rect 9324 23662 9352 24686
rect 11152 24608 11204 24614
rect 11152 24550 11204 24556
rect 11164 24206 11192 24550
rect 11808 24410 11836 24754
rect 11796 24404 11848 24410
rect 11796 24346 11848 24352
rect 11152 24200 11204 24206
rect 11152 24142 11204 24148
rect 10140 24064 10192 24070
rect 10140 24006 10192 24012
rect 10152 23866 10180 24006
rect 10140 23860 10192 23866
rect 10140 23802 10192 23808
rect 11704 23724 11756 23730
rect 11704 23666 11756 23672
rect 9312 23656 9364 23662
rect 9312 23598 9364 23604
rect 11716 23118 11744 23666
rect 11704 23112 11756 23118
rect 11704 23054 11756 23060
rect 11612 22976 11664 22982
rect 11612 22918 11664 22924
rect 7564 22636 7616 22642
rect 7564 22578 7616 22584
rect 11428 22636 11480 22642
rect 11428 22578 11480 22584
rect 6736 17672 6788 17678
rect 6736 17614 6788 17620
rect 6000 15496 6052 15502
rect 6000 15438 6052 15444
rect 6012 15026 6040 15438
rect 6000 15020 6052 15026
rect 6000 14962 6052 14968
rect 5816 14408 5868 14414
rect 5816 14350 5868 14356
rect 5828 4146 5856 14350
rect 7576 4146 7604 22578
rect 11440 22098 11468 22578
rect 11624 22166 11652 22918
rect 11716 22778 11744 23054
rect 11704 22772 11756 22778
rect 11704 22714 11756 22720
rect 11612 22160 11664 22166
rect 11612 22102 11664 22108
rect 11900 22098 11928 28426
rect 12176 27674 12204 28630
rect 12636 28218 12664 29446
rect 13280 29306 13308 44406
rect 14740 40520 14792 40526
rect 14740 40462 14792 40468
rect 14648 39976 14700 39982
rect 14648 39918 14700 39924
rect 14660 39642 14688 39918
rect 14648 39636 14700 39642
rect 14648 39578 14700 39584
rect 14752 38962 14780 40462
rect 16028 40452 16080 40458
rect 16028 40394 16080 40400
rect 16040 40186 16068 40394
rect 16028 40180 16080 40186
rect 16028 40122 16080 40128
rect 14924 39976 14976 39982
rect 14924 39918 14976 39924
rect 16948 39976 17000 39982
rect 16948 39918 17000 39924
rect 14936 38962 14964 39918
rect 16028 39500 16080 39506
rect 16028 39442 16080 39448
rect 16040 38962 16068 39442
rect 16960 38962 16988 39918
rect 14740 38956 14792 38962
rect 14740 38898 14792 38904
rect 14924 38956 14976 38962
rect 14924 38898 14976 38904
rect 16028 38956 16080 38962
rect 16028 38898 16080 38904
rect 16948 38956 17000 38962
rect 16948 38898 17000 38904
rect 14280 38548 14332 38554
rect 14280 38490 14332 38496
rect 14292 37806 14320 38490
rect 14752 37942 14780 38898
rect 14832 38888 14884 38894
rect 14832 38830 14884 38836
rect 14844 38214 14872 38830
rect 14936 38554 14964 38898
rect 15016 38752 15068 38758
rect 15016 38694 15068 38700
rect 15936 38752 15988 38758
rect 15936 38694 15988 38700
rect 14924 38548 14976 38554
rect 14924 38490 14976 38496
rect 15028 38350 15056 38694
rect 15108 38480 15160 38486
rect 15108 38422 15160 38428
rect 15016 38344 15068 38350
rect 15016 38286 15068 38292
rect 14832 38208 14884 38214
rect 14832 38150 14884 38156
rect 14740 37936 14792 37942
rect 14740 37878 14792 37884
rect 13820 37800 13872 37806
rect 13820 37742 13872 37748
rect 14280 37800 14332 37806
rect 14280 37742 14332 37748
rect 13832 37330 13860 37742
rect 13820 37324 13872 37330
rect 13820 37266 13872 37272
rect 14556 37324 14608 37330
rect 14556 37266 14608 37272
rect 13832 36922 13860 37266
rect 13820 36916 13872 36922
rect 13820 36858 13872 36864
rect 14096 35828 14148 35834
rect 14096 35770 14148 35776
rect 14004 35488 14056 35494
rect 14004 35430 14056 35436
rect 13728 34672 13780 34678
rect 13728 34614 13780 34620
rect 13740 33522 13768 34614
rect 14016 34610 14044 35430
rect 14004 34604 14056 34610
rect 14004 34546 14056 34552
rect 14108 34202 14136 35770
rect 14568 35698 14596 37266
rect 14752 37262 14780 37878
rect 14844 37874 14872 38150
rect 14832 37868 14884 37874
rect 14832 37810 14884 37816
rect 14844 37754 14872 37810
rect 14844 37726 14964 37754
rect 14936 37262 14964 37726
rect 15028 37262 15056 38286
rect 15120 37874 15148 38422
rect 15660 38344 15712 38350
rect 15660 38286 15712 38292
rect 15108 37868 15160 37874
rect 15108 37810 15160 37816
rect 15108 37664 15160 37670
rect 15108 37606 15160 37612
rect 14740 37256 14792 37262
rect 14740 37198 14792 37204
rect 14924 37256 14976 37262
rect 14924 37198 14976 37204
rect 15016 37256 15068 37262
rect 15016 37198 15068 37204
rect 14752 36854 14780 37198
rect 14936 37126 14964 37198
rect 15120 37194 15148 37606
rect 15108 37188 15160 37194
rect 15108 37130 15160 37136
rect 14924 37120 14976 37126
rect 14924 37062 14976 37068
rect 14740 36848 14792 36854
rect 14740 36790 14792 36796
rect 14752 36650 14780 36790
rect 14936 36786 14964 37062
rect 14924 36780 14976 36786
rect 14924 36722 14976 36728
rect 14740 36644 14792 36650
rect 14740 36586 14792 36592
rect 14556 35692 14608 35698
rect 14556 35634 14608 35640
rect 14464 35488 14516 35494
rect 14464 35430 14516 35436
rect 14476 34746 14504 35430
rect 15672 35154 15700 38286
rect 15844 38276 15896 38282
rect 15844 38218 15896 38224
rect 15856 38010 15884 38218
rect 15844 38004 15896 38010
rect 15844 37946 15896 37952
rect 15948 37874 15976 38694
rect 16960 38554 16988 38898
rect 16948 38548 17000 38554
rect 16948 38490 17000 38496
rect 16960 38214 16988 38490
rect 16948 38208 17000 38214
rect 16948 38150 17000 38156
rect 16960 37942 16988 38150
rect 16948 37936 17000 37942
rect 16948 37878 17000 37884
rect 15936 37868 15988 37874
rect 15936 37810 15988 37816
rect 15948 35766 15976 37810
rect 16960 37398 16988 37878
rect 16948 37392 17000 37398
rect 16948 37334 17000 37340
rect 17040 37188 17092 37194
rect 17040 37130 17092 37136
rect 16488 36712 16540 36718
rect 16488 36654 16540 36660
rect 15936 35760 15988 35766
rect 15936 35702 15988 35708
rect 15660 35148 15712 35154
rect 15660 35090 15712 35096
rect 14464 34740 14516 34746
rect 14464 34682 14516 34688
rect 15672 34542 15700 35090
rect 15384 34536 15436 34542
rect 15384 34478 15436 34484
rect 15660 34536 15712 34542
rect 15660 34478 15712 34484
rect 14096 34196 14148 34202
rect 14096 34138 14148 34144
rect 15396 34066 15424 34478
rect 15384 34060 15436 34066
rect 15384 34002 15436 34008
rect 13728 33516 13780 33522
rect 13728 33458 13780 33464
rect 15396 32978 15424 34002
rect 15384 32972 15436 32978
rect 15384 32914 15436 32920
rect 14280 32904 14332 32910
rect 14280 32846 14332 32852
rect 13544 32768 13596 32774
rect 13544 32710 13596 32716
rect 13556 32502 13584 32710
rect 13544 32496 13596 32502
rect 13544 32438 13596 32444
rect 14292 32026 14320 32846
rect 14832 32836 14884 32842
rect 14832 32778 14884 32784
rect 14556 32564 14608 32570
rect 14556 32506 14608 32512
rect 14280 32020 14332 32026
rect 14280 31962 14332 31968
rect 14568 31754 14596 32506
rect 14556 31748 14608 31754
rect 14556 31690 14608 31696
rect 13544 31272 13596 31278
rect 13544 31214 13596 31220
rect 13556 30938 13584 31214
rect 13544 30932 13596 30938
rect 13544 30874 13596 30880
rect 14280 29640 14332 29646
rect 14280 29582 14332 29588
rect 14740 29640 14792 29646
rect 14740 29582 14792 29588
rect 13268 29300 13320 29306
rect 13268 29242 13320 29248
rect 12716 29028 12768 29034
rect 12716 28970 12768 28976
rect 12728 28422 12756 28970
rect 13544 28960 13596 28966
rect 13544 28902 13596 28908
rect 13556 28490 13584 28902
rect 14292 28762 14320 29582
rect 14464 29504 14516 29510
rect 14464 29446 14516 29452
rect 14476 29238 14504 29446
rect 14464 29232 14516 29238
rect 14464 29174 14516 29180
rect 14752 29102 14780 29582
rect 14740 29096 14792 29102
rect 14740 29038 14792 29044
rect 14280 28756 14332 28762
rect 14280 28698 14332 28704
rect 13728 28620 13780 28626
rect 13728 28562 13780 28568
rect 13544 28484 13596 28490
rect 13544 28426 13596 28432
rect 12716 28416 12768 28422
rect 12716 28358 12768 28364
rect 12900 28416 12952 28422
rect 12900 28358 12952 28364
rect 12624 28212 12676 28218
rect 12624 28154 12676 28160
rect 12912 28150 12940 28358
rect 12900 28144 12952 28150
rect 12900 28086 12952 28092
rect 12164 27668 12216 27674
rect 12164 27610 12216 27616
rect 12532 27532 12584 27538
rect 12532 27474 12584 27480
rect 12256 26376 12308 26382
rect 12256 26318 12308 26324
rect 12072 26240 12124 26246
rect 12072 26182 12124 26188
rect 12084 25974 12112 26182
rect 12072 25968 12124 25974
rect 12072 25910 12124 25916
rect 12268 25498 12296 26318
rect 12440 25696 12492 25702
rect 12440 25638 12492 25644
rect 12256 25492 12308 25498
rect 12256 25434 12308 25440
rect 12452 24886 12480 25638
rect 12544 25362 12572 27474
rect 12900 27328 12952 27334
rect 12900 27270 12952 27276
rect 12532 25356 12584 25362
rect 12532 25298 12584 25304
rect 12440 24880 12492 24886
rect 12440 24822 12492 24828
rect 12544 24698 12572 25298
rect 12624 25152 12676 25158
rect 12624 25094 12676 25100
rect 12452 24670 12572 24698
rect 12348 24608 12400 24614
rect 12348 24550 12400 24556
rect 12360 24138 12388 24550
rect 12452 24274 12480 24670
rect 12440 24268 12492 24274
rect 12440 24210 12492 24216
rect 12348 24132 12400 24138
rect 12348 24074 12400 24080
rect 12452 23186 12480 24210
rect 12440 23180 12492 23186
rect 12440 23122 12492 23128
rect 11428 22092 11480 22098
rect 11428 22034 11480 22040
rect 11888 22092 11940 22098
rect 11888 22034 11940 22040
rect 11900 21690 11928 22034
rect 11888 21684 11940 21690
rect 11888 21626 11940 21632
rect 12532 20460 12584 20466
rect 12532 20402 12584 20408
rect 12164 20256 12216 20262
rect 12164 20198 12216 20204
rect 12176 19786 12204 20198
rect 12164 19780 12216 19786
rect 12164 19722 12216 19728
rect 12256 19780 12308 19786
rect 12256 19722 12308 19728
rect 12268 17678 12296 19722
rect 12544 19514 12572 20402
rect 12532 19508 12584 19514
rect 12532 19450 12584 19456
rect 12636 19174 12664 25094
rect 12808 22976 12860 22982
rect 12808 22918 12860 22924
rect 12716 20460 12768 20466
rect 12716 20402 12768 20408
rect 12624 19168 12676 19174
rect 12624 19110 12676 19116
rect 12636 18306 12664 19110
rect 12452 18278 12664 18306
rect 12072 17672 12124 17678
rect 12072 17614 12124 17620
rect 12256 17672 12308 17678
rect 12256 17614 12308 17620
rect 12084 17542 12112 17614
rect 11980 17536 12032 17542
rect 11980 17478 12032 17484
rect 12072 17536 12124 17542
rect 12072 17478 12124 17484
rect 11992 17202 12020 17478
rect 12268 17270 12296 17614
rect 12256 17264 12308 17270
rect 12256 17206 12308 17212
rect 11980 17196 12032 17202
rect 11980 17138 12032 17144
rect 12268 13938 12296 17206
rect 12256 13932 12308 13938
rect 12256 13874 12308 13880
rect 12452 12434 12480 18278
rect 12636 18222 12664 18278
rect 12532 18216 12584 18222
rect 12532 18158 12584 18164
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 12544 17610 12572 18158
rect 12728 18086 12756 20402
rect 12820 20398 12848 22918
rect 12808 20392 12860 20398
rect 12808 20334 12860 20340
rect 12820 20058 12848 20334
rect 12808 20052 12860 20058
rect 12808 19994 12860 20000
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 12728 17898 12756 18022
rect 12636 17882 12756 17898
rect 12624 17876 12756 17882
rect 12676 17870 12756 17876
rect 12624 17818 12676 17824
rect 12532 17604 12584 17610
rect 12532 17546 12584 17552
rect 12452 12406 12664 12434
rect 12532 5228 12584 5234
rect 12532 5170 12584 5176
rect 12544 4146 12572 5170
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 7196 4004 7248 4010
rect 7196 3946 7248 3952
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 6104 3602 6132 3878
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 5540 1692 5592 1698
rect 5540 1634 5592 1640
rect 6472 800 6500 3538
rect 6644 2848 6696 2854
rect 6644 2790 6696 2796
rect 6656 2514 6684 2790
rect 6840 2514 6868 3878
rect 7208 3738 7236 3946
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 7196 3732 7248 3738
rect 7196 3674 7248 3680
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7484 3058 7512 3470
rect 7668 3126 7696 3878
rect 10704 3602 10732 3878
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 10508 3528 10560 3534
rect 10508 3470 10560 3476
rect 7656 3120 7708 3126
rect 7656 3062 7708 3068
rect 10520 3058 10548 3470
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 6644 2508 6696 2514
rect 6644 2450 6696 2456
rect 6828 2508 6880 2514
rect 6828 2450 6880 2456
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 7116 800 7144 2450
rect 7760 800 7788 2926
rect 10980 800 11008 3538
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 11624 800 11652 2994
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12452 2514 12480 2790
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 12544 2378 12572 3878
rect 12636 2650 12664 12406
rect 12820 3738 12848 19994
rect 12912 17678 12940 27270
rect 13084 25696 13136 25702
rect 13084 25638 13136 25644
rect 13096 25294 13124 25638
rect 13084 25288 13136 25294
rect 13084 25230 13136 25236
rect 13556 24954 13584 28426
rect 13740 27538 13768 28562
rect 14648 28552 14700 28558
rect 14648 28494 14700 28500
rect 13728 27532 13780 27538
rect 13728 27474 13780 27480
rect 14556 27464 14608 27470
rect 14556 27406 14608 27412
rect 14372 27328 14424 27334
rect 14372 27270 14424 27276
rect 14384 26994 14412 27270
rect 14372 26988 14424 26994
rect 14372 26930 14424 26936
rect 13636 26920 13688 26926
rect 13636 26862 13688 26868
rect 13544 24948 13596 24954
rect 13544 24890 13596 24896
rect 12992 24812 13044 24818
rect 12992 24754 13044 24760
rect 13004 24410 13032 24754
rect 13648 24750 13676 26862
rect 14568 26586 14596 27406
rect 14556 26580 14608 26586
rect 14556 26522 14608 26528
rect 14556 26376 14608 26382
rect 14556 26318 14608 26324
rect 13636 24744 13688 24750
rect 13636 24686 13688 24692
rect 12992 24404 13044 24410
rect 12992 24346 13044 24352
rect 13648 23662 13676 24686
rect 13912 24608 13964 24614
rect 13912 24550 13964 24556
rect 13924 24206 13952 24550
rect 14568 24342 14596 26318
rect 14556 24336 14608 24342
rect 14556 24278 14608 24284
rect 14568 24206 14596 24278
rect 13912 24200 13964 24206
rect 13912 24142 13964 24148
rect 14556 24200 14608 24206
rect 14556 24142 14608 24148
rect 14464 24064 14516 24070
rect 14464 24006 14516 24012
rect 14280 23724 14332 23730
rect 14280 23666 14332 23672
rect 13084 23656 13136 23662
rect 13084 23598 13136 23604
rect 13636 23656 13688 23662
rect 13636 23598 13688 23604
rect 13096 22574 13124 23598
rect 14292 23322 14320 23666
rect 14280 23316 14332 23322
rect 14280 23258 14332 23264
rect 14476 23118 14504 24006
rect 14464 23112 14516 23118
rect 14464 23054 14516 23060
rect 13084 22568 13136 22574
rect 13084 22510 13136 22516
rect 13096 22098 13124 22510
rect 13084 22092 13136 22098
rect 13084 22034 13136 22040
rect 13096 21554 13124 22034
rect 14464 22024 14516 22030
rect 14464 21966 14516 21972
rect 14280 21888 14332 21894
rect 14280 21830 14332 21836
rect 14292 21622 14320 21830
rect 14280 21616 14332 21622
rect 14280 21558 14332 21564
rect 13084 21548 13136 21554
rect 13084 21490 13136 21496
rect 14476 21146 14504 21966
rect 14464 21140 14516 21146
rect 14464 21082 14516 21088
rect 13820 21004 13872 21010
rect 13820 20946 13872 20952
rect 13452 19712 13504 19718
rect 13452 19654 13504 19660
rect 13360 19440 13412 19446
rect 13360 19382 13412 19388
rect 13372 18290 13400 19382
rect 13464 19378 13492 19654
rect 13452 19372 13504 19378
rect 13452 19314 13504 19320
rect 13832 19310 13860 20946
rect 14568 20942 14596 24142
rect 14660 23254 14688 28494
rect 14752 28082 14780 29038
rect 14740 28076 14792 28082
rect 14740 28018 14792 28024
rect 14844 27606 14872 32778
rect 15016 32224 15068 32230
rect 15016 32166 15068 32172
rect 15028 31958 15056 32166
rect 15396 32026 15424 32914
rect 15568 32904 15620 32910
rect 15568 32846 15620 32852
rect 15580 32366 15608 32846
rect 15568 32360 15620 32366
rect 15568 32302 15620 32308
rect 15384 32020 15436 32026
rect 15384 31962 15436 31968
rect 15016 31952 15068 31958
rect 15016 31894 15068 31900
rect 15292 31816 15344 31822
rect 15292 31758 15344 31764
rect 15304 31414 15332 31758
rect 15660 31748 15712 31754
rect 15660 31690 15712 31696
rect 15292 31408 15344 31414
rect 15292 31350 15344 31356
rect 15672 30938 15700 31690
rect 16500 31346 16528 36654
rect 17052 36174 17080 37130
rect 17316 36644 17368 36650
rect 17316 36586 17368 36592
rect 17328 36378 17356 36586
rect 17316 36372 17368 36378
rect 17316 36314 17368 36320
rect 17040 36168 17092 36174
rect 17040 36110 17092 36116
rect 16672 35080 16724 35086
rect 16672 35022 16724 35028
rect 16580 34944 16632 34950
rect 16580 34886 16632 34892
rect 16592 34746 16620 34886
rect 16580 34740 16632 34746
rect 16580 34682 16632 34688
rect 16684 34610 16712 35022
rect 16856 35012 16908 35018
rect 16856 34954 16908 34960
rect 17224 35012 17276 35018
rect 17224 34954 17276 34960
rect 16868 34746 16896 34954
rect 17132 34944 17184 34950
rect 17132 34886 17184 34892
rect 16856 34740 16908 34746
rect 16856 34682 16908 34688
rect 17144 34610 17172 34886
rect 16672 34604 16724 34610
rect 16672 34546 16724 34552
rect 17132 34604 17184 34610
rect 17132 34546 17184 34552
rect 17236 33318 17264 34954
rect 17328 33930 17356 36314
rect 17316 33924 17368 33930
rect 17316 33866 17368 33872
rect 17224 33312 17276 33318
rect 17224 33254 17276 33260
rect 17236 32434 17264 33254
rect 17224 32428 17276 32434
rect 17224 32370 17276 32376
rect 17328 31754 17356 33866
rect 17420 32570 17448 47126
rect 17512 47054 17540 48198
rect 19352 47054 19380 49200
rect 20444 47184 20496 47190
rect 20444 47126 20496 47132
rect 17500 47048 17552 47054
rect 17500 46990 17552 46996
rect 19340 47048 19392 47054
rect 19340 46990 19392 46996
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 19248 46368 19300 46374
rect 19248 46310 19300 46316
rect 19064 40520 19116 40526
rect 19064 40462 19116 40468
rect 17776 40384 17828 40390
rect 17776 40326 17828 40332
rect 17788 40118 17816 40326
rect 17776 40112 17828 40118
rect 17776 40054 17828 40060
rect 19076 39914 19104 40462
rect 19260 39982 19288 46310
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 20456 41414 20484 47126
rect 22468 47048 22520 47054
rect 22468 46990 22520 46996
rect 22480 46578 22508 46990
rect 22468 46572 22520 46578
rect 22468 46514 22520 46520
rect 23216 46510 23244 49200
rect 23860 47054 23888 49200
rect 24676 47184 24728 47190
rect 24676 47126 24728 47132
rect 23848 47048 23900 47054
rect 23848 46990 23900 46996
rect 22652 46504 22704 46510
rect 22652 46446 22704 46452
rect 23204 46504 23256 46510
rect 23204 46446 23256 46452
rect 22664 46170 22692 46446
rect 22652 46164 22704 46170
rect 22652 46106 22704 46112
rect 24584 45960 24636 45966
rect 24584 45902 24636 45908
rect 22560 45824 22612 45830
rect 22560 45766 22612 45772
rect 22572 45422 22600 45766
rect 24596 45490 24624 45902
rect 24584 45484 24636 45490
rect 24584 45426 24636 45432
rect 22560 45416 22612 45422
rect 22560 45358 22612 45364
rect 20456 41386 20576 41414
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 19248 39976 19300 39982
rect 19248 39918 19300 39924
rect 19064 39908 19116 39914
rect 19064 39850 19116 39856
rect 18880 38956 18932 38962
rect 18880 38898 18932 38904
rect 18052 38888 18104 38894
rect 18052 38830 18104 38836
rect 17960 38752 18012 38758
rect 17960 38694 18012 38700
rect 17972 37874 18000 38694
rect 17960 37868 18012 37874
rect 17960 37810 18012 37816
rect 17972 37330 18000 37810
rect 17960 37324 18012 37330
rect 17960 37266 18012 37272
rect 17960 35624 18012 35630
rect 17960 35566 18012 35572
rect 17684 35556 17736 35562
rect 17684 35498 17736 35504
rect 17500 35148 17552 35154
rect 17500 35090 17552 35096
rect 17512 34678 17540 35090
rect 17696 35086 17724 35498
rect 17972 35222 18000 35566
rect 18064 35494 18092 38830
rect 18892 38554 18920 38898
rect 18880 38548 18932 38554
rect 18880 38490 18932 38496
rect 18696 38276 18748 38282
rect 18696 38218 18748 38224
rect 18708 38010 18736 38218
rect 18696 38004 18748 38010
rect 18696 37946 18748 37952
rect 18892 37942 18920 38490
rect 18880 37936 18932 37942
rect 18880 37878 18932 37884
rect 18972 37936 19024 37942
rect 18972 37878 19024 37884
rect 18236 37868 18288 37874
rect 18236 37810 18288 37816
rect 18144 37732 18196 37738
rect 18144 37674 18196 37680
rect 18052 35488 18104 35494
rect 18052 35430 18104 35436
rect 17960 35216 18012 35222
rect 17960 35158 18012 35164
rect 17684 35080 17736 35086
rect 17684 35022 17736 35028
rect 17500 34672 17552 34678
rect 17500 34614 17552 34620
rect 17512 34202 17540 34614
rect 17500 34196 17552 34202
rect 17500 34138 17552 34144
rect 17512 33998 17540 34138
rect 17500 33992 17552 33998
rect 17500 33934 17552 33940
rect 17696 33454 17724 35022
rect 17972 34542 18000 35158
rect 18064 35086 18092 35430
rect 18052 35080 18104 35086
rect 18052 35022 18104 35028
rect 18156 34610 18184 37674
rect 18248 37466 18276 37810
rect 18604 37800 18656 37806
rect 18604 37742 18656 37748
rect 18236 37460 18288 37466
rect 18236 37402 18288 37408
rect 18616 37262 18644 37742
rect 18984 37330 19012 37878
rect 18972 37324 19024 37330
rect 18972 37266 19024 37272
rect 18604 37256 18656 37262
rect 18604 37198 18656 37204
rect 18616 37126 18644 37198
rect 18604 37120 18656 37126
rect 18604 37062 18656 37068
rect 18236 36780 18288 36786
rect 18236 36722 18288 36728
rect 18144 34604 18196 34610
rect 18144 34546 18196 34552
rect 17960 34536 18012 34542
rect 17960 34478 18012 34484
rect 17788 34134 17816 34165
rect 17776 34128 17828 34134
rect 18144 34128 18196 34134
rect 17828 34076 18000 34082
rect 17776 34070 18000 34076
rect 18144 34070 18196 34076
rect 17788 34054 18000 34070
rect 17788 33998 17816 34054
rect 17776 33992 17828 33998
rect 17776 33934 17828 33940
rect 17776 33856 17828 33862
rect 17776 33798 17828 33804
rect 17788 33590 17816 33798
rect 17776 33584 17828 33590
rect 17776 33526 17828 33532
rect 17684 33448 17736 33454
rect 17684 33390 17736 33396
rect 17972 33386 18000 34054
rect 18156 33590 18184 34070
rect 18144 33584 18196 33590
rect 18144 33526 18196 33532
rect 18052 33516 18104 33522
rect 18052 33458 18104 33464
rect 17960 33380 18012 33386
rect 17960 33322 18012 33328
rect 18064 32570 18092 33458
rect 18144 33312 18196 33318
rect 18144 33254 18196 33260
rect 17408 32564 17460 32570
rect 17408 32506 17460 32512
rect 18052 32564 18104 32570
rect 18052 32506 18104 32512
rect 18156 32434 18184 33254
rect 18144 32428 18196 32434
rect 18144 32370 18196 32376
rect 17592 32360 17644 32366
rect 17592 32302 17644 32308
rect 17604 31890 17632 32302
rect 17592 31884 17644 31890
rect 17644 31844 17816 31872
rect 17592 31826 17644 31832
rect 17328 31726 17632 31754
rect 16580 31680 16632 31686
rect 16580 31622 16632 31628
rect 17040 31680 17092 31686
rect 17040 31622 17092 31628
rect 16592 31482 16620 31622
rect 16580 31476 16632 31482
rect 16580 31418 16632 31424
rect 16488 31340 16540 31346
rect 16488 31282 16540 31288
rect 17052 31210 17080 31622
rect 17040 31204 17092 31210
rect 17040 31146 17092 31152
rect 17500 31204 17552 31210
rect 17500 31146 17552 31152
rect 15936 31136 15988 31142
rect 15936 31078 15988 31084
rect 15660 30932 15712 30938
rect 15660 30874 15712 30880
rect 15948 30734 15976 31078
rect 15936 30728 15988 30734
rect 15936 30670 15988 30676
rect 16580 30592 16632 30598
rect 16580 30534 16632 30540
rect 15476 30252 15528 30258
rect 15476 30194 15528 30200
rect 15384 30048 15436 30054
rect 15384 29990 15436 29996
rect 15396 29578 15424 29990
rect 15384 29572 15436 29578
rect 15384 29514 15436 29520
rect 15488 29306 15516 30194
rect 16592 30190 16620 30534
rect 16580 30184 16632 30190
rect 16580 30126 16632 30132
rect 17512 29782 17540 31146
rect 17500 29776 17552 29782
rect 17500 29718 17552 29724
rect 17224 29504 17276 29510
rect 17224 29446 17276 29452
rect 15476 29300 15528 29306
rect 15476 29242 15528 29248
rect 15660 29300 15712 29306
rect 15660 29242 15712 29248
rect 15672 29170 15700 29242
rect 15660 29164 15712 29170
rect 15660 29106 15712 29112
rect 16856 29164 16908 29170
rect 16856 29106 16908 29112
rect 16868 28762 16896 29106
rect 16856 28756 16908 28762
rect 16856 28698 16908 28704
rect 17236 28558 17264 29446
rect 17224 28552 17276 28558
rect 17224 28494 17276 28500
rect 17132 28212 17184 28218
rect 17132 28154 17184 28160
rect 14832 27600 14884 27606
rect 14832 27542 14884 27548
rect 14844 27470 14872 27542
rect 15016 27532 15068 27538
rect 15016 27474 15068 27480
rect 14832 27464 14884 27470
rect 14832 27406 14884 27412
rect 15028 27402 15056 27474
rect 15016 27396 15068 27402
rect 15016 27338 15068 27344
rect 14924 26376 14976 26382
rect 14924 26318 14976 26324
rect 14832 25152 14884 25158
rect 14832 25094 14884 25100
rect 14844 24886 14872 25094
rect 14832 24880 14884 24886
rect 14832 24822 14884 24828
rect 14740 24268 14792 24274
rect 14740 24210 14792 24216
rect 14648 23248 14700 23254
rect 14648 23190 14700 23196
rect 14648 23112 14700 23118
rect 14648 23054 14700 23060
rect 14660 22234 14688 23054
rect 14648 22228 14700 22234
rect 14648 22170 14700 22176
rect 14556 20936 14608 20942
rect 14476 20896 14556 20924
rect 14476 19446 14504 20896
rect 14556 20878 14608 20884
rect 14660 20602 14688 22170
rect 14752 22030 14780 24210
rect 14936 24206 14964 26318
rect 14924 24200 14976 24206
rect 14924 24142 14976 24148
rect 14740 22024 14792 22030
rect 14740 21966 14792 21972
rect 14936 21146 14964 24142
rect 15028 23118 15056 27338
rect 16212 26988 16264 26994
rect 16212 26930 16264 26936
rect 15200 26784 15252 26790
rect 15200 26726 15252 26732
rect 15212 26382 15240 26726
rect 16224 26382 16252 26930
rect 17144 26926 17172 28154
rect 17408 28076 17460 28082
rect 17408 28018 17460 28024
rect 17420 27674 17448 28018
rect 17408 27668 17460 27674
rect 17408 27610 17460 27616
rect 17604 27606 17632 31726
rect 17788 29714 17816 31844
rect 17960 31680 18012 31686
rect 17960 31622 18012 31628
rect 17972 31346 18000 31622
rect 17960 31340 18012 31346
rect 17960 31282 18012 31288
rect 17868 31136 17920 31142
rect 17868 31078 17920 31084
rect 17880 30734 17908 31078
rect 17868 30728 17920 30734
rect 17868 30670 17920 30676
rect 17868 30184 17920 30190
rect 17868 30126 17920 30132
rect 17776 29708 17828 29714
rect 17776 29650 17828 29656
rect 17788 28762 17816 29650
rect 17880 29578 17908 30126
rect 17868 29572 17920 29578
rect 17868 29514 17920 29520
rect 17776 28756 17828 28762
rect 17776 28698 17828 28704
rect 17788 28626 17816 28698
rect 17776 28620 17828 28626
rect 17776 28562 17828 28568
rect 18248 28558 18276 36722
rect 18420 34604 18472 34610
rect 18420 34546 18472 34552
rect 18604 34604 18656 34610
rect 18604 34546 18656 34552
rect 18788 34604 18840 34610
rect 18788 34546 18840 34552
rect 18432 34490 18460 34546
rect 18432 34462 18552 34490
rect 18420 34400 18472 34406
rect 18420 34342 18472 34348
rect 18432 34066 18460 34342
rect 18420 34060 18472 34066
rect 18420 34002 18472 34008
rect 18524 33998 18552 34462
rect 18512 33992 18564 33998
rect 18512 33934 18564 33940
rect 18524 33522 18552 33934
rect 18616 33844 18644 34546
rect 18800 33998 18828 34546
rect 18880 34536 18932 34542
rect 18880 34478 18932 34484
rect 18892 34202 18920 34478
rect 18880 34196 18932 34202
rect 18880 34138 18932 34144
rect 18788 33992 18840 33998
rect 18788 33934 18840 33940
rect 18696 33856 18748 33862
rect 18616 33816 18696 33844
rect 18696 33798 18748 33804
rect 18512 33516 18564 33522
rect 18512 33458 18564 33464
rect 18708 33386 18736 33798
rect 18800 33658 18828 33934
rect 18788 33652 18840 33658
rect 18788 33594 18840 33600
rect 18512 33380 18564 33386
rect 18512 33322 18564 33328
rect 18696 33380 18748 33386
rect 18696 33322 18748 33328
rect 18328 32836 18380 32842
rect 18328 32778 18380 32784
rect 18340 30326 18368 32778
rect 18420 30728 18472 30734
rect 18420 30670 18472 30676
rect 18328 30320 18380 30326
rect 18328 30262 18380 30268
rect 18340 30122 18368 30262
rect 18432 30190 18460 30670
rect 18420 30184 18472 30190
rect 18420 30126 18472 30132
rect 18328 30116 18380 30122
rect 18328 30058 18380 30064
rect 18432 29646 18460 30126
rect 18420 29640 18472 29646
rect 18420 29582 18472 29588
rect 18524 29458 18552 33322
rect 18604 29640 18656 29646
rect 18604 29582 18656 29588
rect 18432 29430 18552 29458
rect 18328 28960 18380 28966
rect 18328 28902 18380 28908
rect 18340 28558 18368 28902
rect 18236 28552 18288 28558
rect 18236 28494 18288 28500
rect 18328 28552 18380 28558
rect 18328 28494 18380 28500
rect 18052 28416 18104 28422
rect 18052 28358 18104 28364
rect 17592 27600 17644 27606
rect 17592 27542 17644 27548
rect 18064 27538 18092 28358
rect 17224 27532 17276 27538
rect 17224 27474 17276 27480
rect 18052 27532 18104 27538
rect 18052 27474 18104 27480
rect 17132 26920 17184 26926
rect 17132 26862 17184 26868
rect 17144 26382 17172 26862
rect 15200 26376 15252 26382
rect 15200 26318 15252 26324
rect 16212 26376 16264 26382
rect 17132 26376 17184 26382
rect 16212 26318 16264 26324
rect 16960 26336 17132 26364
rect 16224 25294 16252 26318
rect 16960 25294 16988 26336
rect 17132 26318 17184 26324
rect 17040 26240 17092 26246
rect 17040 26182 17092 26188
rect 17052 25362 17080 26182
rect 17040 25356 17092 25362
rect 17040 25298 17092 25304
rect 15292 25288 15344 25294
rect 15292 25230 15344 25236
rect 15936 25288 15988 25294
rect 15936 25230 15988 25236
rect 16212 25288 16264 25294
rect 16212 25230 16264 25236
rect 16948 25288 17000 25294
rect 16948 25230 17000 25236
rect 15304 24138 15332 25230
rect 15948 24342 15976 25230
rect 16120 25220 16172 25226
rect 16120 25162 16172 25168
rect 16132 24954 16160 25162
rect 16120 24948 16172 24954
rect 16120 24890 16172 24896
rect 15384 24336 15436 24342
rect 15384 24278 15436 24284
rect 15936 24336 15988 24342
rect 15936 24278 15988 24284
rect 15396 24206 15424 24278
rect 16132 24206 16160 24890
rect 16488 24744 16540 24750
rect 16488 24686 16540 24692
rect 16500 24342 16528 24686
rect 16684 24410 16988 24426
rect 16672 24404 16988 24410
rect 16724 24398 16988 24404
rect 16672 24346 16724 24352
rect 16960 24342 16988 24398
rect 16488 24336 16540 24342
rect 16488 24278 16540 24284
rect 16948 24336 17000 24342
rect 16948 24278 17000 24284
rect 16396 24268 16448 24274
rect 16396 24210 16448 24216
rect 15384 24200 15436 24206
rect 15384 24142 15436 24148
rect 16120 24200 16172 24206
rect 16120 24142 16172 24148
rect 15292 24132 15344 24138
rect 15292 24074 15344 24080
rect 15396 23866 15424 24142
rect 15384 23860 15436 23866
rect 16408 23848 16436 24210
rect 17132 24064 17184 24070
rect 17132 24006 17184 24012
rect 17144 23866 17172 24006
rect 17132 23860 17184 23866
rect 16408 23820 16528 23848
rect 15384 23802 15436 23808
rect 15016 23112 15068 23118
rect 15016 23054 15068 23060
rect 16212 22976 16264 22982
rect 16212 22918 16264 22924
rect 15568 22568 15620 22574
rect 15568 22510 15620 22516
rect 15580 22098 15608 22510
rect 15568 22092 15620 22098
rect 15568 22034 15620 22040
rect 14924 21140 14976 21146
rect 14924 21082 14976 21088
rect 14648 20596 14700 20602
rect 14648 20538 14700 20544
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 15108 20460 15160 20466
rect 15108 20402 15160 20408
rect 15292 20460 15344 20466
rect 15292 20402 15344 20408
rect 14556 20256 14608 20262
rect 14556 20198 14608 20204
rect 14568 19786 14596 20198
rect 14556 19780 14608 19786
rect 14556 19722 14608 19728
rect 14660 19514 14688 20402
rect 15120 19718 15148 20402
rect 15304 20058 15332 20402
rect 16224 20262 16252 22918
rect 16304 22636 16356 22642
rect 16304 22578 16356 22584
rect 16396 22636 16448 22642
rect 16396 22578 16448 22584
rect 16316 20602 16344 22578
rect 16408 21486 16436 22578
rect 16500 22234 16528 23820
rect 17132 23802 17184 23808
rect 17040 22636 17092 22642
rect 17040 22578 17092 22584
rect 16764 22432 16816 22438
rect 16764 22374 16816 22380
rect 16488 22228 16540 22234
rect 16488 22170 16540 22176
rect 16396 21480 16448 21486
rect 16396 21422 16448 21428
rect 16408 20942 16436 21422
rect 16396 20936 16448 20942
rect 16396 20878 16448 20884
rect 16304 20596 16356 20602
rect 16304 20538 16356 20544
rect 15752 20256 15804 20262
rect 15752 20198 15804 20204
rect 16212 20256 16264 20262
rect 16212 20198 16264 20204
rect 15292 20052 15344 20058
rect 15292 19994 15344 20000
rect 15108 19712 15160 19718
rect 15108 19654 15160 19660
rect 14648 19508 14700 19514
rect 14648 19450 14700 19456
rect 14464 19440 14516 19446
rect 14464 19382 14516 19388
rect 13544 19304 13596 19310
rect 13544 19246 13596 19252
rect 13820 19304 13872 19310
rect 13820 19246 13872 19252
rect 13556 18290 13584 19246
rect 13360 18284 13412 18290
rect 13360 18226 13412 18232
rect 13544 18284 13596 18290
rect 13544 18226 13596 18232
rect 13728 18284 13780 18290
rect 13728 18226 13780 18232
rect 13740 17882 13768 18226
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 12900 17672 12952 17678
rect 12900 17614 12952 17620
rect 13268 17536 13320 17542
rect 13268 17478 13320 17484
rect 13280 17338 13308 17478
rect 13268 17332 13320 17338
rect 13268 17274 13320 17280
rect 13280 15502 13308 17274
rect 13740 17270 13768 17818
rect 14476 17678 14504 19382
rect 14924 19304 14976 19310
rect 14924 19246 14976 19252
rect 14740 18216 14792 18222
rect 14740 18158 14792 18164
rect 14752 17678 14780 18158
rect 14464 17672 14516 17678
rect 14464 17614 14516 17620
rect 14740 17672 14792 17678
rect 14740 17614 14792 17620
rect 13728 17264 13780 17270
rect 13728 17206 13780 17212
rect 13740 16658 13768 17206
rect 13728 16652 13780 16658
rect 13728 16594 13780 16600
rect 14648 16108 14700 16114
rect 14648 16050 14700 16056
rect 14832 16108 14884 16114
rect 14832 16050 14884 16056
rect 14280 15700 14332 15706
rect 14280 15642 14332 15648
rect 13268 15496 13320 15502
rect 13268 15438 13320 15444
rect 13280 15026 13308 15438
rect 14292 15162 14320 15642
rect 14660 15570 14688 16050
rect 14844 15706 14872 16050
rect 14832 15700 14884 15706
rect 14832 15642 14884 15648
rect 14648 15564 14700 15570
rect 14648 15506 14700 15512
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 14280 15156 14332 15162
rect 14280 15098 14332 15104
rect 14384 15026 14412 15438
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 14372 15020 14424 15026
rect 14372 14962 14424 14968
rect 14384 14482 14412 14962
rect 14936 14482 14964 19246
rect 15120 19242 15148 19654
rect 15304 19446 15332 19994
rect 15764 19514 15792 20198
rect 16316 19854 16344 20538
rect 16304 19848 16356 19854
rect 16304 19790 16356 19796
rect 15752 19508 15804 19514
rect 15752 19450 15804 19456
rect 15292 19440 15344 19446
rect 15292 19382 15344 19388
rect 15108 19236 15160 19242
rect 15108 19178 15160 19184
rect 15120 18834 15148 19178
rect 15108 18828 15160 18834
rect 15108 18770 15160 18776
rect 15304 18766 15332 19382
rect 16500 19310 16528 22170
rect 16580 21888 16632 21894
rect 16580 21830 16632 21836
rect 16592 21554 16620 21830
rect 16580 21548 16632 21554
rect 16580 21490 16632 21496
rect 16592 20874 16620 21490
rect 16776 20942 16804 22374
rect 17052 21962 17080 22578
rect 16856 21956 16908 21962
rect 16856 21898 16908 21904
rect 17040 21956 17092 21962
rect 17040 21898 17092 21904
rect 16868 21486 16896 21898
rect 16948 21616 17000 21622
rect 16948 21558 17000 21564
rect 16856 21480 16908 21486
rect 16856 21422 16908 21428
rect 16960 20942 16988 21558
rect 17236 21554 17264 27474
rect 17592 27464 17644 27470
rect 17592 27406 17644 27412
rect 17776 27464 17828 27470
rect 17776 27406 17828 27412
rect 17604 27130 17632 27406
rect 17592 27124 17644 27130
rect 17592 27066 17644 27072
rect 17788 26586 17816 27406
rect 18144 26988 18196 26994
rect 18144 26930 18196 26936
rect 17868 26920 17920 26926
rect 17868 26862 17920 26868
rect 17776 26580 17828 26586
rect 17776 26522 17828 26528
rect 17788 26450 17816 26522
rect 17776 26444 17828 26450
rect 17776 26386 17828 26392
rect 17880 26382 17908 26862
rect 18156 26450 18184 26930
rect 18144 26444 18196 26450
rect 18144 26386 18196 26392
rect 17868 26376 17920 26382
rect 17868 26318 17920 26324
rect 17880 25906 17908 26318
rect 17868 25900 17920 25906
rect 17868 25842 17920 25848
rect 18156 25770 18184 26386
rect 18144 25764 18196 25770
rect 18144 25706 18196 25712
rect 17868 25288 17920 25294
rect 17868 25230 17920 25236
rect 17316 25152 17368 25158
rect 17316 25094 17368 25100
rect 17500 25152 17552 25158
rect 17500 25094 17552 25100
rect 17328 24682 17356 25094
rect 17316 24676 17368 24682
rect 17316 24618 17368 24624
rect 17512 24274 17540 25094
rect 17880 24954 17908 25230
rect 18248 25226 18276 28494
rect 18432 28490 18460 29430
rect 18616 28966 18644 29582
rect 18604 28960 18656 28966
rect 18604 28902 18656 28908
rect 18604 28552 18656 28558
rect 18604 28494 18656 28500
rect 18420 28484 18472 28490
rect 18420 28426 18472 28432
rect 18432 28150 18460 28426
rect 18616 28218 18644 28494
rect 18604 28212 18656 28218
rect 18604 28154 18656 28160
rect 18420 28144 18472 28150
rect 18420 28086 18472 28092
rect 18512 25968 18564 25974
rect 18512 25910 18564 25916
rect 18524 25430 18552 25910
rect 18880 25900 18932 25906
rect 18880 25842 18932 25848
rect 18604 25696 18656 25702
rect 18604 25638 18656 25644
rect 18616 25498 18644 25638
rect 18604 25492 18656 25498
rect 18604 25434 18656 25440
rect 18512 25424 18564 25430
rect 18512 25366 18564 25372
rect 18892 25294 18920 25842
rect 18880 25288 18932 25294
rect 18880 25230 18932 25236
rect 18236 25220 18288 25226
rect 18288 25180 18368 25208
rect 18236 25162 18288 25168
rect 18144 25152 18196 25158
rect 18144 25094 18196 25100
rect 17868 24948 17920 24954
rect 17868 24890 17920 24896
rect 17684 24812 17736 24818
rect 17684 24754 17736 24760
rect 17696 24410 17724 24754
rect 17868 24608 17920 24614
rect 17868 24550 17920 24556
rect 17684 24404 17736 24410
rect 17684 24346 17736 24352
rect 17500 24268 17552 24274
rect 17500 24210 17552 24216
rect 17592 24200 17644 24206
rect 17592 24142 17644 24148
rect 17604 22982 17632 24142
rect 17592 22976 17644 22982
rect 17592 22918 17644 22924
rect 17880 22094 17908 24550
rect 18156 22094 18184 25094
rect 18236 22228 18288 22234
rect 18236 22170 18288 22176
rect 17604 22066 17908 22094
rect 18064 22066 18184 22094
rect 17224 21548 17276 21554
rect 17224 21490 17276 21496
rect 17604 21486 17632 22066
rect 17868 22024 17920 22030
rect 17868 21966 17920 21972
rect 17776 21888 17828 21894
rect 17880 21876 17908 21966
rect 17880 21848 18000 21876
rect 17776 21830 17828 21836
rect 17788 21554 17816 21830
rect 17972 21622 18000 21848
rect 17960 21616 18012 21622
rect 17960 21558 18012 21564
rect 18064 21570 18092 22066
rect 18248 21978 18276 22170
rect 18340 22166 18368 25180
rect 19076 24750 19104 39850
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 19248 38820 19300 38826
rect 19248 38762 19300 38768
rect 19260 37874 19288 38762
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 19248 37868 19300 37874
rect 19248 37810 19300 37816
rect 19260 35698 19288 37810
rect 19432 37664 19484 37670
rect 19432 37606 19484 37612
rect 19800 37664 19852 37670
rect 19800 37606 19852 37612
rect 19340 37256 19392 37262
rect 19340 37198 19392 37204
rect 19352 36786 19380 37198
rect 19340 36780 19392 36786
rect 19340 36722 19392 36728
rect 19444 36718 19472 37606
rect 19812 37262 19840 37606
rect 19800 37256 19852 37262
rect 19800 37198 19852 37204
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19524 36780 19576 36786
rect 19524 36722 19576 36728
rect 19432 36712 19484 36718
rect 19432 36654 19484 36660
rect 19536 36378 19564 36722
rect 20352 36644 20404 36650
rect 20352 36586 20404 36592
rect 19524 36372 19576 36378
rect 19524 36314 19576 36320
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19248 35692 19300 35698
rect 19248 35634 19300 35640
rect 19260 34610 19288 35634
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19248 34604 19300 34610
rect 19248 34546 19300 34552
rect 19260 34134 19288 34546
rect 19248 34128 19300 34134
rect 19248 34070 19300 34076
rect 19260 32910 19288 34070
rect 19340 34060 19392 34066
rect 19340 34002 19392 34008
rect 19352 33522 19380 34002
rect 19432 33992 19484 33998
rect 19432 33934 19484 33940
rect 20168 33992 20220 33998
rect 20168 33934 20220 33940
rect 19444 33538 19472 33934
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19444 33522 19748 33538
rect 20180 33522 20208 33934
rect 19340 33516 19392 33522
rect 19444 33516 19760 33522
rect 19444 33510 19708 33516
rect 19340 33458 19392 33464
rect 19708 33458 19760 33464
rect 20168 33516 20220 33522
rect 20168 33458 20220 33464
rect 19248 32904 19300 32910
rect 19248 32846 19300 32852
rect 19260 32434 19288 32846
rect 19248 32428 19300 32434
rect 19248 32370 19300 32376
rect 19352 32366 19380 33458
rect 19720 32842 19748 33458
rect 19708 32836 19760 32842
rect 19708 32778 19760 32784
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19340 32360 19392 32366
rect 19340 32302 19392 32308
rect 19352 32026 19380 32302
rect 20180 32298 20208 33458
rect 20260 32496 20312 32502
rect 20260 32438 20312 32444
rect 20168 32292 20220 32298
rect 20168 32234 20220 32240
rect 19984 32224 20036 32230
rect 19984 32166 20036 32172
rect 19340 32020 19392 32026
rect 19340 31962 19392 31968
rect 19352 31346 19380 31962
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19996 31346 20024 32166
rect 20168 31748 20220 31754
rect 20168 31690 20220 31696
rect 20180 31482 20208 31690
rect 20168 31476 20220 31482
rect 20168 31418 20220 31424
rect 19340 31340 19392 31346
rect 19340 31282 19392 31288
rect 19984 31340 20036 31346
rect 19984 31282 20036 31288
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19248 29708 19300 29714
rect 19248 29650 19300 29656
rect 19260 29186 19288 29650
rect 19984 29504 20036 29510
rect 19984 29446 20036 29452
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19432 29232 19484 29238
rect 19260 29170 19380 29186
rect 19432 29174 19484 29180
rect 19260 29164 19392 29170
rect 19260 29158 19340 29164
rect 19340 29106 19392 29112
rect 19444 28762 19472 29174
rect 19432 28756 19484 28762
rect 19432 28698 19484 28704
rect 19996 28626 20024 29446
rect 20076 29164 20128 29170
rect 20076 29106 20128 29112
rect 19984 28620 20036 28626
rect 19984 28562 20036 28568
rect 19432 28484 19484 28490
rect 19432 28426 19484 28432
rect 19444 27606 19472 28426
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 20088 28218 20116 29106
rect 20272 28506 20300 32438
rect 20364 31278 20392 36586
rect 20444 33516 20496 33522
rect 20444 33458 20496 33464
rect 20456 32774 20484 33458
rect 20444 32768 20496 32774
rect 20444 32710 20496 32716
rect 20456 32230 20484 32710
rect 20444 32224 20496 32230
rect 20444 32166 20496 32172
rect 20456 32026 20484 32166
rect 20444 32020 20496 32026
rect 20444 31962 20496 31968
rect 20352 31272 20404 31278
rect 20352 31214 20404 31220
rect 20444 28756 20496 28762
rect 20444 28698 20496 28704
rect 20272 28478 20392 28506
rect 20260 28416 20312 28422
rect 20260 28358 20312 28364
rect 20076 28212 20128 28218
rect 20076 28154 20128 28160
rect 20272 28082 20300 28358
rect 20260 28076 20312 28082
rect 20260 28018 20312 28024
rect 20364 28014 20392 28478
rect 20456 28082 20484 28698
rect 20444 28076 20496 28082
rect 20444 28018 20496 28024
rect 20352 28008 20404 28014
rect 20352 27950 20404 27956
rect 19432 27600 19484 27606
rect 19432 27542 19484 27548
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19984 26240 20036 26246
rect 19984 26182 20036 26188
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19996 25974 20024 26182
rect 19984 25968 20036 25974
rect 19984 25910 20036 25916
rect 19524 25764 19576 25770
rect 19524 25706 19576 25712
rect 19536 25498 19564 25706
rect 19616 25696 19668 25702
rect 19616 25638 19668 25644
rect 20352 25696 20404 25702
rect 20352 25638 20404 25644
rect 19524 25492 19576 25498
rect 19524 25434 19576 25440
rect 19628 25362 19656 25638
rect 19616 25356 19668 25362
rect 19616 25298 19668 25304
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19616 24812 19668 24818
rect 19616 24754 19668 24760
rect 19064 24744 19116 24750
rect 19064 24686 19116 24692
rect 19340 24608 19392 24614
rect 19340 24550 19392 24556
rect 19352 23730 19380 24550
rect 19628 24410 19656 24754
rect 19984 24744 20036 24750
rect 19984 24686 20036 24692
rect 19616 24404 19668 24410
rect 19616 24346 19668 24352
rect 19800 24200 19852 24206
rect 19800 24142 19852 24148
rect 19812 24070 19840 24142
rect 19800 24064 19852 24070
rect 19800 24006 19852 24012
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19340 23724 19392 23730
rect 19340 23666 19392 23672
rect 19996 23186 20024 24686
rect 20076 24404 20128 24410
rect 20076 24346 20128 24352
rect 20088 24206 20116 24346
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 19984 23180 20036 23186
rect 19984 23122 20036 23128
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 18972 22432 19024 22438
rect 18972 22374 19024 22380
rect 18328 22160 18380 22166
rect 18380 22120 18460 22148
rect 18328 22102 18380 22108
rect 18328 22024 18380 22030
rect 18248 21972 18328 21978
rect 18248 21966 18380 21972
rect 18248 21950 18368 21966
rect 18248 21894 18276 21950
rect 18236 21888 18288 21894
rect 18236 21830 18288 21836
rect 17776 21548 17828 21554
rect 18064 21542 18184 21570
rect 17776 21490 17828 21496
rect 18156 21486 18184 21542
rect 17040 21480 17092 21486
rect 17040 21422 17092 21428
rect 17500 21480 17552 21486
rect 17500 21422 17552 21428
rect 17592 21480 17644 21486
rect 17592 21422 17644 21428
rect 18144 21480 18196 21486
rect 18144 21422 18196 21428
rect 17052 21078 17080 21422
rect 17040 21072 17092 21078
rect 17040 21014 17092 21020
rect 16764 20936 16816 20942
rect 16764 20878 16816 20884
rect 16948 20936 17000 20942
rect 16948 20878 17000 20884
rect 16580 20868 16632 20874
rect 16580 20810 16632 20816
rect 16672 20460 16724 20466
rect 16672 20402 16724 20408
rect 16684 20369 16712 20402
rect 16670 20360 16726 20369
rect 16670 20295 16726 20304
rect 16672 19440 16724 19446
rect 16672 19382 16724 19388
rect 16488 19304 16540 19310
rect 16488 19246 16540 19252
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 16304 18284 16356 18290
rect 16304 18226 16356 18232
rect 16132 17882 16160 18226
rect 16316 17882 16344 18226
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 15936 17876 15988 17882
rect 15936 17818 15988 17824
rect 16120 17876 16172 17882
rect 16120 17818 16172 17824
rect 16304 17876 16356 17882
rect 16304 17818 16356 17824
rect 15108 17672 15160 17678
rect 15108 17614 15160 17620
rect 15120 17338 15148 17614
rect 15200 17604 15252 17610
rect 15200 17546 15252 17552
rect 15108 17332 15160 17338
rect 15108 17274 15160 17280
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 15028 16590 15056 17138
rect 15016 16584 15068 16590
rect 15016 16526 15068 16532
rect 15212 16454 15240 17546
rect 15948 17270 15976 17818
rect 16316 17270 16344 17818
rect 15936 17264 15988 17270
rect 15936 17206 15988 17212
rect 16304 17264 16356 17270
rect 16304 17206 16356 17212
rect 15948 16590 15976 17206
rect 16304 16992 16356 16998
rect 16304 16934 16356 16940
rect 16316 16658 16344 16934
rect 16592 16658 16620 18022
rect 16684 17678 16712 19382
rect 16776 18834 16804 20878
rect 16948 20528 17000 20534
rect 17052 20505 17080 21014
rect 17512 20806 17540 21422
rect 17604 20942 17632 21422
rect 17868 21344 17920 21350
rect 17868 21286 17920 21292
rect 17880 21010 17908 21286
rect 17868 21004 17920 21010
rect 17868 20946 17920 20952
rect 17592 20936 17644 20942
rect 17592 20878 17644 20884
rect 17408 20800 17460 20806
rect 17408 20742 17460 20748
rect 17500 20800 17552 20806
rect 17500 20742 17552 20748
rect 16948 20470 17000 20476
rect 17038 20496 17094 20505
rect 16960 19922 16988 20470
rect 17420 20466 17448 20742
rect 17500 20528 17552 20534
rect 17500 20470 17552 20476
rect 17038 20431 17040 20440
rect 17092 20431 17094 20440
rect 17408 20460 17460 20466
rect 17040 20402 17092 20408
rect 17408 20402 17460 20408
rect 17052 20371 17080 20402
rect 17132 20392 17184 20398
rect 17420 20346 17448 20402
rect 17512 20398 17540 20470
rect 17132 20334 17184 20340
rect 17144 20058 17172 20334
rect 17236 20330 17448 20346
rect 17500 20392 17552 20398
rect 17500 20334 17552 20340
rect 17224 20324 17448 20330
rect 17276 20318 17448 20324
rect 17224 20266 17276 20272
rect 17132 20052 17184 20058
rect 17132 19994 17184 20000
rect 16948 19916 17000 19922
rect 16948 19858 17000 19864
rect 16960 19378 16988 19858
rect 17420 19496 17448 20318
rect 17500 19780 17552 19786
rect 17500 19722 17552 19728
rect 17328 19468 17448 19496
rect 16948 19372 17000 19378
rect 16948 19314 17000 19320
rect 17224 19372 17276 19378
rect 17328 19360 17356 19468
rect 17276 19332 17356 19360
rect 17408 19372 17460 19378
rect 17224 19314 17276 19320
rect 17408 19314 17460 19320
rect 16764 18828 16816 18834
rect 16764 18770 16816 18776
rect 16960 18766 16988 19314
rect 16948 18760 17000 18766
rect 16948 18702 17000 18708
rect 17420 18698 17448 19314
rect 17408 18692 17460 18698
rect 17408 18634 17460 18640
rect 16856 18624 16908 18630
rect 16856 18566 16908 18572
rect 16868 17746 16896 18566
rect 17132 18284 17184 18290
rect 17132 18226 17184 18232
rect 17144 17882 17172 18226
rect 17132 17876 17184 17882
rect 17132 17818 17184 17824
rect 16856 17740 16908 17746
rect 16856 17682 16908 17688
rect 16672 17672 16724 17678
rect 16672 17614 16724 17620
rect 16684 17202 16712 17614
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 16868 17066 16896 17682
rect 16948 17536 17000 17542
rect 16948 17478 17000 17484
rect 16960 17338 16988 17478
rect 16948 17332 17000 17338
rect 16948 17274 17000 17280
rect 17144 17270 17172 17818
rect 17132 17264 17184 17270
rect 17132 17206 17184 17212
rect 16856 17060 16908 17066
rect 16856 17002 16908 17008
rect 17316 16992 17368 16998
rect 17316 16934 17368 16940
rect 17328 16794 17356 16934
rect 17316 16788 17368 16794
rect 17316 16730 17368 16736
rect 16028 16652 16080 16658
rect 16028 16594 16080 16600
rect 16304 16652 16356 16658
rect 16304 16594 16356 16600
rect 16580 16652 16632 16658
rect 16580 16594 16632 16600
rect 15936 16584 15988 16590
rect 15936 16526 15988 16532
rect 15844 16516 15896 16522
rect 15844 16458 15896 16464
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 15212 16182 15240 16390
rect 15200 16176 15252 16182
rect 15200 16118 15252 16124
rect 15856 16046 15884 16458
rect 16040 16114 16068 16594
rect 16316 16250 16344 16594
rect 16304 16244 16356 16250
rect 16304 16186 16356 16192
rect 16028 16108 16080 16114
rect 16028 16050 16080 16056
rect 15844 16040 15896 16046
rect 15844 15982 15896 15988
rect 15856 15502 15884 15982
rect 16948 15904 17000 15910
rect 16948 15846 17000 15852
rect 16960 15570 16988 15846
rect 16948 15564 17000 15570
rect 16948 15506 17000 15512
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 16028 15360 16080 15366
rect 16028 15302 16080 15308
rect 16040 14482 16068 15302
rect 17512 15026 17540 19722
rect 17604 19446 17632 20878
rect 18156 20874 18184 21422
rect 17776 20868 17828 20874
rect 17776 20810 17828 20816
rect 18144 20868 18196 20874
rect 18144 20810 18196 20816
rect 17684 20528 17736 20534
rect 17684 20470 17736 20476
rect 17696 20058 17724 20470
rect 17684 20052 17736 20058
rect 17684 19994 17736 20000
rect 17684 19848 17736 19854
rect 17684 19790 17736 19796
rect 17696 19514 17724 19790
rect 17684 19508 17736 19514
rect 17684 19450 17736 19456
rect 17592 19440 17644 19446
rect 17592 19382 17644 19388
rect 17788 17338 17816 20810
rect 18052 20800 18104 20806
rect 18052 20742 18104 20748
rect 17958 20360 18014 20369
rect 17958 20295 18014 20304
rect 17972 20262 18000 20295
rect 17960 20256 18012 20262
rect 17960 20198 18012 20204
rect 18064 17354 18092 20742
rect 18142 20496 18198 20505
rect 18142 20431 18144 20440
rect 18196 20431 18198 20440
rect 18144 20402 18196 20408
rect 18432 20398 18460 22120
rect 18984 22098 19012 22374
rect 20088 22114 20116 24142
rect 20168 24064 20220 24070
rect 20168 24006 20220 24012
rect 20260 24064 20312 24070
rect 20260 24006 20312 24012
rect 18972 22092 19024 22098
rect 18972 22034 19024 22040
rect 19996 22086 20116 22114
rect 19996 21962 20024 22086
rect 20180 21978 20208 24006
rect 20272 23866 20300 24006
rect 20260 23860 20312 23866
rect 20260 23802 20312 23808
rect 20364 23798 20392 25638
rect 20456 24614 20484 28018
rect 20444 24608 20496 24614
rect 20444 24550 20496 24556
rect 20352 23792 20404 23798
rect 20352 23734 20404 23740
rect 20364 22574 20392 23734
rect 20352 22568 20404 22574
rect 20352 22510 20404 22516
rect 20456 22438 20484 24550
rect 20548 23526 20576 41386
rect 23664 40520 23716 40526
rect 23848 40520 23900 40526
rect 23716 40468 23796 40474
rect 23664 40462 23796 40468
rect 23848 40462 23900 40468
rect 23676 40446 23796 40462
rect 22284 40384 22336 40390
rect 22284 40326 22336 40332
rect 22192 40112 22244 40118
rect 22192 40054 22244 40060
rect 21732 40044 21784 40050
rect 21732 39986 21784 39992
rect 20904 39908 20956 39914
rect 20904 39850 20956 39856
rect 20916 39030 20944 39850
rect 21744 39438 21772 39986
rect 21732 39432 21784 39438
rect 21732 39374 21784 39380
rect 20904 39024 20956 39030
rect 20904 38966 20956 38972
rect 20628 38888 20680 38894
rect 20628 38830 20680 38836
rect 20640 37806 20668 38830
rect 20628 37800 20680 37806
rect 20628 37742 20680 37748
rect 20640 37466 20668 37742
rect 20720 37732 20772 37738
rect 20720 37674 20772 37680
rect 20628 37460 20680 37466
rect 20628 37402 20680 37408
rect 20640 36854 20668 37402
rect 20628 36848 20680 36854
rect 20628 36790 20680 36796
rect 20732 36786 20760 37674
rect 20916 37346 20944 38966
rect 21744 38894 21772 39374
rect 22204 39370 22232 40054
rect 22296 39982 22324 40326
rect 22284 39976 22336 39982
rect 22284 39918 22336 39924
rect 22192 39364 22244 39370
rect 22192 39306 22244 39312
rect 22204 38962 22232 39306
rect 22296 38962 22324 39918
rect 23020 39908 23072 39914
rect 23020 39850 23072 39856
rect 23032 39506 23060 39850
rect 23664 39840 23716 39846
rect 23664 39782 23716 39788
rect 23020 39500 23072 39506
rect 23020 39442 23072 39448
rect 23676 39438 23704 39782
rect 23768 39574 23796 40446
rect 23860 39642 23888 40462
rect 24400 40180 24452 40186
rect 24400 40122 24452 40128
rect 24032 40112 24084 40118
rect 24032 40054 24084 40060
rect 23940 39976 23992 39982
rect 23940 39918 23992 39924
rect 23848 39636 23900 39642
rect 23848 39578 23900 39584
rect 23756 39568 23808 39574
rect 23808 39516 23888 39522
rect 23756 39510 23888 39516
rect 23768 39494 23888 39510
rect 22376 39432 22428 39438
rect 22376 39374 22428 39380
rect 23664 39432 23716 39438
rect 23664 39374 23716 39380
rect 23756 39432 23808 39438
rect 23756 39374 23808 39380
rect 22192 38956 22244 38962
rect 22192 38898 22244 38904
rect 22284 38956 22336 38962
rect 22284 38898 22336 38904
rect 21732 38888 21784 38894
rect 21732 38830 21784 38836
rect 20824 37318 20944 37346
rect 20824 37262 20852 37318
rect 20812 37256 20864 37262
rect 20812 37198 20864 37204
rect 20720 36780 20772 36786
rect 20720 36722 20772 36728
rect 20824 35306 20852 37198
rect 20904 37188 20956 37194
rect 20904 37130 20956 37136
rect 20916 36922 20944 37130
rect 22204 36922 22232 38898
rect 22296 38350 22324 38898
rect 22388 38554 22416 39374
rect 23572 39296 23624 39302
rect 23572 39238 23624 39244
rect 23584 38962 23612 39238
rect 23572 38956 23624 38962
rect 23572 38898 23624 38904
rect 23480 38888 23532 38894
rect 23480 38830 23532 38836
rect 23388 38752 23440 38758
rect 23388 38694 23440 38700
rect 22376 38548 22428 38554
rect 22376 38490 22428 38496
rect 22284 38344 22336 38350
rect 22284 38286 22336 38292
rect 23400 37874 23428 38694
rect 23492 38554 23520 38830
rect 23572 38820 23624 38826
rect 23572 38762 23624 38768
rect 23480 38548 23532 38554
rect 23480 38490 23532 38496
rect 23584 38350 23612 38762
rect 23572 38344 23624 38350
rect 23572 38286 23624 38292
rect 23676 38282 23704 39374
rect 23768 39030 23796 39374
rect 23756 39024 23808 39030
rect 23756 38966 23808 38972
rect 23768 38826 23796 38966
rect 23756 38820 23808 38826
rect 23756 38762 23808 38768
rect 23664 38276 23716 38282
rect 23664 38218 23716 38224
rect 23860 38214 23888 39494
rect 23952 38894 23980 39918
rect 24044 39438 24072 40054
rect 24032 39432 24084 39438
rect 24032 39374 24084 39380
rect 23940 38888 23992 38894
rect 23940 38830 23992 38836
rect 23940 38752 23992 38758
rect 23940 38694 23992 38700
rect 23848 38208 23900 38214
rect 23848 38150 23900 38156
rect 23388 37868 23440 37874
rect 23388 37810 23440 37816
rect 22284 37664 22336 37670
rect 22284 37606 22336 37612
rect 20904 36916 20956 36922
rect 20904 36858 20956 36864
rect 22192 36916 22244 36922
rect 22192 36858 22244 36864
rect 21732 36848 21784 36854
rect 21732 36790 21784 36796
rect 21548 36780 21600 36786
rect 21548 36722 21600 36728
rect 21560 36174 21588 36722
rect 21744 36242 21772 36790
rect 22296 36786 22324 37606
rect 23848 37256 23900 37262
rect 23848 37198 23900 37204
rect 22468 37188 22520 37194
rect 22468 37130 22520 37136
rect 22284 36780 22336 36786
rect 22284 36722 22336 36728
rect 22480 36718 22508 37130
rect 22468 36712 22520 36718
rect 22468 36654 22520 36660
rect 21732 36236 21784 36242
rect 21732 36178 21784 36184
rect 21548 36168 21600 36174
rect 21548 36110 21600 36116
rect 21456 35488 21508 35494
rect 21456 35430 21508 35436
rect 20824 35278 20944 35306
rect 20812 35148 20864 35154
rect 20812 35090 20864 35096
rect 20720 34944 20772 34950
rect 20720 34886 20772 34892
rect 20732 34474 20760 34886
rect 20824 34610 20852 35090
rect 20916 35018 20944 35278
rect 21468 35154 21496 35430
rect 21560 35290 21588 36110
rect 21744 35834 21772 36178
rect 21732 35828 21784 35834
rect 21732 35770 21784 35776
rect 22008 35692 22060 35698
rect 22008 35634 22060 35640
rect 21548 35284 21600 35290
rect 21548 35226 21600 35232
rect 21456 35148 21508 35154
rect 21456 35090 21508 35096
rect 20904 35012 20956 35018
rect 20904 34954 20956 34960
rect 20916 34746 20944 34954
rect 21548 34944 21600 34950
rect 21548 34886 21600 34892
rect 20904 34740 20956 34746
rect 20904 34682 20956 34688
rect 20812 34604 20864 34610
rect 20812 34546 20864 34552
rect 20720 34468 20772 34474
rect 20720 34410 20772 34416
rect 20732 34202 20760 34410
rect 20720 34196 20772 34202
rect 20720 34138 20772 34144
rect 20916 33454 20944 34682
rect 21560 34678 21588 34886
rect 21548 34672 21600 34678
rect 21548 34614 21600 34620
rect 21824 34604 21876 34610
rect 21824 34546 21876 34552
rect 21180 33924 21232 33930
rect 21180 33866 21232 33872
rect 20996 33856 21048 33862
rect 20996 33798 21048 33804
rect 21008 33590 21036 33798
rect 21192 33658 21220 33866
rect 21180 33652 21232 33658
rect 21180 33594 21232 33600
rect 20996 33584 21048 33590
rect 20996 33526 21048 33532
rect 21088 33516 21140 33522
rect 21088 33458 21140 33464
rect 20904 33448 20956 33454
rect 20904 33390 20956 33396
rect 21100 33114 21128 33458
rect 21088 33108 21140 33114
rect 21088 33050 21140 33056
rect 21192 32910 21220 33594
rect 21272 33516 21324 33522
rect 21272 33458 21324 33464
rect 21284 32978 21312 33458
rect 21272 32972 21324 32978
rect 21272 32914 21324 32920
rect 21180 32904 21232 32910
rect 21180 32846 21232 32852
rect 21284 32434 21312 32914
rect 21836 32910 21864 34546
rect 22020 34542 22048 35634
rect 22008 34536 22060 34542
rect 22008 34478 22060 34484
rect 22020 33998 22048 34478
rect 22008 33992 22060 33998
rect 22008 33934 22060 33940
rect 21824 32904 21876 32910
rect 21824 32846 21876 32852
rect 21272 32428 21324 32434
rect 21272 32370 21324 32376
rect 21272 32224 21324 32230
rect 21272 32166 21324 32172
rect 21284 31414 21312 32166
rect 21836 31754 21864 32846
rect 22192 32768 22244 32774
rect 22192 32710 22244 32716
rect 22100 32428 22152 32434
rect 22100 32370 22152 32376
rect 22008 32360 22060 32366
rect 22008 32302 22060 32308
rect 22020 31890 22048 32302
rect 22112 32026 22140 32370
rect 22100 32020 22152 32026
rect 22100 31962 22152 31968
rect 22008 31884 22060 31890
rect 22008 31826 22060 31832
rect 22204 31822 22232 32710
rect 22480 31890 22508 36654
rect 23480 36168 23532 36174
rect 23480 36110 23532 36116
rect 23492 35698 23520 36110
rect 23480 35692 23532 35698
rect 23480 35634 23532 35640
rect 23204 35624 23256 35630
rect 23204 35566 23256 35572
rect 23216 35290 23244 35566
rect 23204 35284 23256 35290
rect 23204 35226 23256 35232
rect 23216 34542 23244 35226
rect 23492 35018 23520 35634
rect 23756 35488 23808 35494
rect 23756 35430 23808 35436
rect 23480 35012 23532 35018
rect 23480 34954 23532 34960
rect 23664 35012 23716 35018
rect 23664 34954 23716 34960
rect 23676 34746 23704 34954
rect 23480 34740 23532 34746
rect 23480 34682 23532 34688
rect 23664 34740 23716 34746
rect 23664 34682 23716 34688
rect 23204 34536 23256 34542
rect 23204 34478 23256 34484
rect 23492 33998 23520 34682
rect 23768 34610 23796 35430
rect 23860 35086 23888 37198
rect 23952 37194 23980 38694
rect 23940 37188 23992 37194
rect 23940 37130 23992 37136
rect 23940 36576 23992 36582
rect 23940 36518 23992 36524
rect 23848 35080 23900 35086
rect 23848 35022 23900 35028
rect 23756 34604 23808 34610
rect 23756 34546 23808 34552
rect 23480 33992 23532 33998
rect 23480 33934 23532 33940
rect 23860 33454 23888 35022
rect 23952 34678 23980 36518
rect 24044 35894 24072 39374
rect 24412 38962 24440 40122
rect 24492 39976 24544 39982
rect 24492 39918 24544 39924
rect 24504 39438 24532 39918
rect 24492 39432 24544 39438
rect 24492 39374 24544 39380
rect 24400 38956 24452 38962
rect 24400 38898 24452 38904
rect 24492 38888 24544 38894
rect 24492 38830 24544 38836
rect 24504 38010 24532 38830
rect 24584 38344 24636 38350
rect 24584 38286 24636 38292
rect 24492 38004 24544 38010
rect 24492 37946 24544 37952
rect 24596 37942 24624 38286
rect 24584 37936 24636 37942
rect 24584 37878 24636 37884
rect 24596 37262 24624 37878
rect 24584 37256 24636 37262
rect 24584 37198 24636 37204
rect 24044 35866 24164 35894
rect 24032 35828 24084 35834
rect 24032 35770 24084 35776
rect 24044 34678 24072 35770
rect 24136 35630 24164 35866
rect 24124 35624 24176 35630
rect 24124 35566 24176 35572
rect 23940 34672 23992 34678
rect 23940 34614 23992 34620
rect 24032 34672 24084 34678
rect 24032 34614 24084 34620
rect 23848 33448 23900 33454
rect 23848 33390 23900 33396
rect 23860 32978 23888 33390
rect 23848 32972 23900 32978
rect 23848 32914 23900 32920
rect 23388 32836 23440 32842
rect 23388 32778 23440 32784
rect 23400 32230 23428 32778
rect 23860 32502 23888 32914
rect 24044 32910 24072 34614
rect 24032 32904 24084 32910
rect 24032 32846 24084 32852
rect 24044 32570 24072 32846
rect 24136 32774 24164 35566
rect 24688 33386 24716 47126
rect 24952 46504 25004 46510
rect 24952 46446 25004 46452
rect 24964 45626 24992 46446
rect 25148 46034 25176 49200
rect 25320 47048 25372 47054
rect 25320 46990 25372 46996
rect 25332 46646 25360 46990
rect 25320 46640 25372 46646
rect 25320 46582 25372 46588
rect 25792 46510 25820 49200
rect 25780 46504 25832 46510
rect 25780 46446 25832 46452
rect 27080 46374 27108 49200
rect 29656 46510 29684 49200
rect 29736 47048 29788 47054
rect 29736 46990 29788 46996
rect 29368 46504 29420 46510
rect 29368 46446 29420 46452
rect 29644 46504 29696 46510
rect 29644 46446 29696 46452
rect 27068 46368 27120 46374
rect 27068 46310 27120 46316
rect 29380 46170 29408 46446
rect 29368 46164 29420 46170
rect 29368 46106 29420 46112
rect 25228 46096 25280 46102
rect 25228 46038 25280 46044
rect 25136 46028 25188 46034
rect 25136 45970 25188 45976
rect 24952 45620 25004 45626
rect 24952 45562 25004 45568
rect 25240 45490 25268 46038
rect 29748 46034 29776 46990
rect 30300 46034 30328 49200
rect 31588 47138 31616 49200
rect 31588 47110 31800 47138
rect 31772 47054 31800 47110
rect 31760 47048 31812 47054
rect 31760 46990 31812 46996
rect 33140 47048 33192 47054
rect 33140 46990 33192 46996
rect 32496 46912 32548 46918
rect 32496 46854 32548 46860
rect 29736 46028 29788 46034
rect 29736 45970 29788 45976
rect 30288 46028 30340 46034
rect 30288 45970 30340 45976
rect 29000 45960 29052 45966
rect 29000 45902 29052 45908
rect 25320 45824 25372 45830
rect 25320 45766 25372 45772
rect 25332 45626 25360 45766
rect 25320 45620 25372 45626
rect 25320 45562 25372 45568
rect 25228 45484 25280 45490
rect 25228 45426 25280 45432
rect 25240 45286 25268 45426
rect 29012 45354 29040 45902
rect 29920 45892 29972 45898
rect 29920 45834 29972 45840
rect 29932 45558 29960 45834
rect 29920 45552 29972 45558
rect 29920 45494 29972 45500
rect 29828 45484 29880 45490
rect 29828 45426 29880 45432
rect 29000 45348 29052 45354
rect 29000 45290 29052 45296
rect 25228 45280 25280 45286
rect 25228 45222 25280 45228
rect 29012 44198 29040 45290
rect 29000 44192 29052 44198
rect 29000 44134 29052 44140
rect 29644 44192 29696 44198
rect 29644 44134 29696 44140
rect 24952 40044 25004 40050
rect 24952 39986 25004 39992
rect 24964 39370 24992 39986
rect 25596 39432 25648 39438
rect 25596 39374 25648 39380
rect 24952 39364 25004 39370
rect 24952 39306 25004 39312
rect 25608 39030 25636 39374
rect 25596 39024 25648 39030
rect 25596 38966 25648 38972
rect 24860 38752 24912 38758
rect 24860 38694 24912 38700
rect 24872 38350 24900 38694
rect 25608 38554 25636 38966
rect 28448 38956 28500 38962
rect 28448 38898 28500 38904
rect 25596 38548 25648 38554
rect 25596 38490 25648 38496
rect 24860 38344 24912 38350
rect 24860 38286 24912 38292
rect 28460 37330 28488 38898
rect 28448 37324 28500 37330
rect 28448 37266 28500 37272
rect 27712 37256 27764 37262
rect 27712 37198 27764 37204
rect 28080 37256 28132 37262
rect 28080 37198 28132 37204
rect 28172 37256 28224 37262
rect 28172 37198 28224 37204
rect 24768 37120 24820 37126
rect 24768 37062 24820 37068
rect 26056 37120 26108 37126
rect 26056 37062 26108 37068
rect 24780 36582 24808 37062
rect 24952 36780 25004 36786
rect 24952 36722 25004 36728
rect 25596 36780 25648 36786
rect 25596 36722 25648 36728
rect 24860 36712 24912 36718
rect 24860 36654 24912 36660
rect 24768 36576 24820 36582
rect 24768 36518 24820 36524
rect 24780 35834 24808 36518
rect 24872 36378 24900 36654
rect 24860 36372 24912 36378
rect 24860 36314 24912 36320
rect 24872 35834 24900 36314
rect 24768 35828 24820 35834
rect 24768 35770 24820 35776
rect 24860 35828 24912 35834
rect 24860 35770 24912 35776
rect 24964 35698 24992 36722
rect 25228 36100 25280 36106
rect 25228 36042 25280 36048
rect 25044 36032 25096 36038
rect 25044 35974 25096 35980
rect 24952 35692 25004 35698
rect 24952 35634 25004 35640
rect 24964 35562 24992 35634
rect 24768 35556 24820 35562
rect 24768 35498 24820 35504
rect 24952 35556 25004 35562
rect 24952 35498 25004 35504
rect 24780 34610 24808 35498
rect 24860 34944 24912 34950
rect 24860 34886 24912 34892
rect 24872 34610 24900 34886
rect 24964 34746 24992 35498
rect 25056 35290 25084 35974
rect 25240 35834 25268 36042
rect 25228 35828 25280 35834
rect 25228 35770 25280 35776
rect 25608 35698 25636 36722
rect 25688 36644 25740 36650
rect 25688 36586 25740 36592
rect 25596 35692 25648 35698
rect 25596 35634 25648 35640
rect 25136 35488 25188 35494
rect 25136 35430 25188 35436
rect 25148 35290 25176 35430
rect 25044 35284 25096 35290
rect 25044 35226 25096 35232
rect 25136 35284 25188 35290
rect 25136 35226 25188 35232
rect 24952 34740 25004 34746
rect 24952 34682 25004 34688
rect 24768 34604 24820 34610
rect 24768 34546 24820 34552
rect 24860 34604 24912 34610
rect 24860 34546 24912 34552
rect 25700 34134 25728 36586
rect 26068 36038 26096 37062
rect 27724 36786 27752 37198
rect 27712 36780 27764 36786
rect 27712 36722 27764 36728
rect 27988 36780 28040 36786
rect 27988 36722 28040 36728
rect 27712 36576 27764 36582
rect 27712 36518 27764 36524
rect 26332 36372 26384 36378
rect 26332 36314 26384 36320
rect 26148 36100 26200 36106
rect 26148 36042 26200 36048
rect 26056 36032 26108 36038
rect 26056 35974 26108 35980
rect 25780 35760 25832 35766
rect 25780 35702 25832 35708
rect 25792 35290 25820 35702
rect 26160 35698 26188 36042
rect 26344 35698 26372 36314
rect 27724 36174 27752 36518
rect 28000 36378 28028 36722
rect 27988 36372 28040 36378
rect 27988 36314 28040 36320
rect 28092 36310 28120 37198
rect 28184 36922 28212 37198
rect 28172 36916 28224 36922
rect 28172 36858 28224 36864
rect 28080 36304 28132 36310
rect 28080 36246 28132 36252
rect 28460 36174 28488 37266
rect 27436 36168 27488 36174
rect 27436 36110 27488 36116
rect 27712 36168 27764 36174
rect 27712 36110 27764 36116
rect 28448 36168 28500 36174
rect 28448 36110 28500 36116
rect 26516 36032 26568 36038
rect 26516 35974 26568 35980
rect 26528 35766 26556 35974
rect 26516 35760 26568 35766
rect 26516 35702 26568 35708
rect 26148 35692 26200 35698
rect 26148 35634 26200 35640
rect 26332 35692 26384 35698
rect 26332 35634 26384 35640
rect 27344 35692 27396 35698
rect 27344 35634 27396 35640
rect 26056 35556 26108 35562
rect 26056 35498 26108 35504
rect 25780 35284 25832 35290
rect 25780 35226 25832 35232
rect 25872 35080 25924 35086
rect 25872 35022 25924 35028
rect 26068 35034 26096 35498
rect 26160 35154 26188 35634
rect 26148 35148 26200 35154
rect 26148 35090 26200 35096
rect 26240 35080 26292 35086
rect 26068 35028 26240 35034
rect 26068 35022 26292 35028
rect 25780 34672 25832 34678
rect 25780 34614 25832 34620
rect 25884 34626 25912 35022
rect 26068 35006 26280 35022
rect 26344 34746 26372 35634
rect 27068 35624 27120 35630
rect 27068 35566 27120 35572
rect 26332 34740 26384 34746
rect 26332 34682 26384 34688
rect 25688 34128 25740 34134
rect 25688 34070 25740 34076
rect 25596 33856 25648 33862
rect 25596 33798 25648 33804
rect 25608 33590 25636 33798
rect 25700 33590 25728 34070
rect 25596 33584 25648 33590
rect 25596 33526 25648 33532
rect 25688 33584 25740 33590
rect 25688 33526 25740 33532
rect 25792 33522 25820 34614
rect 25884 34598 26372 34626
rect 27080 34610 27108 35566
rect 27160 34944 27212 34950
rect 27160 34886 27212 34892
rect 27172 34610 27200 34886
rect 26240 34536 26292 34542
rect 26240 34478 26292 34484
rect 24860 33516 24912 33522
rect 24860 33458 24912 33464
rect 25780 33516 25832 33522
rect 25780 33458 25832 33464
rect 24676 33380 24728 33386
rect 24676 33322 24728 33328
rect 24124 32768 24176 32774
rect 24124 32710 24176 32716
rect 24032 32564 24084 32570
rect 24032 32506 24084 32512
rect 23848 32496 23900 32502
rect 23848 32438 23900 32444
rect 23388 32224 23440 32230
rect 23388 32166 23440 32172
rect 23400 31890 23428 32166
rect 22468 31884 22520 31890
rect 22468 31826 22520 31832
rect 23388 31884 23440 31890
rect 23388 31826 23440 31832
rect 22192 31816 22244 31822
rect 22192 31758 22244 31764
rect 21836 31726 21956 31754
rect 21272 31408 21324 31414
rect 21272 31350 21324 31356
rect 21548 30048 21600 30054
rect 21548 29990 21600 29996
rect 20904 29708 20956 29714
rect 20904 29650 20956 29656
rect 20628 29640 20680 29646
rect 20628 29582 20680 29588
rect 20640 29170 20668 29582
rect 20628 29164 20680 29170
rect 20628 29106 20680 29112
rect 20640 28558 20668 29106
rect 20916 28626 20944 29650
rect 21560 29578 21588 29990
rect 21548 29572 21600 29578
rect 21548 29514 21600 29520
rect 21180 28960 21232 28966
rect 21180 28902 21232 28908
rect 20904 28620 20956 28626
rect 20904 28562 20956 28568
rect 21192 28558 21220 28902
rect 20628 28552 20680 28558
rect 20628 28494 20680 28500
rect 21180 28552 21232 28558
rect 21180 28494 21232 28500
rect 21192 27130 21220 28494
rect 21180 27124 21232 27130
rect 21180 27066 21232 27072
rect 20996 26920 21048 26926
rect 20996 26862 21048 26868
rect 21364 26920 21416 26926
rect 21364 26862 21416 26868
rect 20812 26784 20864 26790
rect 20812 26726 20864 26732
rect 20824 26382 20852 26726
rect 20812 26376 20864 26382
rect 20812 26318 20864 26324
rect 21008 25430 21036 26862
rect 21376 26518 21404 26862
rect 21364 26512 21416 26518
rect 21364 26454 21416 26460
rect 20996 25424 21048 25430
rect 20996 25366 21048 25372
rect 20628 25288 20680 25294
rect 20628 25230 20680 25236
rect 20640 24954 20668 25230
rect 20628 24948 20680 24954
rect 20628 24890 20680 24896
rect 21376 24274 21404 26454
rect 21456 26240 21508 26246
rect 21456 26182 21508 26188
rect 21468 26042 21496 26182
rect 21456 26036 21508 26042
rect 21456 25978 21508 25984
rect 21468 25294 21496 25978
rect 21640 25832 21692 25838
rect 21640 25774 21692 25780
rect 21652 25294 21680 25774
rect 21456 25288 21508 25294
rect 21456 25230 21508 25236
rect 21640 25288 21692 25294
rect 21640 25230 21692 25236
rect 21364 24268 21416 24274
rect 21364 24210 21416 24216
rect 20628 24132 20680 24138
rect 20628 24074 20680 24080
rect 20640 23866 20668 24074
rect 20628 23860 20680 23866
rect 20628 23802 20680 23808
rect 20536 23520 20588 23526
rect 20536 23462 20588 23468
rect 21272 23316 21324 23322
rect 21272 23258 21324 23264
rect 21284 22642 21312 23258
rect 20996 22636 21048 22642
rect 20996 22578 21048 22584
rect 21272 22636 21324 22642
rect 21272 22578 21324 22584
rect 20720 22500 20772 22506
rect 20720 22442 20772 22448
rect 20444 22432 20496 22438
rect 20444 22374 20496 22380
rect 20088 21962 20208 21978
rect 19984 21956 20036 21962
rect 19984 21898 20036 21904
rect 20076 21956 20208 21962
rect 20128 21950 20208 21956
rect 20076 21898 20128 21904
rect 20088 21842 20116 21898
rect 19996 21814 20116 21842
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19340 20800 19392 20806
rect 19340 20742 19392 20748
rect 19352 20466 19380 20742
rect 19340 20460 19392 20466
rect 19340 20402 19392 20408
rect 18420 20392 18472 20398
rect 18420 20334 18472 20340
rect 18432 19334 18460 20334
rect 19444 20058 19472 20878
rect 19996 20806 20024 21814
rect 20456 21350 20484 22374
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 20456 21146 20484 21286
rect 20076 21140 20128 21146
rect 20076 21082 20128 21088
rect 20444 21140 20496 21146
rect 20444 21082 20496 21088
rect 19984 20800 20036 20806
rect 19984 20742 20036 20748
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19432 20052 19484 20058
rect 19432 19994 19484 20000
rect 19996 19854 20024 20742
rect 20088 20312 20116 21082
rect 20444 20936 20496 20942
rect 20444 20878 20496 20884
rect 20260 20324 20312 20330
rect 20088 20284 20260 20312
rect 19984 19848 20036 19854
rect 19984 19790 20036 19796
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 20088 19446 20116 20284
rect 20260 20266 20312 20272
rect 20352 20256 20404 20262
rect 20352 20198 20404 20204
rect 20364 19854 20392 20198
rect 20456 19990 20484 20878
rect 20732 20534 20760 22442
rect 21008 22098 21036 22578
rect 20996 22092 21048 22098
rect 20996 22034 21048 22040
rect 21180 21956 21232 21962
rect 21180 21898 21232 21904
rect 21192 20602 21220 21898
rect 21284 21622 21312 22578
rect 21272 21616 21324 21622
rect 21272 21558 21324 21564
rect 21180 20596 21232 20602
rect 21180 20538 21232 20544
rect 20720 20528 20772 20534
rect 20720 20470 20772 20476
rect 20444 19984 20496 19990
rect 20444 19926 20496 19932
rect 20352 19848 20404 19854
rect 20352 19790 20404 19796
rect 21192 19446 21220 20538
rect 21456 19848 21508 19854
rect 21456 19790 21508 19796
rect 20076 19440 20128 19446
rect 20076 19382 20128 19388
rect 20628 19440 20680 19446
rect 20628 19382 20680 19388
rect 21180 19440 21232 19446
rect 21180 19382 21232 19388
rect 18340 19306 18460 19334
rect 19984 19372 20036 19378
rect 19984 19314 20036 19320
rect 18340 18290 18368 19306
rect 19248 19304 19300 19310
rect 19248 19246 19300 19252
rect 19260 18970 19288 19246
rect 19708 19168 19760 19174
rect 19708 19110 19760 19116
rect 19248 18964 19300 18970
rect 19248 18906 19300 18912
rect 18328 18284 18380 18290
rect 18328 18226 18380 18232
rect 18328 18080 18380 18086
rect 18328 18022 18380 18028
rect 18064 17338 18184 17354
rect 17776 17332 17828 17338
rect 17776 17274 17828 17280
rect 18052 17332 18184 17338
rect 18104 17326 18184 17332
rect 18052 17274 18104 17280
rect 18052 17196 18104 17202
rect 18052 17138 18104 17144
rect 18064 16726 18092 17138
rect 18156 17066 18184 17326
rect 18340 17202 18368 18022
rect 19260 17882 19288 18906
rect 19720 18766 19748 19110
rect 19340 18760 19392 18766
rect 19340 18702 19392 18708
rect 19708 18760 19760 18766
rect 19708 18702 19760 18708
rect 19248 17876 19300 17882
rect 19248 17818 19300 17824
rect 19352 17746 19380 18702
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19996 18426 20024 19314
rect 20640 19242 20668 19382
rect 20628 19236 20680 19242
rect 20628 19178 20680 19184
rect 20536 18624 20588 18630
rect 20536 18566 20588 18572
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 20548 18290 20576 18566
rect 20168 18284 20220 18290
rect 20168 18226 20220 18232
rect 20536 18284 20588 18290
rect 20536 18226 20588 18232
rect 19340 17740 19392 17746
rect 19340 17682 19392 17688
rect 19432 17672 19484 17678
rect 19432 17614 19484 17620
rect 18512 17604 18564 17610
rect 18512 17546 18564 17552
rect 18524 17338 18552 17546
rect 19444 17542 19472 17614
rect 19432 17536 19484 17542
rect 19432 17478 19484 17484
rect 18512 17332 18564 17338
rect 18512 17274 18564 17280
rect 19444 17270 19472 17478
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 20180 17270 20208 18226
rect 20548 18170 20576 18226
rect 20364 18142 20576 18170
rect 20260 17672 20312 17678
rect 20260 17614 20312 17620
rect 20272 17338 20300 17614
rect 20260 17332 20312 17338
rect 20260 17274 20312 17280
rect 19432 17264 19484 17270
rect 19432 17206 19484 17212
rect 20168 17264 20220 17270
rect 20168 17206 20220 17212
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 18144 17060 18196 17066
rect 18144 17002 18196 17008
rect 18052 16720 18104 16726
rect 18052 16662 18104 16668
rect 19444 15570 19472 17206
rect 20260 16516 20312 16522
rect 20260 16458 20312 16464
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19432 15564 19484 15570
rect 19432 15506 19484 15512
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 18236 15496 18288 15502
rect 18236 15438 18288 15444
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 17880 15094 17908 15302
rect 17868 15088 17920 15094
rect 17868 15030 17920 15036
rect 17500 15020 17552 15026
rect 17500 14962 17552 14968
rect 18064 14618 18092 15438
rect 18052 14612 18104 14618
rect 18052 14554 18104 14560
rect 14372 14476 14424 14482
rect 14372 14418 14424 14424
rect 14924 14476 14976 14482
rect 14924 14418 14976 14424
rect 16028 14476 16080 14482
rect 16028 14418 16080 14424
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13464 13938 13492 14214
rect 14384 14074 14412 14418
rect 17500 14408 17552 14414
rect 17500 14350 17552 14356
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 16212 14000 16264 14006
rect 16212 13942 16264 13948
rect 13452 13932 13504 13938
rect 13452 13874 13504 13880
rect 16224 13326 16252 13942
rect 16212 13320 16264 13326
rect 16212 13262 16264 13268
rect 16224 12434 16252 13262
rect 17040 13252 17092 13258
rect 17040 13194 17092 13200
rect 17052 12986 17080 13194
rect 17040 12980 17092 12986
rect 17040 12922 17092 12928
rect 17512 12442 17540 14350
rect 18052 13184 18104 13190
rect 18052 13126 18104 13132
rect 18064 12850 18092 13126
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 18248 12714 18276 15438
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 18788 14816 18840 14822
rect 18788 14758 18840 14764
rect 18800 14414 18828 14758
rect 18328 14408 18380 14414
rect 18328 14350 18380 14356
rect 18512 14408 18564 14414
rect 18512 14350 18564 14356
rect 18788 14408 18840 14414
rect 18788 14350 18840 14356
rect 18340 13394 18368 14350
rect 18328 13388 18380 13394
rect 18328 13330 18380 13336
rect 18524 13326 18552 14350
rect 19444 14074 19472 14962
rect 19984 14408 20036 14414
rect 19984 14350 20036 14356
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 18512 13320 18564 13326
rect 18512 13262 18564 13268
rect 18328 13252 18380 13258
rect 18328 13194 18380 13200
rect 18236 12708 18288 12714
rect 18236 12650 18288 12656
rect 17960 12640 18012 12646
rect 17960 12582 18012 12588
rect 17500 12436 17552 12442
rect 16224 12406 16344 12434
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16224 11082 16252 11494
rect 16316 11082 16344 12406
rect 17500 12378 17552 12384
rect 17972 12238 18000 12582
rect 18248 12434 18276 12650
rect 18156 12406 18276 12434
rect 17960 12232 18012 12238
rect 17960 12174 18012 12180
rect 17040 12096 17092 12102
rect 17040 12038 17092 12044
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 17052 11762 17080 12038
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 17328 11354 17356 12038
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 18156 11286 18184 12406
rect 18340 12238 18368 13194
rect 18328 12232 18380 12238
rect 18328 12174 18380 12180
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 18248 11626 18276 12038
rect 18236 11620 18288 11626
rect 18236 11562 18288 11568
rect 18144 11280 18196 11286
rect 18144 11222 18196 11228
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17960 11144 18012 11150
rect 17960 11086 18012 11092
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 16212 11076 16264 11082
rect 16212 11018 16264 11024
rect 16304 11076 16356 11082
rect 16304 11018 16356 11024
rect 17328 10674 17356 11086
rect 17776 11008 17828 11014
rect 17776 10950 17828 10956
rect 17788 10742 17816 10950
rect 17776 10736 17828 10742
rect 17776 10678 17828 10684
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17972 10266 18000 11086
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 13188 3670 13216 4082
rect 13360 3936 13412 3942
rect 13360 3878 13412 3884
rect 13176 3664 13228 3670
rect 13176 3606 13228 3612
rect 13176 3528 13228 3534
rect 13176 3470 13228 3476
rect 13188 3058 13216 3470
rect 13372 3126 13400 3878
rect 17604 3670 17632 5646
rect 18248 4690 18276 11086
rect 18524 10062 18552 13262
rect 18972 12096 19024 12102
rect 18972 12038 19024 12044
rect 18984 11830 19012 12038
rect 18972 11824 19024 11830
rect 18972 11766 19024 11772
rect 19352 10810 19380 13806
rect 19444 11898 19472 14010
rect 19892 14000 19944 14006
rect 19892 13942 19944 13948
rect 19904 13326 19932 13942
rect 19996 13938 20024 14350
rect 20088 14346 20116 16390
rect 20272 16250 20300 16458
rect 20260 16244 20312 16250
rect 20260 16186 20312 16192
rect 20260 15360 20312 15366
rect 20260 15302 20312 15308
rect 20168 15020 20220 15026
rect 20168 14962 20220 14968
rect 20180 14618 20208 14962
rect 20168 14612 20220 14618
rect 20168 14554 20220 14560
rect 20076 14340 20128 14346
rect 20076 14282 20128 14288
rect 20088 14074 20116 14282
rect 20076 14068 20128 14074
rect 20076 14010 20128 14016
rect 19984 13932 20036 13938
rect 19984 13874 20036 13880
rect 19996 13546 20024 13874
rect 19996 13518 20116 13546
rect 19984 13456 20036 13462
rect 19984 13398 20036 13404
rect 19892 13320 19944 13326
rect 19892 13262 19944 13268
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19996 12306 20024 13398
rect 20088 13326 20116 13518
rect 20272 13326 20300 15302
rect 20364 14278 20392 18142
rect 20444 17672 20496 17678
rect 20444 17614 20496 17620
rect 20456 17218 20484 17614
rect 20640 17218 20668 19178
rect 21468 18630 21496 19790
rect 21456 18624 21508 18630
rect 21456 18566 21508 18572
rect 21468 18358 21496 18566
rect 21456 18352 21508 18358
rect 21456 18294 21508 18300
rect 21272 18216 21324 18222
rect 21272 18158 21324 18164
rect 21088 17876 21140 17882
rect 21088 17818 21140 17824
rect 20456 17190 20668 17218
rect 20536 17060 20588 17066
rect 20536 17002 20588 17008
rect 20444 16448 20496 16454
rect 20444 16390 20496 16396
rect 20456 16114 20484 16390
rect 20548 16250 20576 17002
rect 20640 16794 20668 17190
rect 20996 16992 21048 16998
rect 20996 16934 21048 16940
rect 20628 16788 20680 16794
rect 20628 16730 20680 16736
rect 20536 16244 20588 16250
rect 20536 16186 20588 16192
rect 20444 16108 20496 16114
rect 20444 16050 20496 16056
rect 20444 15496 20496 15502
rect 20444 15438 20496 15444
rect 20456 15162 20484 15438
rect 20444 15156 20496 15162
rect 20444 15098 20496 15104
rect 20444 14544 20496 14550
rect 20444 14486 20496 14492
rect 20352 14272 20404 14278
rect 20352 14214 20404 14220
rect 20076 13320 20128 13326
rect 20076 13262 20128 13268
rect 20260 13320 20312 13326
rect 20260 13262 20312 13268
rect 20272 12866 20300 13262
rect 20272 12838 20392 12866
rect 20456 12850 20484 14486
rect 20640 14006 20668 16730
rect 20812 15904 20864 15910
rect 20812 15846 20864 15852
rect 20824 15502 20852 15846
rect 21008 15570 21036 16934
rect 20996 15564 21048 15570
rect 20996 15506 21048 15512
rect 20812 15496 20864 15502
rect 20812 15438 20864 15444
rect 20824 15026 20852 15438
rect 20812 15020 20864 15026
rect 20812 14962 20864 14968
rect 21008 14822 21036 15506
rect 20996 14816 21048 14822
rect 20996 14758 21048 14764
rect 21100 14618 21128 17818
rect 21284 17338 21312 18158
rect 21640 18148 21692 18154
rect 21640 18090 21692 18096
rect 21272 17332 21324 17338
rect 21272 17274 21324 17280
rect 21284 17202 21312 17274
rect 21272 17196 21324 17202
rect 21272 17138 21324 17144
rect 21548 17196 21600 17202
rect 21548 17138 21600 17144
rect 21560 16522 21588 17138
rect 21652 16590 21680 18090
rect 21732 17536 21784 17542
rect 21732 17478 21784 17484
rect 21744 17202 21772 17478
rect 21732 17196 21784 17202
rect 21732 17138 21784 17144
rect 21640 16584 21692 16590
rect 21640 16526 21692 16532
rect 21548 16516 21600 16522
rect 21548 16458 21600 16464
rect 21456 16108 21508 16114
rect 21456 16050 21508 16056
rect 21468 15706 21496 16050
rect 21456 15700 21508 15706
rect 21456 15642 21508 15648
rect 21456 15496 21508 15502
rect 21456 15438 21508 15444
rect 21468 15162 21496 15438
rect 21456 15156 21508 15162
rect 21456 15098 21508 15104
rect 21088 14612 21140 14618
rect 21088 14554 21140 14560
rect 21100 14498 21128 14554
rect 21100 14470 21220 14498
rect 21088 14408 21140 14414
rect 21088 14350 21140 14356
rect 20904 14272 20956 14278
rect 20904 14214 20956 14220
rect 20628 14000 20680 14006
rect 20628 13942 20680 13948
rect 20916 13938 20944 14214
rect 20904 13932 20956 13938
rect 20904 13874 20956 13880
rect 21100 13530 21128 14350
rect 21192 14074 21220 14470
rect 21364 14408 21416 14414
rect 21364 14350 21416 14356
rect 21180 14068 21232 14074
rect 21180 14010 21232 14016
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 21180 13320 21232 13326
rect 21180 13262 21232 13268
rect 21192 12850 21220 13262
rect 21376 12918 21404 14350
rect 21640 13728 21692 13734
rect 21640 13670 21692 13676
rect 21652 13326 21680 13670
rect 21640 13320 21692 13326
rect 21640 13262 21692 13268
rect 21652 12986 21680 13262
rect 21640 12980 21692 12986
rect 21640 12922 21692 12928
rect 21364 12912 21416 12918
rect 21364 12854 21416 12860
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 20272 12374 20300 12718
rect 20260 12368 20312 12374
rect 20260 12310 20312 12316
rect 19984 12300 20036 12306
rect 19984 12242 20036 12248
rect 19984 12164 20036 12170
rect 19984 12106 20036 12112
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 19996 11762 20024 12106
rect 20364 11898 20392 12838
rect 20444 12844 20496 12850
rect 20444 12786 20496 12792
rect 21180 12844 21232 12850
rect 21180 12786 21232 12792
rect 20536 12436 20588 12442
rect 20536 12378 20588 12384
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 19984 11756 20036 11762
rect 19984 11698 20036 11704
rect 19984 11144 20036 11150
rect 19984 11086 20036 11092
rect 19432 11008 19484 11014
rect 19432 10950 19484 10956
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 19444 10742 19472 10950
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19432 10736 19484 10742
rect 19432 10678 19484 10684
rect 18880 10464 18932 10470
rect 18880 10406 18932 10412
rect 18892 10062 18920 10406
rect 19996 10266 20024 11086
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 20548 10130 20576 12378
rect 20812 12096 20864 12102
rect 20812 12038 20864 12044
rect 20720 10668 20772 10674
rect 20720 10610 20772 10616
rect 20732 10470 20760 10610
rect 20720 10464 20772 10470
rect 20720 10406 20772 10412
rect 20732 10266 20760 10406
rect 20720 10260 20772 10266
rect 20720 10202 20772 10208
rect 20536 10124 20588 10130
rect 20536 10066 20588 10072
rect 20732 10062 20760 10202
rect 18420 10056 18472 10062
rect 18420 9998 18472 10004
rect 18512 10056 18564 10062
rect 18512 9998 18564 10004
rect 18880 10056 18932 10062
rect 18880 9998 18932 10004
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 18432 9722 18460 9998
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 18420 9716 18472 9722
rect 18420 9658 18472 9664
rect 20732 9654 20760 9998
rect 20824 9994 20852 12038
rect 21928 11830 21956 31726
rect 22376 31748 22428 31754
rect 22376 31690 22428 31696
rect 22100 30252 22152 30258
rect 22100 30194 22152 30200
rect 22008 30184 22060 30190
rect 22008 30126 22060 30132
rect 22020 29646 22048 30126
rect 22008 29640 22060 29646
rect 22008 29582 22060 29588
rect 22020 28014 22048 29582
rect 22112 29170 22140 30194
rect 22388 30172 22416 31690
rect 22480 31210 22508 31826
rect 23940 31816 23992 31822
rect 23940 31758 23992 31764
rect 22468 31204 22520 31210
rect 22468 31146 22520 31152
rect 23572 30592 23624 30598
rect 23572 30534 23624 30540
rect 23296 30252 23348 30258
rect 23296 30194 23348 30200
rect 22468 30184 22520 30190
rect 22388 30144 22468 30172
rect 22468 30126 22520 30132
rect 22376 30048 22428 30054
rect 22376 29990 22428 29996
rect 22100 29164 22152 29170
rect 22100 29106 22152 29112
rect 22388 28762 22416 29990
rect 22480 29714 22508 30126
rect 23308 29782 23336 30194
rect 23296 29776 23348 29782
rect 23296 29718 23348 29724
rect 22468 29708 22520 29714
rect 22468 29650 22520 29656
rect 23480 29640 23532 29646
rect 23480 29582 23532 29588
rect 22560 29164 22612 29170
rect 22560 29106 22612 29112
rect 22376 28756 22428 28762
rect 22376 28698 22428 28704
rect 22572 28626 22600 29106
rect 22928 29096 22980 29102
rect 22928 29038 22980 29044
rect 22560 28620 22612 28626
rect 22560 28562 22612 28568
rect 22376 28552 22428 28558
rect 22376 28494 22428 28500
rect 22284 28416 22336 28422
rect 22284 28358 22336 28364
rect 22296 28082 22324 28358
rect 22284 28076 22336 28082
rect 22284 28018 22336 28024
rect 22008 28008 22060 28014
rect 22008 27950 22060 27956
rect 22020 27538 22048 27950
rect 22388 27674 22416 28494
rect 22376 27668 22428 27674
rect 22376 27610 22428 27616
rect 22572 27606 22600 28562
rect 22652 28552 22704 28558
rect 22652 28494 22704 28500
rect 22664 28150 22692 28494
rect 22652 28144 22704 28150
rect 22652 28086 22704 28092
rect 22560 27600 22612 27606
rect 22560 27542 22612 27548
rect 22008 27532 22060 27538
rect 22008 27474 22060 27480
rect 22020 26042 22048 27474
rect 22940 27470 22968 29038
rect 23492 28762 23520 29582
rect 23584 29510 23612 30534
rect 23572 29504 23624 29510
rect 23572 29446 23624 29452
rect 23848 29504 23900 29510
rect 23848 29446 23900 29452
rect 23584 29170 23612 29446
rect 23572 29164 23624 29170
rect 23572 29106 23624 29112
rect 23756 29028 23808 29034
rect 23756 28970 23808 28976
rect 23480 28756 23532 28762
rect 23480 28698 23532 28704
rect 23768 28626 23796 28970
rect 23756 28620 23808 28626
rect 23756 28562 23808 28568
rect 23572 28552 23624 28558
rect 23572 28494 23624 28500
rect 23388 28416 23440 28422
rect 23388 28358 23440 28364
rect 23400 28218 23428 28358
rect 23388 28212 23440 28218
rect 23388 28154 23440 28160
rect 23020 27600 23072 27606
rect 23020 27542 23072 27548
rect 23032 27470 23060 27542
rect 23400 27470 23428 28154
rect 22928 27464 22980 27470
rect 22928 27406 22980 27412
rect 23020 27464 23072 27470
rect 23020 27406 23072 27412
rect 23388 27464 23440 27470
rect 23388 27406 23440 27412
rect 22376 26444 22428 26450
rect 22376 26386 22428 26392
rect 22008 26036 22060 26042
rect 22008 25978 22060 25984
rect 22008 24608 22060 24614
rect 22008 24550 22060 24556
rect 22020 24274 22048 24550
rect 22008 24268 22060 24274
rect 22008 24210 22060 24216
rect 22388 23186 22416 26386
rect 22836 24268 22888 24274
rect 22836 24210 22888 24216
rect 22376 23180 22428 23186
rect 22376 23122 22428 23128
rect 22008 22568 22060 22574
rect 22008 22510 22060 22516
rect 22020 22098 22048 22510
rect 22008 22092 22060 22098
rect 22388 22094 22416 23122
rect 22652 22976 22704 22982
rect 22652 22918 22704 22924
rect 22744 22976 22796 22982
rect 22744 22918 22796 22924
rect 22560 22636 22612 22642
rect 22560 22578 22612 22584
rect 22572 22234 22600 22578
rect 22664 22234 22692 22918
rect 22560 22228 22612 22234
rect 22560 22170 22612 22176
rect 22652 22228 22704 22234
rect 22652 22170 22704 22176
rect 22008 22034 22060 22040
rect 22296 22066 22416 22094
rect 22296 21894 22324 22066
rect 22756 22030 22784 22918
rect 22744 22024 22796 22030
rect 22744 21966 22796 21972
rect 22284 21888 22336 21894
rect 22284 21830 22336 21836
rect 22376 21888 22428 21894
rect 22376 21830 22428 21836
rect 22388 21690 22416 21830
rect 22376 21684 22428 21690
rect 22376 21626 22428 21632
rect 22388 20942 22416 21626
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 22008 20868 22060 20874
rect 22008 20810 22060 20816
rect 22020 19854 22048 20810
rect 22376 20256 22428 20262
rect 22376 20198 22428 20204
rect 22008 19848 22060 19854
rect 22008 19790 22060 19796
rect 22100 19848 22152 19854
rect 22100 19790 22152 19796
rect 22112 19281 22140 19790
rect 22192 19712 22244 19718
rect 22192 19654 22244 19660
rect 22204 19378 22232 19654
rect 22388 19378 22416 20198
rect 22192 19372 22244 19378
rect 22192 19314 22244 19320
rect 22376 19372 22428 19378
rect 22848 19360 22876 24210
rect 22940 20806 22968 27406
rect 23032 24410 23060 27406
rect 23584 26790 23612 28494
rect 23756 27396 23808 27402
rect 23756 27338 23808 27344
rect 23572 26784 23624 26790
rect 23572 26726 23624 26732
rect 23584 26586 23612 26726
rect 23768 26586 23796 27338
rect 23572 26580 23624 26586
rect 23572 26522 23624 26528
rect 23756 26580 23808 26586
rect 23756 26522 23808 26528
rect 23388 26240 23440 26246
rect 23388 26182 23440 26188
rect 23400 25974 23428 26182
rect 23388 25968 23440 25974
rect 23388 25910 23440 25916
rect 23860 25362 23888 29446
rect 23952 27962 23980 31758
rect 24768 31340 24820 31346
rect 24768 31282 24820 31288
rect 24780 30054 24808 31282
rect 24872 30122 24900 33458
rect 25688 33448 25740 33454
rect 25688 33390 25740 33396
rect 25228 33312 25280 33318
rect 25228 33254 25280 33260
rect 25240 32910 25268 33254
rect 25228 32904 25280 32910
rect 25228 32846 25280 32852
rect 25228 32768 25280 32774
rect 25228 32710 25280 32716
rect 25044 32428 25096 32434
rect 25044 32370 25096 32376
rect 25056 31822 25084 32370
rect 25044 31816 25096 31822
rect 25044 31758 25096 31764
rect 25136 31680 25188 31686
rect 25136 31622 25188 31628
rect 24952 31476 25004 31482
rect 24952 31418 25004 31424
rect 24860 30116 24912 30122
rect 24860 30058 24912 30064
rect 24768 30048 24820 30054
rect 24768 29990 24820 29996
rect 24780 29646 24808 29990
rect 24964 29866 24992 31418
rect 25148 30666 25176 31622
rect 25240 31210 25268 32710
rect 25700 31686 25728 33390
rect 26252 32570 26280 34478
rect 26344 33454 26372 34598
rect 27068 34604 27120 34610
rect 27068 34546 27120 34552
rect 27160 34604 27212 34610
rect 27160 34546 27212 34552
rect 26608 34060 26660 34066
rect 26608 34002 26660 34008
rect 26620 33522 26648 34002
rect 27172 33998 27200 34546
rect 27252 34400 27304 34406
rect 27252 34342 27304 34348
rect 27264 34202 27292 34342
rect 27252 34196 27304 34202
rect 27252 34138 27304 34144
rect 27264 34066 27292 34138
rect 27252 34060 27304 34066
rect 27252 34002 27304 34008
rect 27160 33992 27212 33998
rect 27160 33934 27212 33940
rect 27172 33658 27200 33934
rect 27160 33652 27212 33658
rect 27160 33594 27212 33600
rect 26608 33516 26660 33522
rect 26608 33458 26660 33464
rect 26332 33448 26384 33454
rect 26332 33390 26384 33396
rect 26344 33114 26372 33390
rect 27172 33114 27200 33594
rect 27252 33516 27304 33522
rect 27356 33504 27384 35634
rect 27448 35290 27476 36110
rect 27724 35494 27752 36110
rect 27804 36032 27856 36038
rect 27804 35974 27856 35980
rect 27712 35488 27764 35494
rect 27712 35430 27764 35436
rect 27436 35284 27488 35290
rect 27436 35226 27488 35232
rect 27620 35148 27672 35154
rect 27620 35090 27672 35096
rect 27528 35080 27580 35086
rect 27528 35022 27580 35028
rect 27540 34610 27568 35022
rect 27528 34604 27580 34610
rect 27528 34546 27580 34552
rect 27632 34202 27660 35090
rect 27620 34196 27672 34202
rect 27620 34138 27672 34144
rect 27816 34134 27844 35974
rect 28724 35828 28776 35834
rect 28724 35770 28776 35776
rect 28632 35488 28684 35494
rect 28632 35430 28684 35436
rect 28644 35154 28672 35430
rect 28632 35148 28684 35154
rect 28632 35090 28684 35096
rect 28736 35086 28764 35770
rect 28724 35080 28776 35086
rect 28724 35022 28776 35028
rect 27804 34128 27856 34134
rect 27804 34070 27856 34076
rect 27436 33992 27488 33998
rect 27436 33934 27488 33940
rect 27448 33658 27476 33934
rect 27436 33652 27488 33658
rect 27436 33594 27488 33600
rect 27304 33476 27384 33504
rect 27252 33458 27304 33464
rect 26332 33108 26384 33114
rect 26332 33050 26384 33056
rect 27160 33108 27212 33114
rect 27160 33050 27212 33056
rect 27448 32978 27476 33594
rect 28736 33590 28764 35022
rect 29368 35012 29420 35018
rect 29368 34954 29420 34960
rect 29380 34746 29408 34954
rect 29368 34740 29420 34746
rect 29368 34682 29420 34688
rect 28724 33584 28776 33590
rect 28724 33526 28776 33532
rect 27528 33312 27580 33318
rect 27528 33254 27580 33260
rect 27436 32972 27488 32978
rect 27436 32914 27488 32920
rect 27540 32910 27568 33254
rect 28356 32972 28408 32978
rect 28356 32914 28408 32920
rect 27528 32904 27580 32910
rect 27528 32846 27580 32852
rect 26240 32564 26292 32570
rect 26240 32506 26292 32512
rect 28368 32502 28396 32914
rect 28736 32570 28764 33526
rect 29092 33380 29144 33386
rect 29092 33322 29144 33328
rect 28724 32564 28776 32570
rect 28724 32506 28776 32512
rect 28356 32496 28408 32502
rect 28356 32438 28408 32444
rect 26148 32428 26200 32434
rect 26148 32370 26200 32376
rect 26516 32428 26568 32434
rect 26516 32370 26568 32376
rect 25872 32360 25924 32366
rect 25872 32302 25924 32308
rect 25780 31816 25832 31822
rect 25780 31758 25832 31764
rect 25688 31680 25740 31686
rect 25688 31622 25740 31628
rect 25792 31482 25820 31758
rect 25884 31754 25912 32302
rect 25884 31726 26004 31754
rect 25872 31680 25924 31686
rect 25976 31657 26004 31726
rect 25872 31622 25924 31628
rect 25962 31648 26018 31657
rect 25780 31476 25832 31482
rect 25780 31418 25832 31424
rect 25884 31346 25912 31622
rect 25962 31583 26018 31592
rect 25596 31340 25648 31346
rect 25596 31282 25648 31288
rect 25688 31340 25740 31346
rect 25688 31282 25740 31288
rect 25872 31340 25924 31346
rect 25872 31282 25924 31288
rect 25504 31272 25556 31278
rect 25504 31214 25556 31220
rect 25228 31204 25280 31210
rect 25228 31146 25280 31152
rect 25412 31136 25464 31142
rect 25412 31078 25464 31084
rect 25424 30734 25452 31078
rect 25412 30728 25464 30734
rect 25412 30670 25464 30676
rect 25136 30660 25188 30666
rect 25136 30602 25188 30608
rect 24872 29838 24992 29866
rect 24768 29640 24820 29646
rect 24768 29582 24820 29588
rect 24780 29170 24808 29582
rect 24768 29164 24820 29170
rect 24768 29106 24820 29112
rect 24872 29102 24900 29838
rect 24952 29708 25004 29714
rect 24952 29650 25004 29656
rect 24964 29594 24992 29650
rect 24964 29566 25084 29594
rect 25056 29510 25084 29566
rect 25044 29504 25096 29510
rect 25044 29446 25096 29452
rect 25148 29322 25176 30602
rect 25412 30048 25464 30054
rect 25412 29990 25464 29996
rect 25424 29714 25452 29990
rect 25516 29782 25544 31214
rect 25504 29776 25556 29782
rect 25504 29718 25556 29724
rect 25412 29708 25464 29714
rect 25412 29650 25464 29656
rect 25056 29294 25176 29322
rect 24400 29096 24452 29102
rect 24400 29038 24452 29044
rect 24860 29096 24912 29102
rect 24860 29038 24912 29044
rect 24412 28762 24440 29038
rect 24400 28756 24452 28762
rect 24400 28698 24452 28704
rect 24872 28558 24900 29038
rect 24124 28552 24176 28558
rect 24124 28494 24176 28500
rect 24860 28552 24912 28558
rect 24860 28494 24912 28500
rect 23952 27934 24072 27962
rect 23940 27872 23992 27878
rect 23940 27814 23992 27820
rect 23952 26382 23980 27814
rect 24044 26518 24072 27934
rect 24032 26512 24084 26518
rect 24032 26454 24084 26460
rect 23940 26376 23992 26382
rect 24136 26330 24164 28494
rect 25056 28082 25084 29294
rect 25516 29170 25544 29718
rect 25504 29164 25556 29170
rect 25504 29106 25556 29112
rect 25608 29034 25636 31282
rect 25596 29028 25648 29034
rect 25596 28970 25648 28976
rect 25044 28076 25096 28082
rect 25044 28018 25096 28024
rect 25412 28076 25464 28082
rect 25412 28018 25464 28024
rect 24676 26988 24728 26994
rect 24676 26930 24728 26936
rect 23940 26318 23992 26324
rect 24044 26302 24164 26330
rect 24688 26314 24716 26930
rect 24860 26784 24912 26790
rect 24860 26726 24912 26732
rect 24676 26308 24728 26314
rect 23848 25356 23900 25362
rect 23848 25298 23900 25304
rect 23664 25288 23716 25294
rect 23664 25230 23716 25236
rect 23480 24812 23532 24818
rect 23480 24754 23532 24760
rect 23572 24812 23624 24818
rect 23572 24754 23624 24760
rect 23112 24744 23164 24750
rect 23112 24686 23164 24692
rect 23020 24404 23072 24410
rect 23020 24346 23072 24352
rect 23124 23866 23152 24686
rect 23112 23860 23164 23866
rect 23112 23802 23164 23808
rect 23204 23724 23256 23730
rect 23204 23666 23256 23672
rect 23216 23186 23244 23666
rect 23492 23594 23520 24754
rect 23584 23866 23612 24754
rect 23676 23866 23704 25230
rect 23756 25152 23808 25158
rect 23756 25094 23808 25100
rect 23572 23860 23624 23866
rect 23572 23802 23624 23808
rect 23664 23860 23716 23866
rect 23664 23802 23716 23808
rect 23480 23588 23532 23594
rect 23480 23530 23532 23536
rect 23204 23180 23256 23186
rect 23204 23122 23256 23128
rect 23216 22778 23244 23122
rect 23204 22772 23256 22778
rect 23204 22714 23256 22720
rect 23572 22092 23624 22098
rect 23768 22094 23796 25094
rect 23860 24750 23888 25298
rect 23848 24744 23900 24750
rect 23848 24686 23900 24692
rect 23848 22160 23900 22166
rect 23848 22102 23900 22108
rect 23572 22034 23624 22040
rect 23676 22066 23796 22094
rect 23584 21706 23612 22034
rect 23676 21894 23704 22066
rect 23664 21888 23716 21894
rect 23664 21830 23716 21836
rect 23112 21684 23164 21690
rect 23584 21678 23704 21706
rect 23112 21626 23164 21632
rect 23124 21078 23152 21626
rect 23676 21554 23704 21678
rect 23664 21548 23716 21554
rect 23664 21490 23716 21496
rect 23112 21072 23164 21078
rect 23480 21072 23532 21078
rect 23112 21014 23164 21020
rect 23308 21020 23480 21026
rect 23308 21014 23532 21020
rect 23308 20998 23520 21014
rect 23308 20942 23336 20998
rect 23296 20936 23348 20942
rect 23296 20878 23348 20884
rect 22928 20800 22980 20806
rect 22928 20742 22980 20748
rect 22848 19332 22968 19360
rect 22376 19314 22428 19320
rect 22098 19272 22154 19281
rect 22098 19207 22154 19216
rect 22836 19236 22888 19242
rect 22008 19168 22060 19174
rect 22008 19110 22060 19116
rect 22020 18766 22048 19110
rect 22008 18760 22060 18766
rect 22008 18702 22060 18708
rect 22112 17490 22140 19207
rect 22836 19178 22888 19184
rect 22848 18834 22876 19178
rect 22836 18828 22888 18834
rect 22836 18770 22888 18776
rect 22020 17462 22140 17490
rect 22020 17270 22048 17462
rect 22100 17332 22152 17338
rect 22100 17274 22152 17280
rect 22008 17264 22060 17270
rect 22008 17206 22060 17212
rect 22112 13258 22140 17274
rect 22836 16108 22888 16114
rect 22836 16050 22888 16056
rect 22848 15638 22876 16050
rect 22836 15632 22888 15638
rect 22836 15574 22888 15580
rect 22652 14952 22704 14958
rect 22652 14894 22704 14900
rect 22664 14006 22692 14894
rect 22652 14000 22704 14006
rect 22652 13942 22704 13948
rect 22664 13394 22692 13942
rect 22652 13388 22704 13394
rect 22652 13330 22704 13336
rect 22100 13252 22152 13258
rect 22100 13194 22152 13200
rect 22940 12434 22968 19332
rect 23020 19304 23072 19310
rect 23020 19246 23072 19252
rect 23032 18902 23060 19246
rect 23020 18896 23072 18902
rect 23020 18838 23072 18844
rect 23756 18624 23808 18630
rect 23756 18566 23808 18572
rect 23572 18352 23624 18358
rect 23572 18294 23624 18300
rect 23664 18352 23716 18358
rect 23664 18294 23716 18300
rect 23204 17740 23256 17746
rect 23204 17682 23256 17688
rect 23020 17128 23072 17134
rect 23020 17070 23072 17076
rect 23032 16794 23060 17070
rect 23112 17060 23164 17066
rect 23112 17002 23164 17008
rect 23020 16788 23072 16794
rect 23020 16730 23072 16736
rect 23124 16046 23152 17002
rect 23216 16998 23244 17682
rect 23480 17604 23532 17610
rect 23480 17546 23532 17552
rect 23492 17202 23520 17546
rect 23480 17196 23532 17202
rect 23480 17138 23532 17144
rect 23204 16992 23256 16998
rect 23204 16934 23256 16940
rect 23112 16040 23164 16046
rect 23112 15982 23164 15988
rect 23216 15978 23244 16934
rect 23388 16788 23440 16794
rect 23388 16730 23440 16736
rect 23296 16516 23348 16522
rect 23296 16458 23348 16464
rect 23308 15978 23336 16458
rect 23400 16114 23428 16730
rect 23492 16590 23520 17138
rect 23480 16584 23532 16590
rect 23480 16526 23532 16532
rect 23388 16108 23440 16114
rect 23388 16050 23440 16056
rect 23480 16108 23532 16114
rect 23480 16050 23532 16056
rect 23204 15972 23256 15978
rect 23204 15914 23256 15920
rect 23296 15972 23348 15978
rect 23296 15914 23348 15920
rect 23308 15706 23336 15914
rect 23296 15700 23348 15706
rect 23296 15642 23348 15648
rect 23492 15502 23520 16050
rect 23480 15496 23532 15502
rect 23480 15438 23532 15444
rect 23388 13932 23440 13938
rect 23388 13874 23440 13880
rect 23204 13728 23256 13734
rect 23204 13670 23256 13676
rect 23216 13326 23244 13670
rect 23204 13320 23256 13326
rect 23204 13262 23256 13268
rect 23400 12986 23428 13874
rect 23388 12980 23440 12986
rect 23388 12922 23440 12928
rect 23296 12776 23348 12782
rect 23296 12718 23348 12724
rect 22848 12406 22968 12434
rect 22284 11892 22336 11898
rect 22284 11834 22336 11840
rect 21916 11824 21968 11830
rect 21916 11766 21968 11772
rect 21548 11688 21600 11694
rect 21548 11630 21600 11636
rect 21560 10742 21588 11630
rect 22296 10742 22324 11834
rect 22560 11756 22612 11762
rect 22560 11698 22612 11704
rect 22468 11552 22520 11558
rect 22468 11494 22520 11500
rect 22480 11218 22508 11494
rect 22468 11212 22520 11218
rect 22468 11154 22520 11160
rect 22376 11144 22428 11150
rect 22376 11086 22428 11092
rect 21548 10736 21600 10742
rect 21548 10678 21600 10684
rect 22284 10736 22336 10742
rect 22284 10678 22336 10684
rect 21456 10668 21508 10674
rect 21456 10610 21508 10616
rect 21824 10668 21876 10674
rect 21824 10610 21876 10616
rect 22192 10668 22244 10674
rect 22192 10610 22244 10616
rect 21468 9994 21496 10610
rect 21836 10266 21864 10610
rect 22204 10554 22232 10610
rect 22204 10526 22324 10554
rect 22192 10464 22244 10470
rect 22192 10406 22244 10412
rect 21824 10260 21876 10266
rect 21824 10202 21876 10208
rect 20812 9988 20864 9994
rect 20812 9930 20864 9936
rect 21456 9988 21508 9994
rect 21456 9930 21508 9936
rect 21272 9920 21324 9926
rect 21272 9862 21324 9868
rect 21284 9654 21312 9862
rect 20720 9648 20772 9654
rect 20720 9590 20772 9596
rect 21272 9648 21324 9654
rect 21272 9590 21324 9596
rect 22204 9586 22232 10406
rect 22296 9994 22324 10526
rect 22284 9988 22336 9994
rect 22284 9930 22336 9936
rect 22388 9722 22416 11086
rect 22480 10538 22508 11154
rect 22572 10810 22600 11698
rect 22560 10804 22612 10810
rect 22560 10746 22612 10752
rect 22744 10668 22796 10674
rect 22744 10610 22796 10616
rect 22468 10532 22520 10538
rect 22468 10474 22520 10480
rect 22756 10062 22784 10610
rect 22744 10056 22796 10062
rect 22744 9998 22796 10004
rect 22376 9716 22428 9722
rect 22376 9658 22428 9664
rect 22756 9586 22784 9998
rect 22192 9580 22244 9586
rect 22192 9522 22244 9528
rect 22744 9580 22796 9586
rect 22744 9522 22796 9528
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 22848 6914 22876 12406
rect 23308 12306 23336 12718
rect 23296 12300 23348 12306
rect 23296 12242 23348 12248
rect 22928 12164 22980 12170
rect 22928 12106 22980 12112
rect 22940 11354 22968 12106
rect 22928 11348 22980 11354
rect 22928 11290 22980 11296
rect 23388 11144 23440 11150
rect 23388 11086 23440 11092
rect 23400 10674 23428 11086
rect 23388 10668 23440 10674
rect 23388 10610 23440 10616
rect 23204 10464 23256 10470
rect 23204 10406 23256 10412
rect 23216 10130 23244 10406
rect 23204 10124 23256 10130
rect 23204 10066 23256 10072
rect 23204 9988 23256 9994
rect 23204 9930 23256 9936
rect 23216 9586 23244 9930
rect 23296 9920 23348 9926
rect 23296 9862 23348 9868
rect 23308 9586 23336 9862
rect 23204 9580 23256 9586
rect 23204 9522 23256 9528
rect 23296 9580 23348 9586
rect 23296 9522 23348 9528
rect 22848 6886 22968 6914
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 18236 4684 18288 4690
rect 18236 4626 18288 4632
rect 19432 4548 19484 4554
rect 19432 4490 19484 4496
rect 17592 3664 17644 3670
rect 17592 3606 17644 3612
rect 17604 3534 17632 3606
rect 19444 3534 19472 4490
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 20168 4004 20220 4010
rect 20168 3946 20220 3952
rect 20076 3936 20128 3942
rect 20076 3878 20128 3884
rect 16856 3528 16908 3534
rect 16856 3470 16908 3476
rect 17592 3528 17644 3534
rect 17592 3470 17644 3476
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19984 3528 20036 3534
rect 19984 3470 20036 3476
rect 13360 3120 13412 3126
rect 13360 3062 13412 3068
rect 16868 3058 16896 3470
rect 17040 3392 17092 3398
rect 17040 3334 17092 3340
rect 17052 3126 17080 3334
rect 17040 3120 17092 3126
rect 17040 3062 17092 3068
rect 13176 3052 13228 3058
rect 13176 2994 13228 3000
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 17408 2984 17460 2990
rect 17408 2926 17460 2932
rect 12624 2644 12676 2650
rect 12624 2586 12676 2592
rect 12900 2508 12952 2514
rect 12900 2450 12952 2456
rect 12532 2372 12584 2378
rect 12532 2314 12584 2320
rect 12912 800 12940 2450
rect 13556 800 13584 2926
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 14200 800 14228 2382
rect 17420 800 17448 2926
rect 19352 2514 19380 3470
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 19444 3126 19472 3334
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19432 3120 19484 3126
rect 19432 3062 19484 3068
rect 19340 2508 19392 2514
rect 19340 2450 19392 2456
rect 19616 2508 19668 2514
rect 19616 2450 19668 2456
rect 19628 2394 19656 2450
rect 19352 2366 19656 2394
rect 19352 800 19380 2366
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19996 800 20024 3470
rect 20088 2990 20116 3878
rect 20076 2984 20128 2990
rect 20076 2926 20128 2932
rect 20180 2378 20208 3946
rect 20628 2984 20680 2990
rect 20628 2926 20680 2932
rect 20168 2372 20220 2378
rect 20168 2314 20220 2320
rect 20640 800 20668 2926
rect 22572 870 22784 898
rect 22572 800 22600 870
rect 2778 776 2834 785
rect 2778 711 2834 720
rect 3210 200 3322 800
rect 4498 200 4610 800
rect 5142 200 5254 800
rect 6430 200 6542 800
rect 7074 200 7186 800
rect 7718 200 7830 800
rect 9006 200 9118 800
rect 9650 200 9762 800
rect 10938 200 11050 800
rect 11582 200 11694 800
rect 12870 200 12982 800
rect 13514 200 13626 800
rect 14158 200 14270 800
rect 15446 200 15558 800
rect 16090 200 16202 800
rect 17378 200 17490 800
rect 18022 200 18134 800
rect 19310 200 19422 800
rect 19954 200 20066 800
rect 20598 200 20710 800
rect 21886 200 21998 800
rect 22530 200 22642 800
rect 22756 762 22784 870
rect 22940 762 22968 6886
rect 23584 2922 23612 18294
rect 23676 17882 23704 18294
rect 23664 17876 23716 17882
rect 23664 17818 23716 17824
rect 23768 17678 23796 18566
rect 23860 18086 23888 22102
rect 23940 18760 23992 18766
rect 23940 18702 23992 18708
rect 23952 18426 23980 18702
rect 23940 18420 23992 18426
rect 23940 18362 23992 18368
rect 24044 18290 24072 26302
rect 24676 26250 24728 26256
rect 24124 25288 24176 25294
rect 24124 25230 24176 25236
rect 24136 22642 24164 25230
rect 24584 22976 24636 22982
rect 24584 22918 24636 22924
rect 24596 22710 24624 22918
rect 24584 22704 24636 22710
rect 24584 22646 24636 22652
rect 24124 22636 24176 22642
rect 24124 22578 24176 22584
rect 24136 22030 24164 22578
rect 24688 22030 24716 26250
rect 24872 24886 24900 26726
rect 24952 25900 25004 25906
rect 24952 25842 25004 25848
rect 24964 25498 24992 25842
rect 24952 25492 25004 25498
rect 24952 25434 25004 25440
rect 25056 25378 25084 28018
rect 25228 27872 25280 27878
rect 25228 27814 25280 27820
rect 25240 27402 25268 27814
rect 25228 27396 25280 27402
rect 25228 27338 25280 27344
rect 25424 27130 25452 28018
rect 25412 27124 25464 27130
rect 25412 27066 25464 27072
rect 25228 26376 25280 26382
rect 25228 26318 25280 26324
rect 25240 26042 25268 26318
rect 25594 26208 25650 26217
rect 25594 26143 25650 26152
rect 25228 26036 25280 26042
rect 25228 25978 25280 25984
rect 25608 25838 25636 26143
rect 25700 25906 25728 31282
rect 25780 30252 25832 30258
rect 25780 30194 25832 30200
rect 25792 30122 25820 30194
rect 25780 30116 25832 30122
rect 25780 30058 25832 30064
rect 25780 29640 25832 29646
rect 25780 29582 25832 29588
rect 25792 29102 25820 29582
rect 25780 29096 25832 29102
rect 25780 29038 25832 29044
rect 25792 27674 25820 29038
rect 25884 28626 25912 31282
rect 25976 30734 26004 31583
rect 25964 30728 26016 30734
rect 25964 30670 26016 30676
rect 25964 30184 26016 30190
rect 25964 30126 26016 30132
rect 25976 29714 26004 30126
rect 25964 29708 26016 29714
rect 25964 29650 26016 29656
rect 25872 28620 25924 28626
rect 25872 28562 25924 28568
rect 25780 27668 25832 27674
rect 25780 27610 25832 27616
rect 25964 27600 26016 27606
rect 25964 27542 26016 27548
rect 25976 26994 26004 27542
rect 25964 26988 26016 26994
rect 25964 26930 26016 26936
rect 26160 26382 26188 32370
rect 26240 30592 26292 30598
rect 26240 30534 26292 30540
rect 26252 29646 26280 30534
rect 26240 29640 26292 29646
rect 26240 29582 26292 29588
rect 26240 27940 26292 27946
rect 26240 27882 26292 27888
rect 26252 26586 26280 27882
rect 26240 26580 26292 26586
rect 26240 26522 26292 26528
rect 26148 26376 26200 26382
rect 26200 26324 26372 26330
rect 26148 26318 26372 26324
rect 26160 26302 26372 26318
rect 25688 25900 25740 25906
rect 25688 25842 25740 25848
rect 25596 25832 25648 25838
rect 25596 25774 25648 25780
rect 24964 25350 25084 25378
rect 25608 25362 25636 25774
rect 25596 25356 25648 25362
rect 24860 24880 24912 24886
rect 24860 24822 24912 24828
rect 24768 23112 24820 23118
rect 24768 23054 24820 23060
rect 24780 22234 24808 23054
rect 24872 22234 24900 24822
rect 24768 22228 24820 22234
rect 24768 22170 24820 22176
rect 24860 22228 24912 22234
rect 24860 22170 24912 22176
rect 24964 22094 24992 25350
rect 25596 25298 25648 25304
rect 25504 23656 25556 23662
rect 25504 23598 25556 23604
rect 25044 23112 25096 23118
rect 25044 23054 25096 23060
rect 25056 22438 25084 23054
rect 25516 22438 25544 23598
rect 25044 22432 25096 22438
rect 25044 22374 25096 22380
rect 25504 22432 25556 22438
rect 25504 22374 25556 22380
rect 24872 22066 24992 22094
rect 24124 22024 24176 22030
rect 24124 21966 24176 21972
rect 24676 22024 24728 22030
rect 24676 21966 24728 21972
rect 24308 21548 24360 21554
rect 24308 21490 24360 21496
rect 24320 21146 24348 21490
rect 24688 21350 24716 21966
rect 24676 21344 24728 21350
rect 24676 21286 24728 21292
rect 24308 21140 24360 21146
rect 24308 21082 24360 21088
rect 24768 19168 24820 19174
rect 24768 19110 24820 19116
rect 24780 18766 24808 19110
rect 24768 18760 24820 18766
rect 24768 18702 24820 18708
rect 24780 18290 24808 18702
rect 24872 18698 24900 22066
rect 24952 22024 25004 22030
rect 24952 21966 25004 21972
rect 24964 21690 24992 21966
rect 24952 21684 25004 21690
rect 24952 21626 25004 21632
rect 25056 21554 25084 22374
rect 25516 22030 25544 22374
rect 25504 22024 25556 22030
rect 25504 21966 25556 21972
rect 25044 21548 25096 21554
rect 25044 21490 25096 21496
rect 25228 20936 25280 20942
rect 25280 20884 25360 20890
rect 25228 20878 25360 20884
rect 25240 20862 25360 20878
rect 25228 19848 25280 19854
rect 25228 19790 25280 19796
rect 25240 19530 25268 19790
rect 25148 19514 25268 19530
rect 25148 19508 25280 19514
rect 25148 19502 25228 19508
rect 25044 18964 25096 18970
rect 25044 18906 25096 18912
rect 24860 18692 24912 18698
rect 24860 18634 24912 18640
rect 24032 18284 24084 18290
rect 24032 18226 24084 18232
rect 24768 18284 24820 18290
rect 24768 18226 24820 18232
rect 24872 18154 24900 18634
rect 25056 18426 25084 18906
rect 25148 18630 25176 19502
rect 25228 19450 25280 19456
rect 25228 19372 25280 19378
rect 25228 19314 25280 19320
rect 25240 18970 25268 19314
rect 25228 18964 25280 18970
rect 25228 18906 25280 18912
rect 25228 18760 25280 18766
rect 25228 18702 25280 18708
rect 25136 18624 25188 18630
rect 25136 18566 25188 18572
rect 25044 18420 25096 18426
rect 25044 18362 25096 18368
rect 25148 18358 25176 18566
rect 25136 18352 25188 18358
rect 25136 18294 25188 18300
rect 24860 18148 24912 18154
rect 24860 18090 24912 18096
rect 23848 18080 23900 18086
rect 23848 18022 23900 18028
rect 23940 18080 23992 18086
rect 23940 18022 23992 18028
rect 23756 17672 23808 17678
rect 23756 17614 23808 17620
rect 23664 13864 23716 13870
rect 23664 13806 23716 13812
rect 23676 11082 23704 13806
rect 23756 13252 23808 13258
rect 23756 13194 23808 13200
rect 23768 12850 23796 13194
rect 23756 12844 23808 12850
rect 23756 12786 23808 12792
rect 23860 12306 23888 18022
rect 23952 17678 23980 18022
rect 23940 17672 23992 17678
rect 23940 17614 23992 17620
rect 23952 17134 23980 17614
rect 23940 17128 23992 17134
rect 23940 17070 23992 17076
rect 24032 16992 24084 16998
rect 24032 16934 24084 16940
rect 24044 16046 24072 16934
rect 24872 16658 24900 18090
rect 24860 16652 24912 16658
rect 24860 16594 24912 16600
rect 25240 16590 25268 18702
rect 25228 16584 25280 16590
rect 25228 16526 25280 16532
rect 25228 16448 25280 16454
rect 25228 16390 25280 16396
rect 25240 16114 25268 16390
rect 25228 16108 25280 16114
rect 25228 16050 25280 16056
rect 24032 16040 24084 16046
rect 24032 15982 24084 15988
rect 25332 14906 25360 20862
rect 25608 18766 25636 25298
rect 25872 25220 25924 25226
rect 25872 25162 25924 25168
rect 25884 24818 25912 25162
rect 26240 25152 26292 25158
rect 26240 25094 26292 25100
rect 26252 24818 26280 25094
rect 25872 24812 25924 24818
rect 25872 24754 25924 24760
rect 26240 24812 26292 24818
rect 26240 24754 26292 24760
rect 25884 24206 25912 24754
rect 26148 24676 26200 24682
rect 26148 24618 26200 24624
rect 26160 24410 26188 24618
rect 26148 24404 26200 24410
rect 26148 24346 26200 24352
rect 25872 24200 25924 24206
rect 25872 24142 25924 24148
rect 25688 19712 25740 19718
rect 25688 19654 25740 19660
rect 25596 18760 25648 18766
rect 25596 18702 25648 18708
rect 25596 16584 25648 16590
rect 25596 16526 25648 16532
rect 25412 15904 25464 15910
rect 25412 15846 25464 15852
rect 25424 15094 25452 15846
rect 25608 15638 25636 16526
rect 25596 15632 25648 15638
rect 25596 15574 25648 15580
rect 25504 15564 25556 15570
rect 25504 15506 25556 15512
rect 25412 15088 25464 15094
rect 25412 15030 25464 15036
rect 25332 14878 25452 14906
rect 24032 13184 24084 13190
rect 24032 13126 24084 13132
rect 24044 12850 24072 13126
rect 25320 12980 25372 12986
rect 25320 12922 25372 12928
rect 24032 12844 24084 12850
rect 24032 12786 24084 12792
rect 23848 12300 23900 12306
rect 23848 12242 23900 12248
rect 23860 11762 23888 12242
rect 24044 12238 24072 12786
rect 24032 12232 24084 12238
rect 24032 12174 24084 12180
rect 25332 11898 25360 12922
rect 25424 12434 25452 14878
rect 25516 14278 25544 15506
rect 25608 15502 25636 15574
rect 25596 15496 25648 15502
rect 25596 15438 25648 15444
rect 25608 14890 25636 15438
rect 25596 14884 25648 14890
rect 25596 14826 25648 14832
rect 25700 14482 25728 19654
rect 25780 15020 25832 15026
rect 25780 14962 25832 14968
rect 25688 14476 25740 14482
rect 25688 14418 25740 14424
rect 25504 14272 25556 14278
rect 25504 14214 25556 14220
rect 25516 14006 25544 14214
rect 25504 14000 25556 14006
rect 25504 13942 25556 13948
rect 25700 13938 25728 14418
rect 25792 14074 25820 14962
rect 25780 14068 25832 14074
rect 25780 14010 25832 14016
rect 25688 13932 25740 13938
rect 25688 13874 25740 13880
rect 25884 13258 25912 24142
rect 26056 24064 26108 24070
rect 26056 24006 26108 24012
rect 26068 19786 26096 24006
rect 26160 21146 26188 24346
rect 26344 23866 26372 26302
rect 26528 25974 26556 32370
rect 28368 31346 28396 32438
rect 28356 31340 28408 31346
rect 28356 31282 28408 31288
rect 28908 31340 28960 31346
rect 28908 31282 28960 31288
rect 28920 30938 28948 31282
rect 28908 30932 28960 30938
rect 28908 30874 28960 30880
rect 27344 30796 27396 30802
rect 27344 30738 27396 30744
rect 27356 30258 27384 30738
rect 27344 30252 27396 30258
rect 27344 30194 27396 30200
rect 27356 29782 27384 30194
rect 27528 30184 27580 30190
rect 27528 30126 27580 30132
rect 27344 29776 27396 29782
rect 27344 29718 27396 29724
rect 27356 29102 27384 29718
rect 27540 29170 27568 30126
rect 29000 30116 29052 30122
rect 29000 30058 29052 30064
rect 27620 29504 27672 29510
rect 27620 29446 27672 29452
rect 27528 29164 27580 29170
rect 27528 29106 27580 29112
rect 27344 29096 27396 29102
rect 27344 29038 27396 29044
rect 27160 27872 27212 27878
rect 27160 27814 27212 27820
rect 27172 27402 27200 27814
rect 27160 27396 27212 27402
rect 27160 27338 27212 27344
rect 27540 27334 27568 29106
rect 27632 28014 27660 29446
rect 28816 28960 28868 28966
rect 28816 28902 28868 28908
rect 27804 28076 27856 28082
rect 27804 28018 27856 28024
rect 27620 28008 27672 28014
rect 27620 27950 27672 27956
rect 27528 27328 27580 27334
rect 27528 27270 27580 27276
rect 27540 27062 27568 27270
rect 27816 27130 27844 28018
rect 28828 28014 28856 28902
rect 28816 28008 28868 28014
rect 28816 27950 28868 27956
rect 28828 27470 28856 27950
rect 28816 27464 28868 27470
rect 28816 27406 28868 27412
rect 27804 27124 27856 27130
rect 27804 27066 27856 27072
rect 27528 27056 27580 27062
rect 27528 26998 27580 27004
rect 26884 26920 26936 26926
rect 26884 26862 26936 26868
rect 26896 26314 26924 26862
rect 26976 26580 27028 26586
rect 26976 26522 27028 26528
rect 26884 26308 26936 26314
rect 26884 26250 26936 26256
rect 26516 25968 26568 25974
rect 26516 25910 26568 25916
rect 26424 25696 26476 25702
rect 26424 25638 26476 25644
rect 26436 25294 26464 25638
rect 26424 25288 26476 25294
rect 26424 25230 26476 25236
rect 26332 23860 26384 23866
rect 26332 23802 26384 23808
rect 26528 22098 26556 25910
rect 26792 24200 26844 24206
rect 26792 24142 26844 24148
rect 26700 24064 26752 24070
rect 26700 24006 26752 24012
rect 26608 23520 26660 23526
rect 26608 23462 26660 23468
rect 26620 23050 26648 23462
rect 26712 23322 26740 24006
rect 26700 23316 26752 23322
rect 26700 23258 26752 23264
rect 26608 23044 26660 23050
rect 26608 22986 26660 22992
rect 26620 22642 26648 22986
rect 26804 22710 26832 24142
rect 26792 22704 26844 22710
rect 26792 22646 26844 22652
rect 26608 22636 26660 22642
rect 26608 22578 26660 22584
rect 26516 22092 26568 22098
rect 26516 22034 26568 22040
rect 26240 22024 26292 22030
rect 26240 21966 26292 21972
rect 26252 21690 26280 21966
rect 26424 21888 26476 21894
rect 26424 21830 26476 21836
rect 26240 21684 26292 21690
rect 26240 21626 26292 21632
rect 26252 21146 26280 21626
rect 26436 21554 26464 21830
rect 26424 21548 26476 21554
rect 26424 21490 26476 21496
rect 26528 21486 26556 22034
rect 26620 21894 26648 22578
rect 26896 22094 26924 26250
rect 26988 23186 27016 26522
rect 27160 25900 27212 25906
rect 27160 25842 27212 25848
rect 27172 24682 27200 25842
rect 27344 25152 27396 25158
rect 27344 25094 27396 25100
rect 27356 24954 27384 25094
rect 27344 24948 27396 24954
rect 27344 24890 27396 24896
rect 27436 24812 27488 24818
rect 27436 24754 27488 24760
rect 27160 24676 27212 24682
rect 27160 24618 27212 24624
rect 27448 24410 27476 24754
rect 29012 24682 29040 30058
rect 29104 29510 29132 33322
rect 29656 33318 29684 44134
rect 29840 43314 29868 45426
rect 29828 43308 29880 43314
rect 29828 43250 29880 43256
rect 32404 35692 32456 35698
rect 32404 35634 32456 35640
rect 32312 35216 32364 35222
rect 32312 35158 32364 35164
rect 32324 35086 32352 35158
rect 29736 35080 29788 35086
rect 29736 35022 29788 35028
rect 30472 35080 30524 35086
rect 30472 35022 30524 35028
rect 32312 35080 32364 35086
rect 32312 35022 32364 35028
rect 29644 33312 29696 33318
rect 29644 33254 29696 33260
rect 29748 32978 29776 35022
rect 30196 35012 30248 35018
rect 30196 34954 30248 34960
rect 30208 34406 30236 34954
rect 30484 34610 30512 35022
rect 31208 34944 31260 34950
rect 31208 34886 31260 34892
rect 30472 34604 30524 34610
rect 30472 34546 30524 34552
rect 30748 34604 30800 34610
rect 30748 34546 30800 34552
rect 30932 34604 30984 34610
rect 30932 34546 30984 34552
rect 30196 34400 30248 34406
rect 30196 34342 30248 34348
rect 30208 33998 30236 34342
rect 30104 33992 30156 33998
rect 30104 33934 30156 33940
rect 30196 33992 30248 33998
rect 30196 33934 30248 33940
rect 30380 33992 30432 33998
rect 30380 33934 30432 33940
rect 30012 33856 30064 33862
rect 30012 33798 30064 33804
rect 29736 32972 29788 32978
rect 29736 32914 29788 32920
rect 30024 32910 30052 33798
rect 30116 33658 30144 33934
rect 30104 33652 30156 33658
rect 30104 33594 30156 33600
rect 30012 32904 30064 32910
rect 30012 32846 30064 32852
rect 30208 32722 30236 33934
rect 30392 33114 30420 33934
rect 30484 33522 30512 34546
rect 30760 33590 30788 34546
rect 30748 33584 30800 33590
rect 30748 33526 30800 33532
rect 30472 33516 30524 33522
rect 30472 33458 30524 33464
rect 30380 33108 30432 33114
rect 30380 33050 30432 33056
rect 30024 32694 30236 32722
rect 29736 31748 29788 31754
rect 29736 31690 29788 31696
rect 29748 31142 29776 31690
rect 29736 31136 29788 31142
rect 29736 31078 29788 31084
rect 29748 30258 29776 31078
rect 29828 30592 29880 30598
rect 29828 30534 29880 30540
rect 29736 30252 29788 30258
rect 29736 30194 29788 30200
rect 29644 29708 29696 29714
rect 29644 29650 29696 29656
rect 29092 29504 29144 29510
rect 29092 29446 29144 29452
rect 29104 28626 29132 29446
rect 29656 29306 29684 29650
rect 29840 29646 29868 30534
rect 29828 29640 29880 29646
rect 29828 29582 29880 29588
rect 29840 29306 29868 29582
rect 29644 29300 29696 29306
rect 29644 29242 29696 29248
rect 29828 29300 29880 29306
rect 29828 29242 29880 29248
rect 29092 28620 29144 28626
rect 29092 28562 29144 28568
rect 29656 27470 29684 29242
rect 29920 28552 29972 28558
rect 29920 28494 29972 28500
rect 29736 28416 29788 28422
rect 29736 28358 29788 28364
rect 29748 28150 29776 28358
rect 29736 28144 29788 28150
rect 29736 28086 29788 28092
rect 29932 27674 29960 28494
rect 29920 27668 29972 27674
rect 29920 27610 29972 27616
rect 30024 27538 30052 32694
rect 30288 31136 30340 31142
rect 30288 31078 30340 31084
rect 30196 30592 30248 30598
rect 30196 30534 30248 30540
rect 30208 30394 30236 30534
rect 30196 30388 30248 30394
rect 30196 30330 30248 30336
rect 30300 30190 30328 31078
rect 30288 30184 30340 30190
rect 30288 30126 30340 30132
rect 30104 29640 30156 29646
rect 30104 29582 30156 29588
rect 30116 29034 30144 29582
rect 30472 29504 30524 29510
rect 30472 29446 30524 29452
rect 30484 29170 30512 29446
rect 30944 29170 30972 34546
rect 31220 34542 31248 34886
rect 32324 34678 32352 35022
rect 32312 34672 32364 34678
rect 32312 34614 32364 34620
rect 31024 34536 31076 34542
rect 31024 34478 31076 34484
rect 31208 34536 31260 34542
rect 31208 34478 31260 34484
rect 31036 32502 31064 34478
rect 31208 34196 31260 34202
rect 31208 34138 31260 34144
rect 31220 33522 31248 34138
rect 32324 33810 32352 34614
rect 32416 34542 32444 35634
rect 32508 34610 32536 46854
rect 33152 46714 33180 46990
rect 33140 46708 33192 46714
rect 33140 46650 33192 46656
rect 33520 46510 33548 49200
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 33232 46504 33284 46510
rect 33232 46446 33284 46452
rect 33508 46504 33560 46510
rect 33508 46446 33560 46452
rect 33244 46170 33272 46446
rect 35348 46368 35400 46374
rect 35348 46310 35400 46316
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 33232 46164 33284 46170
rect 33232 46106 33284 46112
rect 35360 46034 35388 46310
rect 36096 46034 36124 49200
rect 36740 46442 36768 49200
rect 37648 46504 37700 46510
rect 37648 46446 37700 46452
rect 36728 46436 36780 46442
rect 36728 46378 36780 46384
rect 35348 46028 35400 46034
rect 35348 45970 35400 45976
rect 36084 46028 36136 46034
rect 36084 45970 36136 45976
rect 33140 45960 33192 45966
rect 33140 45902 33192 45908
rect 33152 44334 33180 45902
rect 35624 45892 35676 45898
rect 35624 45834 35676 45840
rect 35636 45558 35664 45834
rect 37660 45558 37688 46446
rect 38672 46442 38700 49200
rect 39764 47116 39816 47122
rect 39764 47058 39816 47064
rect 38936 47048 38988 47054
rect 38936 46990 38988 46996
rect 38660 46436 38712 46442
rect 38660 46378 38712 46384
rect 38292 45960 38344 45966
rect 38292 45902 38344 45908
rect 38384 45960 38436 45966
rect 38384 45902 38436 45908
rect 35624 45552 35676 45558
rect 35624 45494 35676 45500
rect 37648 45552 37700 45558
rect 37648 45494 37700 45500
rect 38304 45490 38332 45902
rect 38396 45626 38424 45902
rect 38384 45620 38436 45626
rect 38384 45562 38436 45568
rect 38948 45490 38976 46990
rect 39776 46578 39804 47058
rect 40132 47048 40184 47054
rect 40132 46990 40184 46996
rect 39764 46572 39816 46578
rect 39764 46514 39816 46520
rect 39948 46504 40000 46510
rect 39948 46446 40000 46452
rect 39960 46170 39988 46446
rect 39948 46164 40000 46170
rect 39948 46106 40000 46112
rect 40144 46034 40172 46990
rect 40604 46034 40632 49200
rect 41512 47048 41564 47054
rect 41512 46990 41564 46996
rect 41524 46578 41552 46990
rect 41512 46572 41564 46578
rect 41512 46514 41564 46520
rect 41892 46442 41920 49200
rect 42536 47054 42564 49200
rect 43628 47184 43680 47190
rect 43628 47126 43680 47132
rect 42524 47048 42576 47054
rect 42524 46990 42576 46996
rect 42800 46504 42852 46510
rect 42800 46446 42852 46452
rect 41880 46436 41932 46442
rect 41880 46378 41932 46384
rect 40132 46028 40184 46034
rect 40132 45970 40184 45976
rect 40592 46028 40644 46034
rect 40592 45970 40644 45976
rect 40316 45892 40368 45898
rect 40316 45834 40368 45840
rect 39120 45824 39172 45830
rect 39120 45766 39172 45772
rect 39132 45558 39160 45766
rect 39120 45552 39172 45558
rect 39120 45494 39172 45500
rect 37280 45484 37332 45490
rect 37280 45426 37332 45432
rect 38292 45484 38344 45490
rect 38292 45426 38344 45432
rect 38936 45484 38988 45490
rect 38936 45426 38988 45432
rect 35716 45280 35768 45286
rect 35716 45222 35768 45228
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 33140 44328 33192 44334
rect 33140 44270 33192 44276
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 35728 38962 35756 45222
rect 37292 44402 37320 45426
rect 40132 45416 40184 45422
rect 40132 45358 40184 45364
rect 40144 45082 40172 45358
rect 40328 45082 40356 45834
rect 42812 45558 42840 46446
rect 42800 45552 42852 45558
rect 42800 45494 42852 45500
rect 40132 45076 40184 45082
rect 40132 45018 40184 45024
rect 40316 45076 40368 45082
rect 40316 45018 40368 45024
rect 37280 44396 37332 44402
rect 37280 44338 37332 44344
rect 35716 38956 35768 38962
rect 35716 38898 35768 38904
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 33048 35692 33100 35698
rect 33048 35634 33100 35640
rect 34796 35692 34848 35698
rect 34796 35634 34848 35640
rect 33060 35290 33088 35634
rect 34704 35624 34756 35630
rect 34704 35566 34756 35572
rect 33508 35488 33560 35494
rect 33508 35430 33560 35436
rect 33048 35284 33100 35290
rect 33048 35226 33100 35232
rect 33520 35154 33548 35430
rect 33508 35148 33560 35154
rect 33508 35090 33560 35096
rect 32680 35012 32732 35018
rect 32680 34954 32732 34960
rect 32496 34604 32548 34610
rect 32496 34546 32548 34552
rect 32404 34536 32456 34542
rect 32404 34478 32456 34484
rect 32416 34066 32444 34478
rect 32404 34060 32456 34066
rect 32404 34002 32456 34008
rect 32324 33782 32628 33810
rect 31208 33516 31260 33522
rect 31208 33458 31260 33464
rect 31024 32496 31076 32502
rect 31024 32438 31076 32444
rect 31036 32026 31064 32438
rect 31024 32020 31076 32026
rect 31024 31962 31076 31968
rect 31036 31822 31064 31962
rect 31024 31816 31076 31822
rect 31024 31758 31076 31764
rect 31036 31414 31064 31758
rect 31024 31408 31076 31414
rect 31024 31350 31076 31356
rect 31024 29640 31076 29646
rect 31024 29582 31076 29588
rect 31036 29170 31064 29582
rect 30472 29164 30524 29170
rect 30472 29106 30524 29112
rect 30932 29164 30984 29170
rect 30932 29106 30984 29112
rect 31024 29164 31076 29170
rect 31024 29106 31076 29112
rect 30656 29096 30708 29102
rect 30656 29038 30708 29044
rect 30104 29028 30156 29034
rect 30104 28970 30156 28976
rect 30012 27532 30064 27538
rect 30012 27474 30064 27480
rect 29644 27464 29696 27470
rect 29644 27406 29696 27412
rect 29552 25696 29604 25702
rect 29552 25638 29604 25644
rect 29564 25294 29592 25638
rect 29656 25498 29684 27406
rect 29644 25492 29696 25498
rect 29644 25434 29696 25440
rect 29552 25288 29604 25294
rect 29552 25230 29604 25236
rect 29000 24676 29052 24682
rect 29000 24618 29052 24624
rect 29012 24410 29040 24618
rect 27436 24404 27488 24410
rect 27436 24346 27488 24352
rect 29000 24404 29052 24410
rect 29000 24346 29052 24352
rect 27620 24268 27672 24274
rect 27620 24210 27672 24216
rect 27632 24138 27660 24210
rect 28540 24200 28592 24206
rect 28540 24142 28592 24148
rect 27620 24132 27672 24138
rect 27620 24074 27672 24080
rect 28448 24132 28500 24138
rect 28448 24074 28500 24080
rect 27632 23662 27660 24074
rect 28460 23866 28488 24074
rect 28448 23860 28500 23866
rect 28448 23802 28500 23808
rect 27712 23724 27764 23730
rect 27712 23666 27764 23672
rect 27160 23656 27212 23662
rect 27160 23598 27212 23604
rect 27620 23656 27672 23662
rect 27620 23598 27672 23604
rect 26976 23180 27028 23186
rect 26976 23122 27028 23128
rect 27172 22137 27200 23598
rect 27632 23202 27660 23598
rect 27724 23254 27752 23666
rect 27804 23520 27856 23526
rect 27804 23462 27856 23468
rect 27540 23174 27660 23202
rect 27712 23248 27764 23254
rect 27712 23190 27764 23196
rect 27344 23112 27396 23118
rect 27540 23066 27568 23174
rect 27396 23060 27568 23066
rect 27344 23054 27568 23060
rect 27620 23112 27672 23118
rect 27620 23054 27672 23060
rect 27356 23038 27568 23054
rect 27540 22778 27568 23038
rect 27528 22772 27580 22778
rect 27528 22714 27580 22720
rect 27344 22704 27396 22710
rect 27344 22646 27396 22652
rect 27356 22574 27384 22646
rect 27436 22636 27488 22642
rect 27436 22578 27488 22584
rect 27344 22568 27396 22574
rect 27344 22510 27396 22516
rect 27252 22228 27304 22234
rect 27252 22170 27304 22176
rect 26804 22066 26924 22094
rect 27158 22128 27214 22137
rect 26804 22030 26832 22066
rect 27158 22063 27214 22072
rect 26792 22024 26844 22030
rect 26792 21966 26844 21972
rect 26608 21888 26660 21894
rect 26608 21830 26660 21836
rect 27264 21622 27292 22170
rect 26700 21616 26752 21622
rect 26700 21558 26752 21564
rect 27068 21616 27120 21622
rect 27068 21558 27120 21564
rect 27252 21616 27304 21622
rect 27252 21558 27304 21564
rect 26516 21480 26568 21486
rect 26516 21422 26568 21428
rect 26332 21412 26384 21418
rect 26332 21354 26384 21360
rect 26148 21140 26200 21146
rect 26148 21082 26200 21088
rect 26240 21140 26292 21146
rect 26240 21082 26292 21088
rect 26344 20942 26372 21354
rect 26332 20936 26384 20942
rect 26332 20878 26384 20884
rect 26344 19922 26372 20878
rect 26712 20806 26740 21558
rect 27080 20942 27108 21558
rect 27356 21554 27384 22510
rect 27448 22234 27476 22578
rect 27436 22228 27488 22234
rect 27436 22170 27488 22176
rect 27434 22128 27490 22137
rect 27632 22094 27660 23054
rect 27816 23050 27844 23462
rect 28552 23118 28580 24142
rect 28448 23112 28500 23118
rect 28448 23054 28500 23060
rect 28540 23112 28592 23118
rect 28540 23054 28592 23060
rect 27804 23044 27856 23050
rect 27804 22986 27856 22992
rect 27712 22772 27764 22778
rect 27712 22714 27764 22720
rect 27724 22642 27752 22714
rect 27712 22636 27764 22642
rect 27712 22578 27764 22584
rect 27724 22166 27752 22578
rect 27712 22160 27764 22166
rect 27712 22102 27764 22108
rect 27434 22063 27490 22072
rect 27540 22066 27660 22094
rect 27344 21548 27396 21554
rect 27344 21490 27396 21496
rect 27356 20942 27384 21490
rect 27068 20936 27120 20942
rect 27068 20878 27120 20884
rect 27344 20936 27396 20942
rect 27344 20878 27396 20884
rect 26700 20800 26752 20806
rect 26700 20742 26752 20748
rect 27252 20800 27304 20806
rect 27252 20742 27304 20748
rect 26332 19916 26384 19922
rect 26332 19858 26384 19864
rect 26056 19780 26108 19786
rect 26056 19722 26108 19728
rect 26148 15904 26200 15910
rect 26148 15846 26200 15852
rect 26160 15434 26188 15846
rect 26148 15428 26200 15434
rect 26148 15370 26200 15376
rect 26240 14816 26292 14822
rect 26240 14758 26292 14764
rect 26252 14414 26280 14758
rect 26240 14408 26292 14414
rect 26240 14350 26292 14356
rect 26344 14226 26372 19858
rect 27160 18624 27212 18630
rect 27160 18566 27212 18572
rect 27172 18290 27200 18566
rect 27264 18290 27292 20742
rect 27344 19712 27396 19718
rect 27344 19654 27396 19660
rect 27356 19378 27384 19654
rect 27448 19378 27476 22063
rect 27540 22030 27568 22066
rect 27816 22030 27844 22986
rect 28460 22642 28488 23054
rect 28552 22710 28580 23054
rect 28540 22704 28592 22710
rect 28540 22646 28592 22652
rect 28448 22636 28500 22642
rect 28448 22578 28500 22584
rect 28632 22432 28684 22438
rect 28632 22374 28684 22380
rect 27528 22024 27580 22030
rect 27528 21966 27580 21972
rect 27804 22024 27856 22030
rect 27804 21966 27856 21972
rect 27540 21350 27568 21966
rect 28080 21888 28132 21894
rect 28080 21830 28132 21836
rect 27712 21480 27764 21486
rect 27712 21422 27764 21428
rect 27528 21344 27580 21350
rect 27528 21286 27580 21292
rect 27540 21146 27568 21286
rect 27528 21140 27580 21146
rect 27528 21082 27580 21088
rect 27620 20800 27672 20806
rect 27620 20742 27672 20748
rect 27632 20466 27660 20742
rect 27724 20466 27752 21422
rect 28092 20942 28120 21830
rect 28644 21622 28672 22374
rect 29012 21978 29040 24346
rect 29276 23520 29328 23526
rect 29276 23462 29328 23468
rect 29288 23254 29316 23462
rect 29276 23248 29328 23254
rect 29276 23190 29328 23196
rect 29288 22438 29316 23190
rect 30024 22710 30052 27474
rect 30116 27470 30144 28970
rect 30668 28626 30696 29038
rect 30656 28620 30708 28626
rect 30656 28562 30708 28568
rect 30380 28212 30432 28218
rect 30380 28154 30432 28160
rect 30392 27470 30420 28154
rect 30944 28082 30972 29106
rect 30932 28076 30984 28082
rect 30932 28018 30984 28024
rect 30104 27464 30156 27470
rect 30104 27406 30156 27412
rect 30380 27464 30432 27470
rect 30380 27406 30432 27412
rect 30116 26330 30144 27406
rect 30116 26302 30328 26330
rect 30196 25696 30248 25702
rect 30196 25638 30248 25644
rect 30208 25226 30236 25638
rect 30300 25294 30328 26302
rect 31116 26240 31168 26246
rect 31116 26182 31168 26188
rect 31128 25838 31156 26182
rect 31220 26024 31248 33458
rect 31392 33108 31444 33114
rect 31392 33050 31444 33056
rect 31404 32434 31432 33050
rect 31576 32836 31628 32842
rect 31576 32778 31628 32784
rect 31392 32428 31444 32434
rect 31392 32370 31444 32376
rect 31588 32366 31616 32778
rect 31668 32428 31720 32434
rect 31668 32370 31720 32376
rect 31576 32360 31628 32366
rect 31576 32302 31628 32308
rect 31300 31952 31352 31958
rect 31300 31894 31352 31900
rect 31312 31346 31340 31894
rect 31588 31754 31616 32302
rect 31680 31822 31708 32370
rect 31760 32360 31812 32366
rect 31760 32302 31812 32308
rect 31772 31890 31800 32302
rect 31760 31884 31812 31890
rect 31760 31826 31812 31832
rect 31668 31816 31720 31822
rect 31668 31758 31720 31764
rect 31496 31726 31616 31754
rect 31300 31340 31352 31346
rect 31300 31282 31352 31288
rect 31496 28762 31524 31726
rect 31576 31680 31628 31686
rect 31576 31622 31628 31628
rect 31588 31346 31616 31622
rect 31576 31340 31628 31346
rect 31576 31282 31628 31288
rect 32496 30252 32548 30258
rect 32496 30194 32548 30200
rect 31944 30184 31996 30190
rect 31944 30126 31996 30132
rect 31576 30116 31628 30122
rect 31576 30058 31628 30064
rect 31588 29034 31616 30058
rect 31576 29028 31628 29034
rect 31576 28970 31628 28976
rect 31484 28756 31536 28762
rect 31484 28698 31536 28704
rect 31496 28558 31524 28698
rect 31588 28626 31616 28970
rect 31576 28620 31628 28626
rect 31576 28562 31628 28568
rect 31484 28552 31536 28558
rect 31484 28494 31536 28500
rect 31588 28506 31616 28562
rect 31588 28478 31708 28506
rect 31680 27946 31708 28478
rect 31668 27940 31720 27946
rect 31668 27882 31720 27888
rect 31680 26042 31708 27882
rect 31956 26518 31984 30126
rect 32312 30048 32364 30054
rect 32312 29990 32364 29996
rect 32324 29578 32352 29990
rect 32312 29572 32364 29578
rect 32312 29514 32364 29520
rect 32036 29232 32088 29238
rect 32404 29232 32456 29238
rect 32088 29180 32404 29186
rect 32036 29174 32456 29180
rect 32048 29158 32444 29174
rect 32508 28966 32536 30194
rect 32496 28960 32548 28966
rect 32496 28902 32548 28908
rect 32220 28756 32272 28762
rect 32220 28698 32272 28704
rect 32232 28490 32260 28698
rect 32220 28484 32272 28490
rect 32220 28426 32272 28432
rect 32036 26920 32088 26926
rect 32036 26862 32088 26868
rect 31944 26512 31996 26518
rect 31944 26454 31996 26460
rect 32048 26450 32076 26862
rect 32036 26444 32088 26450
rect 32036 26386 32088 26392
rect 32312 26308 32364 26314
rect 32312 26250 32364 26256
rect 31668 26036 31720 26042
rect 31220 25996 31616 26024
rect 31588 25922 31616 25996
rect 31668 25978 31720 25984
rect 31760 25968 31812 25974
rect 31588 25916 31760 25922
rect 31588 25910 31812 25916
rect 31208 25900 31260 25906
rect 31588 25894 31800 25910
rect 31208 25842 31260 25848
rect 31116 25832 31168 25838
rect 31116 25774 31168 25780
rect 30288 25288 30340 25294
rect 30288 25230 30340 25236
rect 30196 25220 30248 25226
rect 30196 25162 30248 25168
rect 30104 23180 30156 23186
rect 30104 23122 30156 23128
rect 30012 22704 30064 22710
rect 30012 22646 30064 22652
rect 29092 22432 29144 22438
rect 29092 22374 29144 22380
rect 29276 22432 29328 22438
rect 29276 22374 29328 22380
rect 29104 22030 29132 22374
rect 30116 22030 30144 23122
rect 28920 21962 29040 21978
rect 29092 22024 29144 22030
rect 29092 21966 29144 21972
rect 29920 22024 29972 22030
rect 29920 21966 29972 21972
rect 30104 22024 30156 22030
rect 30104 21966 30156 21972
rect 28908 21956 29040 21962
rect 28960 21950 29040 21956
rect 28908 21898 28960 21904
rect 29828 21888 29880 21894
rect 29828 21830 29880 21836
rect 29736 21684 29788 21690
rect 29736 21626 29788 21632
rect 28632 21616 28684 21622
rect 28632 21558 28684 21564
rect 28908 21412 28960 21418
rect 28908 21354 28960 21360
rect 28080 20936 28132 20942
rect 28080 20878 28132 20884
rect 28632 20800 28684 20806
rect 28632 20742 28684 20748
rect 27620 20460 27672 20466
rect 27620 20402 27672 20408
rect 27712 20460 27764 20466
rect 27712 20402 27764 20408
rect 27344 19372 27396 19378
rect 27344 19314 27396 19320
rect 27436 19372 27488 19378
rect 27436 19314 27488 19320
rect 27160 18284 27212 18290
rect 27160 18226 27212 18232
rect 27252 18284 27304 18290
rect 27252 18226 27304 18232
rect 26516 16244 26568 16250
rect 26516 16186 26568 16192
rect 26528 16046 26556 16186
rect 27344 16108 27396 16114
rect 27344 16050 27396 16056
rect 26516 16040 26568 16046
rect 26568 15988 26740 15994
rect 26516 15982 26740 15988
rect 26528 15966 26740 15982
rect 26608 15904 26660 15910
rect 26608 15846 26660 15852
rect 26516 15020 26568 15026
rect 26516 14962 26568 14968
rect 26252 14198 26372 14226
rect 26252 13938 26280 14198
rect 26240 13932 26292 13938
rect 26240 13874 26292 13880
rect 26056 13320 26108 13326
rect 26056 13262 26108 13268
rect 25872 13252 25924 13258
rect 25872 13194 25924 13200
rect 25424 12406 25728 12434
rect 25700 12186 25728 12406
rect 25884 12238 25912 13194
rect 26068 12986 26096 13262
rect 26056 12980 26108 12986
rect 26056 12922 26108 12928
rect 25608 12158 25728 12186
rect 25872 12232 25924 12238
rect 25872 12174 25924 12180
rect 25608 12102 25636 12158
rect 25596 12096 25648 12102
rect 25596 12038 25648 12044
rect 25320 11892 25372 11898
rect 25320 11834 25372 11840
rect 23848 11756 23900 11762
rect 23848 11698 23900 11704
rect 25228 11688 25280 11694
rect 25228 11630 25280 11636
rect 24952 11552 25004 11558
rect 24952 11494 25004 11500
rect 24964 11150 24992 11494
rect 25136 11212 25188 11218
rect 25136 11154 25188 11160
rect 24952 11144 25004 11150
rect 24952 11086 25004 11092
rect 23664 11076 23716 11082
rect 23664 11018 23716 11024
rect 24676 11008 24728 11014
rect 24676 10950 24728 10956
rect 25044 11008 25096 11014
rect 25044 10950 25096 10956
rect 24032 10668 24084 10674
rect 24032 10610 24084 10616
rect 23848 10464 23900 10470
rect 23848 10406 23900 10412
rect 23860 10198 23888 10406
rect 23848 10192 23900 10198
rect 23848 10134 23900 10140
rect 24044 10062 24072 10610
rect 24688 10062 24716 10950
rect 25056 10810 25084 10950
rect 25044 10804 25096 10810
rect 25044 10746 25096 10752
rect 24860 10668 24912 10674
rect 24860 10610 24912 10616
rect 24872 10198 24900 10610
rect 24860 10192 24912 10198
rect 24860 10134 24912 10140
rect 25148 10130 25176 11154
rect 25240 10470 25268 11630
rect 25228 10464 25280 10470
rect 25228 10406 25280 10412
rect 25136 10124 25188 10130
rect 25136 10066 25188 10072
rect 25608 10062 25636 12038
rect 26252 10130 26280 13874
rect 26424 13184 26476 13190
rect 26424 13126 26476 13132
rect 26332 12844 26384 12850
rect 26332 12786 26384 12792
rect 26344 12442 26372 12786
rect 26332 12436 26384 12442
rect 26332 12378 26384 12384
rect 26436 12238 26464 13126
rect 26424 12232 26476 12238
rect 26424 12174 26476 12180
rect 26528 11354 26556 14962
rect 26620 14958 26648 15846
rect 26608 14952 26660 14958
rect 26608 14894 26660 14900
rect 26712 13870 26740 15966
rect 26700 13864 26752 13870
rect 26700 13806 26752 13812
rect 26608 13524 26660 13530
rect 26608 13466 26660 13472
rect 26620 13326 26648 13466
rect 26608 13320 26660 13326
rect 26608 13262 26660 13268
rect 26620 12986 26648 13262
rect 26608 12980 26660 12986
rect 26608 12922 26660 12928
rect 26608 12436 26660 12442
rect 26712 12434 26740 13806
rect 27356 13530 27384 16050
rect 27448 15026 27476 19314
rect 27724 19281 27752 20402
rect 28540 19372 28592 19378
rect 28540 19314 28592 19320
rect 27710 19272 27766 19281
rect 27710 19207 27766 19216
rect 27724 18290 27752 19207
rect 28552 18834 28580 19314
rect 28644 18902 28672 20742
rect 28920 20466 28948 21354
rect 28908 20460 28960 20466
rect 28908 20402 28960 20408
rect 28920 20058 28948 20402
rect 28908 20052 28960 20058
rect 28908 19994 28960 20000
rect 28724 19712 28776 19718
rect 28724 19654 28776 19660
rect 28736 19446 28764 19654
rect 28724 19440 28776 19446
rect 28724 19382 28776 19388
rect 28632 18896 28684 18902
rect 28632 18838 28684 18844
rect 28540 18828 28592 18834
rect 28540 18770 28592 18776
rect 28448 18760 28500 18766
rect 28448 18702 28500 18708
rect 28460 18426 28488 18702
rect 28448 18420 28500 18426
rect 28448 18362 28500 18368
rect 27528 18284 27580 18290
rect 27528 18226 27580 18232
rect 27712 18284 27764 18290
rect 27712 18226 27764 18232
rect 27540 18170 27568 18226
rect 27540 18142 27660 18170
rect 27632 16114 27660 18142
rect 27724 16182 27752 18226
rect 28552 17202 28580 18770
rect 28540 17196 28592 17202
rect 28540 17138 28592 17144
rect 27804 16448 27856 16454
rect 27804 16390 27856 16396
rect 27712 16176 27764 16182
rect 27712 16118 27764 16124
rect 27816 16114 27844 16390
rect 28644 16250 28672 18838
rect 28920 17882 28948 19994
rect 29184 19848 29236 19854
rect 29184 19790 29236 19796
rect 29196 19174 29224 19790
rect 29184 19168 29236 19174
rect 29184 19110 29236 19116
rect 29196 18766 29224 19110
rect 29184 18760 29236 18766
rect 29184 18702 29236 18708
rect 29748 18358 29776 21626
rect 29840 21554 29868 21830
rect 29828 21548 29880 21554
rect 29828 21490 29880 21496
rect 29932 21146 29960 21966
rect 29920 21140 29972 21146
rect 29920 21082 29972 21088
rect 29920 20936 29972 20942
rect 29920 20878 29972 20884
rect 29932 20330 29960 20878
rect 30116 20602 30144 21966
rect 30208 20942 30236 25162
rect 30300 24954 30328 25230
rect 30472 25152 30524 25158
rect 30472 25094 30524 25100
rect 30564 25152 30616 25158
rect 30564 25094 30616 25100
rect 30288 24948 30340 24954
rect 30288 24890 30340 24896
rect 30300 23594 30328 24890
rect 30484 24750 30512 25094
rect 30472 24744 30524 24750
rect 30472 24686 30524 24692
rect 30484 24138 30512 24686
rect 30472 24132 30524 24138
rect 30472 24074 30524 24080
rect 30484 23730 30512 24074
rect 30380 23724 30432 23730
rect 30380 23666 30432 23672
rect 30472 23724 30524 23730
rect 30472 23666 30524 23672
rect 30288 23588 30340 23594
rect 30288 23530 30340 23536
rect 30288 23112 30340 23118
rect 30288 23054 30340 23060
rect 30300 22030 30328 23054
rect 30392 23050 30420 23666
rect 30472 23112 30524 23118
rect 30472 23054 30524 23060
rect 30380 23044 30432 23050
rect 30380 22986 30432 22992
rect 30288 22024 30340 22030
rect 30288 21966 30340 21972
rect 30300 21690 30328 21966
rect 30288 21684 30340 21690
rect 30288 21626 30340 21632
rect 30392 20942 30420 22986
rect 30484 21078 30512 23054
rect 30576 22982 30604 25094
rect 30748 24812 30800 24818
rect 30748 24754 30800 24760
rect 31024 24812 31076 24818
rect 31024 24754 31076 24760
rect 30760 23798 30788 24754
rect 30748 23792 30800 23798
rect 30748 23734 30800 23740
rect 30564 22976 30616 22982
rect 30564 22918 30616 22924
rect 30840 22636 30892 22642
rect 30840 22578 30892 22584
rect 30852 21962 30880 22578
rect 31036 22030 31064 24754
rect 31128 24274 31156 25774
rect 31220 25498 31248 25842
rect 31576 25832 31628 25838
rect 31576 25774 31628 25780
rect 31208 25492 31260 25498
rect 31208 25434 31260 25440
rect 31588 25294 31616 25774
rect 31576 25288 31628 25294
rect 31576 25230 31628 25236
rect 31208 24812 31260 24818
rect 31208 24754 31260 24760
rect 31484 24812 31536 24818
rect 31484 24754 31536 24760
rect 31220 24342 31248 24754
rect 31208 24336 31260 24342
rect 31208 24278 31260 24284
rect 31116 24268 31168 24274
rect 31116 24210 31168 24216
rect 31128 23662 31156 24210
rect 31496 24206 31524 24754
rect 31484 24200 31536 24206
rect 31484 24142 31536 24148
rect 31116 23656 31168 23662
rect 31116 23598 31168 23604
rect 31588 23186 31616 25230
rect 31680 23526 31708 25894
rect 32324 25498 32352 26250
rect 32600 25906 32628 33782
rect 32692 33538 32720 34954
rect 33520 34678 33548 35090
rect 34716 35018 34744 35566
rect 34704 35012 34756 35018
rect 34704 34954 34756 34960
rect 34428 34944 34480 34950
rect 34428 34886 34480 34892
rect 33508 34672 33560 34678
rect 33508 34614 33560 34620
rect 33796 34610 34008 34626
rect 34440 34610 34468 34886
rect 33416 34604 33468 34610
rect 33416 34546 33468 34552
rect 33784 34604 34020 34610
rect 33836 34598 33968 34604
rect 33784 34546 33836 34552
rect 33968 34546 34020 34552
rect 34428 34604 34480 34610
rect 34428 34546 34480 34552
rect 32772 33924 32824 33930
rect 32772 33866 32824 33872
rect 32784 33658 32812 33866
rect 33428 33862 33456 34546
rect 34716 34474 34744 34954
rect 34808 34678 34836 35634
rect 35440 35488 35492 35494
rect 35440 35430 35492 35436
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 35348 35148 35400 35154
rect 35348 35090 35400 35096
rect 34796 34672 34848 34678
rect 34796 34614 34848 34620
rect 34704 34468 34756 34474
rect 34704 34410 34756 34416
rect 34808 33998 34836 34614
rect 35360 34542 35388 35090
rect 35348 34536 35400 34542
rect 35348 34478 35400 34484
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34796 33992 34848 33998
rect 34796 33934 34848 33940
rect 33416 33856 33468 33862
rect 33416 33798 33468 33804
rect 32772 33652 32824 33658
rect 32772 33594 32824 33600
rect 32692 33510 32812 33538
rect 32680 30252 32732 30258
rect 32680 30194 32732 30200
rect 32692 29170 32720 30194
rect 32784 30190 32812 33510
rect 32956 33516 33008 33522
rect 32956 33458 33008 33464
rect 32968 33114 32996 33458
rect 32956 33108 33008 33114
rect 32956 33050 33008 33056
rect 33428 32910 33456 33798
rect 34612 33380 34664 33386
rect 34612 33322 34664 33328
rect 33416 32904 33468 32910
rect 33416 32846 33468 32852
rect 33140 32836 33192 32842
rect 33140 32778 33192 32784
rect 33048 32768 33100 32774
rect 33048 32710 33100 32716
rect 32864 32496 32916 32502
rect 32864 32438 32916 32444
rect 32772 30184 32824 30190
rect 32772 30126 32824 30132
rect 32876 29782 32904 32438
rect 33060 32434 33088 32710
rect 33152 32570 33180 32778
rect 33600 32768 33652 32774
rect 33600 32710 33652 32716
rect 33612 32570 33640 32710
rect 34624 32570 34652 33322
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 35256 32972 35308 32978
rect 35256 32914 35308 32920
rect 33140 32564 33192 32570
rect 33140 32506 33192 32512
rect 33600 32564 33652 32570
rect 33600 32506 33652 32512
rect 34612 32564 34664 32570
rect 34612 32506 34664 32512
rect 35268 32434 35296 32914
rect 33048 32428 33100 32434
rect 33048 32370 33100 32376
rect 34796 32428 34848 32434
rect 34796 32370 34848 32376
rect 35256 32428 35308 32434
rect 35256 32370 35308 32376
rect 34704 32360 34756 32366
rect 34704 32302 34756 32308
rect 34716 31686 34744 32302
rect 34704 31680 34756 31686
rect 34704 31622 34756 31628
rect 33968 31340 34020 31346
rect 33968 31282 34020 31288
rect 33048 31136 33100 31142
rect 33048 31078 33100 31084
rect 32864 29776 32916 29782
rect 32916 29724 32996 29730
rect 32864 29718 32996 29724
rect 32876 29702 32996 29718
rect 32968 29170 32996 29702
rect 32680 29164 32732 29170
rect 32680 29106 32732 29112
rect 32956 29164 33008 29170
rect 32956 29106 33008 29112
rect 33060 28558 33088 31078
rect 33232 30116 33284 30122
rect 33232 30058 33284 30064
rect 33244 29102 33272 30058
rect 33980 29782 34008 31282
rect 34716 30802 34744 31622
rect 34808 31482 34836 32370
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35360 31890 35388 34478
rect 35452 34134 35480 35430
rect 35808 35080 35860 35086
rect 35808 35022 35860 35028
rect 35992 35080 36044 35086
rect 35992 35022 36044 35028
rect 37004 35080 37056 35086
rect 37004 35022 37056 35028
rect 38660 35080 38712 35086
rect 38660 35022 38712 35028
rect 39028 35080 39080 35086
rect 39028 35022 39080 35028
rect 39212 35080 39264 35086
rect 39212 35022 39264 35028
rect 35624 35012 35676 35018
rect 35624 34954 35676 34960
rect 35532 34944 35584 34950
rect 35532 34886 35584 34892
rect 35544 34134 35572 34886
rect 35636 34610 35664 34954
rect 35820 34678 35848 35022
rect 36004 34746 36032 35022
rect 36820 35012 36872 35018
rect 36820 34954 36872 34960
rect 36912 35012 36964 35018
rect 36912 34954 36964 34960
rect 36268 34944 36320 34950
rect 36268 34886 36320 34892
rect 35992 34740 36044 34746
rect 35992 34682 36044 34688
rect 35808 34672 35860 34678
rect 35808 34614 35860 34620
rect 35624 34604 35676 34610
rect 35624 34546 35676 34552
rect 35440 34128 35492 34134
rect 35440 34070 35492 34076
rect 35532 34128 35584 34134
rect 35532 34070 35584 34076
rect 35452 33590 35480 34070
rect 35440 33584 35492 33590
rect 35440 33526 35492 33532
rect 35532 32768 35584 32774
rect 35532 32710 35584 32716
rect 35440 32224 35492 32230
rect 35440 32166 35492 32172
rect 35348 31884 35400 31890
rect 35348 31826 35400 31832
rect 34796 31476 34848 31482
rect 34796 31418 34848 31424
rect 34704 30796 34756 30802
rect 34704 30738 34756 30744
rect 34334 30288 34390 30297
rect 34808 30258 34836 31418
rect 35360 31414 35388 31826
rect 35452 31822 35480 32166
rect 35440 31816 35492 31822
rect 35440 31758 35492 31764
rect 35348 31408 35400 31414
rect 35348 31350 35400 31356
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34334 30223 34336 30232
rect 34388 30223 34390 30232
rect 34612 30252 34664 30258
rect 34336 30194 34388 30200
rect 34612 30194 34664 30200
rect 34796 30252 34848 30258
rect 34796 30194 34848 30200
rect 34624 30122 34652 30194
rect 34612 30116 34664 30122
rect 34612 30058 34664 30064
rect 34060 30048 34112 30054
rect 34060 29990 34112 29996
rect 34704 30048 34756 30054
rect 34704 29990 34756 29996
rect 33968 29776 34020 29782
rect 33968 29718 34020 29724
rect 34072 29646 34100 29990
rect 34060 29640 34112 29646
rect 34060 29582 34112 29588
rect 34336 29640 34388 29646
rect 34336 29582 34388 29588
rect 33508 29572 33560 29578
rect 33508 29514 33560 29520
rect 33324 29504 33376 29510
rect 33324 29446 33376 29452
rect 33416 29504 33468 29510
rect 33416 29446 33468 29452
rect 33336 29306 33364 29446
rect 33324 29300 33376 29306
rect 33324 29242 33376 29248
rect 33232 29096 33284 29102
rect 33232 29038 33284 29044
rect 33336 28642 33364 29242
rect 33428 29102 33456 29446
rect 33520 29170 33548 29514
rect 34348 29322 34376 29582
rect 34164 29306 34376 29322
rect 34152 29300 34376 29306
rect 34204 29294 34376 29300
rect 34152 29242 34204 29248
rect 33508 29164 33560 29170
rect 33508 29106 33560 29112
rect 33416 29096 33468 29102
rect 33416 29038 33468 29044
rect 33428 28762 33456 29038
rect 33416 28756 33468 28762
rect 33416 28698 33468 28704
rect 33336 28614 33548 28642
rect 33048 28552 33100 28558
rect 33048 28494 33100 28500
rect 33232 28552 33284 28558
rect 33232 28494 33284 28500
rect 32864 27464 32916 27470
rect 32864 27406 32916 27412
rect 33140 27464 33192 27470
rect 33140 27406 33192 27412
rect 32680 27328 32732 27334
rect 32680 27270 32732 27276
rect 32692 27062 32720 27270
rect 32680 27056 32732 27062
rect 32680 26998 32732 27004
rect 32876 26042 32904 27406
rect 33152 27130 33180 27406
rect 33140 27124 33192 27130
rect 33140 27066 33192 27072
rect 32864 26036 32916 26042
rect 32864 25978 32916 25984
rect 32588 25900 32640 25906
rect 32588 25842 32640 25848
rect 32864 25900 32916 25906
rect 32864 25842 32916 25848
rect 33140 25900 33192 25906
rect 33140 25842 33192 25848
rect 32600 25498 32628 25842
rect 32680 25832 32732 25838
rect 32680 25774 32732 25780
rect 32312 25492 32364 25498
rect 32312 25434 32364 25440
rect 32588 25492 32640 25498
rect 32588 25434 32640 25440
rect 31760 24608 31812 24614
rect 31760 24550 31812 24556
rect 31852 24608 31904 24614
rect 31852 24550 31904 24556
rect 31772 24342 31800 24550
rect 31760 24336 31812 24342
rect 31760 24278 31812 24284
rect 31864 24138 31892 24550
rect 32496 24404 32548 24410
rect 32496 24346 32548 24352
rect 31852 24132 31904 24138
rect 31852 24074 31904 24080
rect 31668 23520 31720 23526
rect 31668 23462 31720 23468
rect 31576 23180 31628 23186
rect 31576 23122 31628 23128
rect 31680 23118 31708 23462
rect 31668 23112 31720 23118
rect 31668 23054 31720 23060
rect 31300 22976 31352 22982
rect 31300 22918 31352 22924
rect 31312 22642 31340 22918
rect 31300 22636 31352 22642
rect 31300 22578 31352 22584
rect 31208 22432 31260 22438
rect 31208 22374 31260 22380
rect 31220 22030 31248 22374
rect 31024 22024 31076 22030
rect 31024 21966 31076 21972
rect 31208 22024 31260 22030
rect 31208 21966 31260 21972
rect 30840 21956 30892 21962
rect 30840 21898 30892 21904
rect 30656 21412 30708 21418
rect 30656 21354 30708 21360
rect 30472 21072 30524 21078
rect 30472 21014 30524 21020
rect 30196 20936 30248 20942
rect 30380 20936 30432 20942
rect 30196 20878 30248 20884
rect 30300 20884 30380 20890
rect 30300 20878 30432 20884
rect 30300 20862 30420 20878
rect 30104 20596 30156 20602
rect 30104 20538 30156 20544
rect 29920 20324 29972 20330
rect 29920 20266 29972 20272
rect 29932 19854 29960 20266
rect 29920 19848 29972 19854
rect 29920 19790 29972 19796
rect 30196 19848 30248 19854
rect 30300 19836 30328 20862
rect 30248 19808 30328 19836
rect 30380 19848 30432 19854
rect 30196 19790 30248 19796
rect 30380 19790 30432 19796
rect 29828 18760 29880 18766
rect 29828 18702 29880 18708
rect 29736 18352 29788 18358
rect 29736 18294 29788 18300
rect 29840 18290 29868 18702
rect 29828 18284 29880 18290
rect 29828 18226 29880 18232
rect 28908 17876 28960 17882
rect 28908 17818 28960 17824
rect 28632 16244 28684 16250
rect 28632 16186 28684 16192
rect 28724 16176 28776 16182
rect 28724 16118 28776 16124
rect 27620 16108 27672 16114
rect 27620 16050 27672 16056
rect 27804 16108 27856 16114
rect 27804 16050 27856 16056
rect 28632 16108 28684 16114
rect 28632 16050 28684 16056
rect 27436 15020 27488 15026
rect 27436 14962 27488 14968
rect 27344 13524 27396 13530
rect 27344 13466 27396 13472
rect 27632 13394 27660 16050
rect 27816 15706 27844 16050
rect 28644 15706 28672 16050
rect 27804 15700 27856 15706
rect 27804 15642 27856 15648
rect 28632 15700 28684 15706
rect 28632 15642 28684 15648
rect 28736 15502 28764 16118
rect 28920 15706 28948 17818
rect 29460 17740 29512 17746
rect 29460 17682 29512 17688
rect 29000 17536 29052 17542
rect 29000 17478 29052 17484
rect 29184 17536 29236 17542
rect 29184 17478 29236 17484
rect 28908 15700 28960 15706
rect 28908 15642 28960 15648
rect 29012 15570 29040 17478
rect 29196 17270 29224 17478
rect 29184 17264 29236 17270
rect 29184 17206 29236 17212
rect 29472 16590 29500 17682
rect 29460 16584 29512 16590
rect 29460 16526 29512 16532
rect 29472 15910 29500 16526
rect 29460 15904 29512 15910
rect 29460 15846 29512 15852
rect 29000 15564 29052 15570
rect 29000 15506 29052 15512
rect 28724 15496 28776 15502
rect 28724 15438 28776 15444
rect 28736 15026 28764 15438
rect 28724 15020 28776 15026
rect 28724 14962 28776 14968
rect 28736 14414 28764 14962
rect 28724 14408 28776 14414
rect 28724 14350 28776 14356
rect 28736 13394 28764 14350
rect 27620 13388 27672 13394
rect 27620 13330 27672 13336
rect 28724 13388 28776 13394
rect 28724 13330 28776 13336
rect 28356 13320 28408 13326
rect 28356 13262 28408 13268
rect 28632 13320 28684 13326
rect 28632 13262 28684 13268
rect 27988 13184 28040 13190
rect 27988 13126 28040 13132
rect 28000 12850 28028 13126
rect 27988 12844 28040 12850
rect 27988 12786 28040 12792
rect 28368 12442 28396 13262
rect 28540 13252 28592 13258
rect 28540 13194 28592 13200
rect 26660 12406 26740 12434
rect 28356 12436 28408 12442
rect 26608 12378 26660 12384
rect 28356 12378 28408 12384
rect 26608 12300 26660 12306
rect 26608 12242 26660 12248
rect 26516 11348 26568 11354
rect 26516 11290 26568 11296
rect 26620 11218 26648 12242
rect 28552 11762 28580 13194
rect 28540 11756 28592 11762
rect 28540 11698 28592 11704
rect 26608 11212 26660 11218
rect 26608 11154 26660 11160
rect 26700 11144 26752 11150
rect 26700 11086 26752 11092
rect 26712 10266 26740 11086
rect 28264 11076 28316 11082
rect 28264 11018 28316 11024
rect 28276 10674 28304 11018
rect 28264 10668 28316 10674
rect 28264 10610 28316 10616
rect 26884 10464 26936 10470
rect 26884 10406 26936 10412
rect 26700 10260 26752 10266
rect 26700 10202 26752 10208
rect 26240 10124 26292 10130
rect 26240 10066 26292 10072
rect 26896 10062 26924 10406
rect 24032 10056 24084 10062
rect 24032 9998 24084 10004
rect 24676 10056 24728 10062
rect 24676 9998 24728 10004
rect 25320 10056 25372 10062
rect 25320 9998 25372 10004
rect 25596 10056 25648 10062
rect 25596 9998 25648 10004
rect 26884 10056 26936 10062
rect 26884 9998 26936 10004
rect 24044 9722 24072 9998
rect 25332 9722 25360 9998
rect 24032 9716 24084 9722
rect 24032 9658 24084 9664
rect 25320 9716 25372 9722
rect 25320 9658 25372 9664
rect 28552 8430 28580 11698
rect 28644 11150 28672 13262
rect 28736 12918 28764 13330
rect 28724 12912 28776 12918
rect 28724 12854 28776 12860
rect 29092 12640 29144 12646
rect 29092 12582 29144 12588
rect 29104 12374 29132 12582
rect 29092 12368 29144 12374
rect 29092 12310 29144 12316
rect 29104 12238 29132 12310
rect 29092 12232 29144 12238
rect 29092 12174 29144 12180
rect 29000 11892 29052 11898
rect 29000 11834 29052 11840
rect 29012 11150 29040 11834
rect 28632 11144 28684 11150
rect 28632 11086 28684 11092
rect 29000 11144 29052 11150
rect 29000 11086 29052 11092
rect 29092 11144 29144 11150
rect 29092 11086 29144 11092
rect 29104 10674 29132 11086
rect 29092 10668 29144 10674
rect 29092 10610 29144 10616
rect 28540 8424 28592 8430
rect 28540 8366 28592 8372
rect 29472 6914 29500 15846
rect 29644 13252 29696 13258
rect 29644 13194 29696 13200
rect 29656 11694 29684 13194
rect 29840 13138 29868 18226
rect 29932 17678 29960 19790
rect 30208 17678 30236 19790
rect 30392 19514 30420 19790
rect 30380 19508 30432 19514
rect 30380 19450 30432 19456
rect 30484 19258 30512 21014
rect 30668 20942 30696 21354
rect 30748 21344 30800 21350
rect 30748 21286 30800 21292
rect 30656 20936 30708 20942
rect 30656 20878 30708 20884
rect 30656 19372 30708 19378
rect 30656 19314 30708 19320
rect 30484 19230 30604 19258
rect 30472 19168 30524 19174
rect 30472 19110 30524 19116
rect 30484 18698 30512 19110
rect 30472 18692 30524 18698
rect 30472 18634 30524 18640
rect 30576 18290 30604 19230
rect 30668 18426 30696 19314
rect 30656 18420 30708 18426
rect 30656 18362 30708 18368
rect 30760 18290 30788 21286
rect 30852 19378 30880 21898
rect 30932 21888 30984 21894
rect 30932 21830 30984 21836
rect 30944 21622 30972 21830
rect 30932 21616 30984 21622
rect 30932 21558 30984 21564
rect 31036 21350 31064 21966
rect 31668 21888 31720 21894
rect 31668 21830 31720 21836
rect 31024 21344 31076 21350
rect 31024 21286 31076 21292
rect 31680 19922 31708 21830
rect 31668 19916 31720 19922
rect 31668 19858 31720 19864
rect 30840 19372 30892 19378
rect 30840 19314 30892 19320
rect 31300 19372 31352 19378
rect 31300 19314 31352 19320
rect 30564 18284 30616 18290
rect 30564 18226 30616 18232
rect 30748 18284 30800 18290
rect 30748 18226 30800 18232
rect 29920 17672 29972 17678
rect 29920 17614 29972 17620
rect 30196 17672 30248 17678
rect 30196 17614 30248 17620
rect 30104 17536 30156 17542
rect 30104 17478 30156 17484
rect 30116 17338 30144 17478
rect 30104 17332 30156 17338
rect 30104 17274 30156 17280
rect 30208 17218 30236 17614
rect 30288 17604 30340 17610
rect 30288 17546 30340 17552
rect 30116 17190 30236 17218
rect 30012 15700 30064 15706
rect 30012 15642 30064 15648
rect 30024 14550 30052 15642
rect 30116 15570 30144 17190
rect 30104 15564 30156 15570
rect 30104 15506 30156 15512
rect 30012 14544 30064 14550
rect 30012 14486 30064 14492
rect 29920 14272 29972 14278
rect 29920 14214 29972 14220
rect 29932 13326 29960 14214
rect 30024 13938 30052 14486
rect 30116 14414 30144 15506
rect 30300 15502 30328 17546
rect 30576 16522 30604 18226
rect 30760 16590 30788 18226
rect 31312 17678 31340 19314
rect 31576 19304 31628 19310
rect 31576 19246 31628 19252
rect 31588 18970 31616 19246
rect 31576 18964 31628 18970
rect 31576 18906 31628 18912
rect 31680 18766 31708 19858
rect 31864 19378 31892 24074
rect 32508 23866 32536 24346
rect 32496 23860 32548 23866
rect 32496 23802 32548 23808
rect 32600 23322 32628 25434
rect 32692 25294 32720 25774
rect 32680 25288 32732 25294
rect 32680 25230 32732 25236
rect 32588 23316 32640 23322
rect 32588 23258 32640 23264
rect 32220 23248 32272 23254
rect 32220 23190 32272 23196
rect 32232 22234 32260 23190
rect 32220 22228 32272 22234
rect 32220 22170 32272 22176
rect 32496 21616 32548 21622
rect 32496 21558 32548 21564
rect 32312 19780 32364 19786
rect 32312 19722 32364 19728
rect 32324 19514 32352 19722
rect 32312 19508 32364 19514
rect 32312 19450 32364 19456
rect 32404 19508 32456 19514
rect 32404 19450 32456 19456
rect 32416 19378 32444 19450
rect 31852 19372 31904 19378
rect 31852 19314 31904 19320
rect 32404 19372 32456 19378
rect 32404 19314 32456 19320
rect 31668 18760 31720 18766
rect 31668 18702 31720 18708
rect 31760 18692 31812 18698
rect 31760 18634 31812 18640
rect 31116 17672 31168 17678
rect 31116 17614 31168 17620
rect 31300 17672 31352 17678
rect 31300 17614 31352 17620
rect 31576 17672 31628 17678
rect 31576 17614 31628 17620
rect 31128 16794 31156 17614
rect 31116 16788 31168 16794
rect 31116 16730 31168 16736
rect 30748 16584 30800 16590
rect 30748 16526 30800 16532
rect 30564 16516 30616 16522
rect 30564 16458 30616 16464
rect 30576 15722 30604 16458
rect 30576 15694 30696 15722
rect 30564 15632 30616 15638
rect 30564 15574 30616 15580
rect 30288 15496 30340 15502
rect 30288 15438 30340 15444
rect 30300 14414 30328 15438
rect 30472 15428 30524 15434
rect 30472 15370 30524 15376
rect 30484 15178 30512 15370
rect 30392 15162 30512 15178
rect 30392 15156 30524 15162
rect 30392 15150 30472 15156
rect 30104 14408 30156 14414
rect 30104 14350 30156 14356
rect 30288 14408 30340 14414
rect 30288 14350 30340 14356
rect 30012 13932 30064 13938
rect 30012 13874 30064 13880
rect 30024 13530 30052 13874
rect 30012 13524 30064 13530
rect 30012 13466 30064 13472
rect 30012 13388 30064 13394
rect 30012 13330 30064 13336
rect 29920 13320 29972 13326
rect 29920 13262 29972 13268
rect 29840 13110 29960 13138
rect 29828 12844 29880 12850
rect 29828 12786 29880 12792
rect 29644 11688 29696 11694
rect 29644 11630 29696 11636
rect 29656 11218 29684 11630
rect 29644 11212 29696 11218
rect 29644 11154 29696 11160
rect 29840 11150 29868 12786
rect 29828 11144 29880 11150
rect 29828 11086 29880 11092
rect 29552 11076 29604 11082
rect 29552 11018 29604 11024
rect 29564 10810 29592 11018
rect 29736 11008 29788 11014
rect 29736 10950 29788 10956
rect 29552 10804 29604 10810
rect 29552 10746 29604 10752
rect 29748 10674 29776 10950
rect 29736 10668 29788 10674
rect 29736 10610 29788 10616
rect 29932 6914 29960 13110
rect 30024 12850 30052 13330
rect 30012 12844 30064 12850
rect 30012 12786 30064 12792
rect 30116 12170 30144 14350
rect 30196 13932 30248 13938
rect 30196 13874 30248 13880
rect 30208 12442 30236 13874
rect 30196 12436 30248 12442
rect 30196 12378 30248 12384
rect 30300 12238 30328 14350
rect 30392 14346 30420 15150
rect 30472 15098 30524 15104
rect 30576 15026 30604 15574
rect 30668 15094 30696 15694
rect 30656 15088 30708 15094
rect 30656 15030 30708 15036
rect 30760 15042 30788 16526
rect 30840 15904 30892 15910
rect 30840 15846 30892 15852
rect 30852 15502 30880 15846
rect 31588 15502 31616 17614
rect 31772 16522 31800 18634
rect 32508 17338 32536 21558
rect 32692 21010 32720 25230
rect 32772 24948 32824 24954
rect 32772 24890 32824 24896
rect 32680 21004 32732 21010
rect 32680 20946 32732 20952
rect 32496 17332 32548 17338
rect 32496 17274 32548 17280
rect 32784 17270 32812 24890
rect 32876 24818 32904 25842
rect 33152 24834 33180 25842
rect 32864 24812 32916 24818
rect 32864 24754 32916 24760
rect 33060 24806 33180 24834
rect 33060 23866 33088 24806
rect 33244 24614 33272 28494
rect 33324 28484 33376 28490
rect 33324 28426 33376 28432
rect 33416 28484 33468 28490
rect 33416 28426 33468 28432
rect 33336 27878 33364 28426
rect 33428 28218 33456 28426
rect 33416 28212 33468 28218
rect 33416 28154 33468 28160
rect 33324 27872 33376 27878
rect 33324 27814 33376 27820
rect 33232 24608 33284 24614
rect 33232 24550 33284 24556
rect 33140 24132 33192 24138
rect 33140 24074 33192 24080
rect 33048 23860 33100 23866
rect 33048 23802 33100 23808
rect 32956 23044 33008 23050
rect 32956 22986 33008 22992
rect 32968 22710 32996 22986
rect 32956 22704 33008 22710
rect 32956 22646 33008 22652
rect 32864 19712 32916 19718
rect 32864 19654 32916 19660
rect 32876 19378 32904 19654
rect 32864 19372 32916 19378
rect 32864 19314 32916 19320
rect 33060 18698 33088 23802
rect 33152 23322 33180 24074
rect 33232 23520 33284 23526
rect 33232 23462 33284 23468
rect 33140 23316 33192 23322
rect 33140 23258 33192 23264
rect 33244 23118 33272 23462
rect 33232 23112 33284 23118
rect 33232 23054 33284 23060
rect 33336 22094 33364 27814
rect 33416 27056 33468 27062
rect 33416 26998 33468 27004
rect 33428 26586 33456 26998
rect 33416 26580 33468 26586
rect 33416 26522 33468 26528
rect 33520 24970 33548 28614
rect 34716 28082 34744 29990
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35360 29714 35388 31350
rect 35544 31346 35572 32710
rect 35636 32366 35664 34546
rect 36280 34202 36308 34886
rect 36832 34610 36860 34954
rect 36924 34746 36952 34954
rect 37016 34746 37044 35022
rect 37648 34944 37700 34950
rect 37648 34886 37700 34892
rect 36912 34740 36964 34746
rect 36912 34682 36964 34688
rect 37004 34740 37056 34746
rect 37004 34682 37056 34688
rect 36820 34604 36872 34610
rect 36820 34546 36872 34552
rect 36268 34196 36320 34202
rect 36268 34138 36320 34144
rect 36280 34082 36308 34138
rect 36188 34054 36308 34082
rect 37016 34066 37044 34682
rect 37660 34610 37688 34886
rect 37648 34604 37700 34610
rect 37648 34546 37700 34552
rect 37556 34536 37608 34542
rect 37556 34478 37608 34484
rect 38016 34536 38068 34542
rect 38016 34478 38068 34484
rect 37568 34202 37596 34478
rect 37556 34196 37608 34202
rect 37556 34138 37608 34144
rect 37004 34060 37056 34066
rect 36188 33930 36216 34054
rect 37004 34002 37056 34008
rect 36268 33992 36320 33998
rect 36268 33934 36320 33940
rect 36176 33924 36228 33930
rect 36176 33866 36228 33872
rect 36188 32910 36216 33866
rect 36280 33266 36308 33934
rect 37372 33924 37424 33930
rect 37372 33866 37424 33872
rect 36544 33856 36596 33862
rect 36544 33798 36596 33804
rect 36556 33454 36584 33798
rect 36544 33448 36596 33454
rect 36544 33390 36596 33396
rect 36280 33238 36400 33266
rect 36176 32904 36228 32910
rect 36176 32846 36228 32852
rect 36188 32434 36216 32846
rect 36372 32842 36400 33238
rect 36360 32836 36412 32842
rect 36360 32778 36412 32784
rect 36372 32502 36400 32778
rect 36360 32496 36412 32502
rect 36360 32438 36412 32444
rect 35992 32428 36044 32434
rect 35992 32370 36044 32376
rect 36176 32428 36228 32434
rect 36176 32370 36228 32376
rect 35624 32360 35676 32366
rect 35624 32302 35676 32308
rect 35636 32026 35664 32302
rect 35624 32020 35676 32026
rect 35624 31962 35676 31968
rect 35808 31748 35860 31754
rect 35808 31690 35860 31696
rect 35820 31346 35848 31690
rect 36004 31482 36032 32370
rect 36912 32292 36964 32298
rect 36912 32234 36964 32240
rect 36176 32224 36228 32230
rect 36176 32166 36228 32172
rect 36084 31680 36136 31686
rect 36084 31622 36136 31628
rect 35992 31476 36044 31482
rect 35992 31418 36044 31424
rect 35532 31340 35584 31346
rect 35532 31282 35584 31288
rect 35808 31340 35860 31346
rect 35808 31282 35860 31288
rect 36096 30666 36124 31622
rect 36188 31414 36216 32166
rect 36176 31408 36228 31414
rect 36176 31350 36228 31356
rect 36924 30734 36952 32234
rect 36912 30728 36964 30734
rect 36912 30670 36964 30676
rect 37188 30728 37240 30734
rect 37188 30670 37240 30676
rect 36084 30660 36136 30666
rect 36084 30602 36136 30608
rect 36268 30660 36320 30666
rect 36268 30602 36320 30608
rect 35438 30288 35494 30297
rect 35438 30223 35440 30232
rect 35492 30223 35494 30232
rect 35440 30194 35492 30200
rect 35348 29708 35400 29714
rect 35348 29650 35400 29656
rect 34796 29572 34848 29578
rect 34796 29514 34848 29520
rect 34704 28076 34756 28082
rect 34704 28018 34756 28024
rect 34520 28008 34572 28014
rect 34520 27950 34572 27956
rect 34152 27056 34204 27062
rect 34152 26998 34204 27004
rect 33692 25696 33744 25702
rect 33692 25638 33744 25644
rect 33704 25294 33732 25638
rect 33784 25492 33836 25498
rect 33784 25434 33836 25440
rect 33692 25288 33744 25294
rect 33692 25230 33744 25236
rect 33428 24942 33548 24970
rect 33428 22506 33456 24942
rect 33508 24880 33560 24886
rect 33508 24822 33560 24828
rect 33520 23730 33548 24822
rect 33600 24812 33652 24818
rect 33600 24754 33652 24760
rect 33508 23724 33560 23730
rect 33508 23666 33560 23672
rect 33612 23186 33640 24754
rect 33704 23662 33732 25230
rect 33796 24818 33824 25434
rect 34164 25294 34192 26998
rect 34244 26376 34296 26382
rect 34244 26318 34296 26324
rect 34256 25838 34284 26318
rect 34244 25832 34296 25838
rect 34244 25774 34296 25780
rect 33968 25288 34020 25294
rect 33968 25230 34020 25236
rect 34152 25288 34204 25294
rect 34152 25230 34204 25236
rect 33980 24886 34008 25230
rect 33968 24880 34020 24886
rect 33968 24822 34020 24828
rect 33784 24812 33836 24818
rect 33784 24754 33836 24760
rect 33796 24290 33824 24754
rect 34152 24744 34204 24750
rect 34152 24686 34204 24692
rect 34164 24614 34192 24686
rect 34152 24608 34204 24614
rect 34152 24550 34204 24556
rect 33796 24274 34008 24290
rect 33796 24268 34020 24274
rect 33796 24262 33968 24268
rect 33968 24210 34020 24216
rect 34256 24206 34284 25774
rect 34532 24410 34560 27950
rect 34808 25906 34836 29514
rect 35360 29238 35388 29650
rect 35348 29232 35400 29238
rect 35348 29174 35400 29180
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 35360 28762 35388 29174
rect 35452 29170 35480 30194
rect 35440 29164 35492 29170
rect 35440 29106 35492 29112
rect 36280 29102 36308 30602
rect 36452 30252 36504 30258
rect 36452 30194 36504 30200
rect 36464 29646 36492 30194
rect 36636 30048 36688 30054
rect 36636 29990 36688 29996
rect 36452 29640 36504 29646
rect 36452 29582 36504 29588
rect 36268 29096 36320 29102
rect 36268 29038 36320 29044
rect 36464 28762 36492 29582
rect 36648 29170 36676 29990
rect 36636 29164 36688 29170
rect 36636 29106 36688 29112
rect 35348 28756 35400 28762
rect 35348 28698 35400 28704
rect 36452 28756 36504 28762
rect 36452 28698 36504 28704
rect 37200 28694 37228 30670
rect 37384 29714 37412 33866
rect 37740 33856 37792 33862
rect 37740 33798 37792 33804
rect 37556 31816 37608 31822
rect 37556 31758 37608 31764
rect 37648 31816 37700 31822
rect 37648 31758 37700 31764
rect 37464 31136 37516 31142
rect 37464 31078 37516 31084
rect 37476 30734 37504 31078
rect 37568 30938 37596 31758
rect 37660 31278 37688 31758
rect 37752 31278 37780 33798
rect 37832 32768 37884 32774
rect 37832 32710 37884 32716
rect 37844 31346 37872 32710
rect 37924 32564 37976 32570
rect 37924 32506 37976 32512
rect 37936 31890 37964 32506
rect 38028 32434 38056 34478
rect 38016 32428 38068 32434
rect 38016 32370 38068 32376
rect 38292 32428 38344 32434
rect 38292 32370 38344 32376
rect 38028 31890 38056 32370
rect 38304 32026 38332 32370
rect 38292 32020 38344 32026
rect 38292 31962 38344 31968
rect 37924 31884 37976 31890
rect 37924 31826 37976 31832
rect 38016 31884 38068 31890
rect 38016 31826 38068 31832
rect 38016 31748 38068 31754
rect 38016 31690 38068 31696
rect 37924 31680 37976 31686
rect 37924 31622 37976 31628
rect 37936 31414 37964 31622
rect 37924 31408 37976 31414
rect 37924 31350 37976 31356
rect 37832 31340 37884 31346
rect 37832 31282 37884 31288
rect 37648 31272 37700 31278
rect 37648 31214 37700 31220
rect 37740 31272 37792 31278
rect 37740 31214 37792 31220
rect 37556 30932 37608 30938
rect 37556 30874 37608 30880
rect 37464 30728 37516 30734
rect 37464 30670 37516 30676
rect 37372 29708 37424 29714
rect 37372 29650 37424 29656
rect 37280 29232 37332 29238
rect 37280 29174 37332 29180
rect 37188 28688 37240 28694
rect 37188 28630 37240 28636
rect 34980 28484 35032 28490
rect 34980 28426 35032 28432
rect 34992 28218 35020 28426
rect 34980 28212 35032 28218
rect 34980 28154 35032 28160
rect 37096 27940 37148 27946
rect 37096 27882 37148 27888
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 36360 27464 36412 27470
rect 36360 27406 36412 27412
rect 36544 27464 36596 27470
rect 36544 27406 36596 27412
rect 36372 27062 36400 27406
rect 36556 27130 36584 27406
rect 36544 27124 36596 27130
rect 36544 27066 36596 27072
rect 36360 27056 36412 27062
rect 36360 26998 36412 27004
rect 35440 26988 35492 26994
rect 35440 26930 35492 26936
rect 35348 26784 35400 26790
rect 35348 26726 35400 26732
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35360 26314 35388 26726
rect 35348 26308 35400 26314
rect 35348 26250 35400 26256
rect 35452 26042 35480 26930
rect 36268 26920 36320 26926
rect 36268 26862 36320 26868
rect 35808 26784 35860 26790
rect 35808 26726 35860 26732
rect 35820 26042 35848 26726
rect 36280 26586 36308 26862
rect 36268 26580 36320 26586
rect 36268 26522 36320 26528
rect 36372 26246 36400 26998
rect 36556 26994 36584 27066
rect 36544 26988 36596 26994
rect 36544 26930 36596 26936
rect 36452 26920 36504 26926
rect 36452 26862 36504 26868
rect 36360 26240 36412 26246
rect 36360 26182 36412 26188
rect 35440 26036 35492 26042
rect 35440 25978 35492 25984
rect 35808 26036 35860 26042
rect 35808 25978 35860 25984
rect 36372 25906 36400 26182
rect 34796 25900 34848 25906
rect 34796 25842 34848 25848
rect 36360 25900 36412 25906
rect 36360 25842 36412 25848
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 36464 24954 36492 26862
rect 36636 25832 36688 25838
rect 36636 25774 36688 25780
rect 36452 24948 36504 24954
rect 36452 24890 36504 24896
rect 34704 24608 34756 24614
rect 34704 24550 34756 24556
rect 36452 24608 36504 24614
rect 36452 24550 36504 24556
rect 34520 24404 34572 24410
rect 34520 24346 34572 24352
rect 34244 24200 34296 24206
rect 34244 24142 34296 24148
rect 33784 24064 33836 24070
rect 33784 24006 33836 24012
rect 33796 23730 33824 24006
rect 34256 23730 34284 24142
rect 33784 23724 33836 23730
rect 33784 23666 33836 23672
rect 34244 23724 34296 23730
rect 34244 23666 34296 23672
rect 33692 23656 33744 23662
rect 33692 23598 33744 23604
rect 33600 23180 33652 23186
rect 33600 23122 33652 23128
rect 33416 22500 33468 22506
rect 33416 22442 33468 22448
rect 33612 22094 33640 23122
rect 34716 23118 34744 24550
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 36176 24132 36228 24138
rect 36176 24074 36228 24080
rect 34888 24064 34940 24070
rect 34888 24006 34940 24012
rect 34900 23730 34928 24006
rect 36188 23866 36216 24074
rect 36176 23860 36228 23866
rect 36176 23802 36228 23808
rect 34796 23724 34848 23730
rect 34796 23666 34848 23672
rect 34888 23724 34940 23730
rect 34888 23666 34940 23672
rect 34808 23322 34836 23666
rect 36464 23662 36492 24550
rect 36648 23730 36676 25774
rect 36728 24064 36780 24070
rect 36728 24006 36780 24012
rect 36636 23724 36688 23730
rect 36636 23666 36688 23672
rect 36452 23656 36504 23662
rect 36452 23598 36504 23604
rect 35624 23520 35676 23526
rect 35624 23462 35676 23468
rect 36084 23520 36136 23526
rect 36084 23462 36136 23468
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34796 23316 34848 23322
rect 34796 23258 34848 23264
rect 35636 23186 35664 23462
rect 35624 23180 35676 23186
rect 35624 23122 35676 23128
rect 34704 23112 34756 23118
rect 34704 23054 34756 23060
rect 34152 22704 34204 22710
rect 34152 22646 34204 22652
rect 33784 22636 33836 22642
rect 33784 22578 33836 22584
rect 33796 22234 33824 22578
rect 34060 22500 34112 22506
rect 34060 22442 34112 22448
rect 33784 22228 33836 22234
rect 33784 22170 33836 22176
rect 33336 22066 33456 22094
rect 33324 21956 33376 21962
rect 33324 21898 33376 21904
rect 33336 21690 33364 21898
rect 33140 21684 33192 21690
rect 33140 21626 33192 21632
rect 33324 21684 33376 21690
rect 33324 21626 33376 21632
rect 33152 20058 33180 21626
rect 33140 20052 33192 20058
rect 33140 19994 33192 20000
rect 33140 19712 33192 19718
rect 33140 19654 33192 19660
rect 33152 19378 33180 19654
rect 33324 19508 33376 19514
rect 33324 19450 33376 19456
rect 33140 19372 33192 19378
rect 33140 19314 33192 19320
rect 33336 19156 33364 19450
rect 33428 19446 33456 22066
rect 33520 22066 33640 22094
rect 33416 19440 33468 19446
rect 33416 19382 33468 19388
rect 33244 19128 33364 19156
rect 33048 18692 33100 18698
rect 33048 18634 33100 18640
rect 33048 17332 33100 17338
rect 33048 17274 33100 17280
rect 32772 17264 32824 17270
rect 32772 17206 32824 17212
rect 31760 16516 31812 16522
rect 31760 16458 31812 16464
rect 31772 16182 31800 16458
rect 31760 16176 31812 16182
rect 31760 16118 31812 16124
rect 32312 16108 32364 16114
rect 32312 16050 32364 16056
rect 32404 16108 32456 16114
rect 32404 16050 32456 16056
rect 31760 15904 31812 15910
rect 31760 15846 31812 15852
rect 31772 15502 31800 15846
rect 30840 15496 30892 15502
rect 30840 15438 30892 15444
rect 31484 15496 31536 15502
rect 31484 15438 31536 15444
rect 31576 15496 31628 15502
rect 31576 15438 31628 15444
rect 31760 15496 31812 15502
rect 31760 15438 31812 15444
rect 31496 15162 31524 15438
rect 31484 15156 31536 15162
rect 31484 15098 31536 15104
rect 30472 15020 30524 15026
rect 30472 14962 30524 14968
rect 30564 15020 30616 15026
rect 30564 14962 30616 14968
rect 30484 14618 30512 14962
rect 30472 14612 30524 14618
rect 30472 14554 30524 14560
rect 30380 14340 30432 14346
rect 30380 14282 30432 14288
rect 30564 13864 30616 13870
rect 30564 13806 30616 13812
rect 30380 13728 30432 13734
rect 30380 13670 30432 13676
rect 30392 12918 30420 13670
rect 30472 13456 30524 13462
rect 30472 13398 30524 13404
rect 30484 13326 30512 13398
rect 30472 13320 30524 13326
rect 30472 13262 30524 13268
rect 30380 12912 30432 12918
rect 30380 12854 30432 12860
rect 30576 12306 30604 13806
rect 30668 13258 30696 15030
rect 30760 15026 30880 15042
rect 30760 15020 30892 15026
rect 30760 15014 30840 15020
rect 30760 13462 30788 15014
rect 30840 14962 30892 14968
rect 30748 13456 30800 13462
rect 30748 13398 30800 13404
rect 31024 13456 31076 13462
rect 31024 13398 31076 13404
rect 30656 13252 30708 13258
rect 30656 13194 30708 13200
rect 30564 12300 30616 12306
rect 30564 12242 30616 12248
rect 30288 12232 30340 12238
rect 30288 12174 30340 12180
rect 30104 12164 30156 12170
rect 30104 12106 30156 12112
rect 30300 12102 30328 12174
rect 30288 12096 30340 12102
rect 30288 12038 30340 12044
rect 30576 11744 30604 12242
rect 31036 11898 31064 13398
rect 31392 12640 31444 12646
rect 31392 12582 31444 12588
rect 31404 12238 31432 12582
rect 31392 12232 31444 12238
rect 31392 12174 31444 12180
rect 31024 11892 31076 11898
rect 31024 11834 31076 11840
rect 31036 11762 31064 11834
rect 30656 11756 30708 11762
rect 30576 11716 30656 11744
rect 30656 11698 30708 11704
rect 31024 11756 31076 11762
rect 31024 11698 31076 11704
rect 29472 6886 29684 6914
rect 29932 6886 30328 6914
rect 24860 4616 24912 4622
rect 24860 4558 24912 4564
rect 24872 4078 24900 4558
rect 27160 4140 27212 4146
rect 27160 4082 27212 4088
rect 24860 4072 24912 4078
rect 24860 4014 24912 4020
rect 24768 3936 24820 3942
rect 24768 3878 24820 3884
rect 25964 3936 26016 3942
rect 25964 3878 26016 3884
rect 24780 3058 24808 3878
rect 25976 3602 26004 3878
rect 27172 3738 27200 4082
rect 27344 3936 27396 3942
rect 27344 3878 27396 3884
rect 27160 3732 27212 3738
rect 27160 3674 27212 3680
rect 25964 3596 26016 3602
rect 25964 3538 26016 3544
rect 26424 3596 26476 3602
rect 26424 3538 26476 3544
rect 24768 3052 24820 3058
rect 24768 2994 24820 3000
rect 24952 2984 25004 2990
rect 24952 2926 25004 2932
rect 25780 2984 25832 2990
rect 25780 2926 25832 2932
rect 23572 2916 23624 2922
rect 23572 2858 23624 2864
rect 24964 2650 24992 2926
rect 24952 2644 25004 2650
rect 24952 2586 25004 2592
rect 25792 800 25820 2926
rect 26436 800 26464 3538
rect 27160 3528 27212 3534
rect 27160 3470 27212 3476
rect 27172 3058 27200 3470
rect 27356 3126 27384 3878
rect 27344 3120 27396 3126
rect 27344 3062 27396 3068
rect 27160 3052 27212 3058
rect 27160 2994 27212 3000
rect 27712 2984 27764 2990
rect 27712 2926 27764 2932
rect 27724 800 27752 2926
rect 29656 2650 29684 6886
rect 30300 3670 30328 6886
rect 30288 3664 30340 3670
rect 30288 3606 30340 3612
rect 29644 2644 29696 2650
rect 29644 2586 29696 2592
rect 29000 2372 29052 2378
rect 29000 2314 29052 2320
rect 29012 800 29040 2314
rect 30668 2310 30696 11698
rect 31588 11626 31616 15438
rect 32324 15026 32352 16050
rect 32416 15706 32444 16050
rect 32404 15700 32456 15706
rect 32404 15642 32456 15648
rect 33060 15434 33088 17274
rect 33048 15428 33100 15434
rect 33048 15370 33100 15376
rect 32312 15020 32364 15026
rect 32312 14962 32364 14968
rect 32588 15020 32640 15026
rect 32588 14962 32640 14968
rect 32600 14618 32628 14962
rect 32588 14612 32640 14618
rect 32588 14554 32640 14560
rect 33048 14272 33100 14278
rect 33048 14214 33100 14220
rect 33060 13938 33088 14214
rect 33048 13932 33100 13938
rect 33048 13874 33100 13880
rect 33140 13388 33192 13394
rect 33140 13330 33192 13336
rect 33152 11762 33180 13330
rect 33244 12850 33272 19128
rect 33520 18902 33548 22066
rect 33796 21554 33824 22170
rect 33876 22092 33928 22098
rect 33876 22034 33928 22040
rect 33784 21548 33836 21554
rect 33784 21490 33836 21496
rect 33888 21486 33916 22034
rect 33876 21480 33928 21486
rect 33876 21422 33928 21428
rect 33692 20460 33744 20466
rect 33692 20402 33744 20408
rect 33704 19922 33732 20402
rect 33784 20256 33836 20262
rect 33784 20198 33836 20204
rect 33876 20256 33928 20262
rect 33876 20198 33928 20204
rect 33796 19990 33824 20198
rect 33784 19984 33836 19990
rect 33784 19926 33836 19932
rect 33600 19916 33652 19922
rect 33600 19858 33652 19864
rect 33692 19916 33744 19922
rect 33692 19858 33744 19864
rect 33508 18896 33560 18902
rect 33508 18838 33560 18844
rect 33324 15360 33376 15366
rect 33324 15302 33376 15308
rect 33336 14414 33364 15302
rect 33612 14618 33640 19858
rect 33704 19174 33732 19858
rect 33888 19854 33916 20198
rect 33876 19848 33928 19854
rect 33876 19790 33928 19796
rect 33784 19780 33836 19786
rect 33784 19722 33836 19728
rect 33796 19378 33824 19722
rect 33888 19446 33916 19790
rect 33876 19440 33928 19446
rect 33876 19382 33928 19388
rect 33784 19372 33836 19378
rect 33784 19314 33836 19320
rect 33692 19168 33744 19174
rect 33692 19110 33744 19116
rect 33784 18284 33836 18290
rect 33784 18226 33836 18232
rect 33796 17882 33824 18226
rect 33968 18080 34020 18086
rect 33968 18022 34020 18028
rect 33784 17876 33836 17882
rect 33784 17818 33836 17824
rect 33796 17678 33824 17818
rect 33784 17672 33836 17678
rect 33784 17614 33836 17620
rect 33980 17202 34008 18022
rect 33968 17196 34020 17202
rect 33968 17138 34020 17144
rect 33692 15904 33744 15910
rect 33692 15846 33744 15852
rect 33704 15638 33732 15846
rect 33692 15632 33744 15638
rect 33692 15574 33744 15580
rect 33968 14884 34020 14890
rect 33968 14826 34020 14832
rect 33876 14816 33928 14822
rect 33876 14758 33928 14764
rect 33600 14612 33652 14618
rect 33600 14554 33652 14560
rect 33888 14482 33916 14758
rect 33876 14476 33928 14482
rect 33876 14418 33928 14424
rect 33980 14414 34008 14826
rect 33324 14408 33376 14414
rect 33324 14350 33376 14356
rect 33416 14408 33468 14414
rect 33416 14350 33468 14356
rect 33968 14408 34020 14414
rect 33968 14350 34020 14356
rect 33428 13938 33456 14350
rect 33416 13932 33468 13938
rect 33416 13874 33468 13880
rect 33784 13932 33836 13938
rect 33784 13874 33836 13880
rect 33428 13530 33456 13874
rect 33416 13524 33468 13530
rect 33416 13466 33468 13472
rect 33324 13456 33376 13462
rect 33324 13398 33376 13404
rect 33336 12918 33364 13398
rect 33428 13326 33456 13466
rect 33416 13320 33468 13326
rect 33416 13262 33468 13268
rect 33796 12986 33824 13874
rect 33784 12980 33836 12986
rect 33784 12922 33836 12928
rect 33324 12912 33376 12918
rect 33324 12854 33376 12860
rect 33232 12844 33284 12850
rect 33232 12786 33284 12792
rect 33140 11756 33192 11762
rect 33140 11698 33192 11704
rect 33048 11688 33100 11694
rect 33048 11630 33100 11636
rect 31576 11620 31628 11626
rect 31576 11562 31628 11568
rect 31116 11008 31168 11014
rect 31116 10950 31168 10956
rect 31128 10674 31156 10950
rect 31116 10668 31168 10674
rect 31116 10610 31168 10616
rect 31588 10606 31616 11562
rect 32312 11552 32364 11558
rect 32312 11494 32364 11500
rect 32324 11150 32352 11494
rect 33060 11354 33088 11630
rect 33048 11348 33100 11354
rect 33048 11290 33100 11296
rect 31668 11144 31720 11150
rect 31668 11086 31720 11092
rect 32312 11144 32364 11150
rect 32312 11086 32364 11092
rect 31680 10674 31708 11086
rect 31668 10668 31720 10674
rect 31668 10610 31720 10616
rect 31576 10600 31628 10606
rect 31576 10542 31628 10548
rect 32220 6860 32272 6866
rect 32220 6802 32272 6808
rect 30656 2304 30708 2310
rect 30656 2246 30708 2252
rect 32232 800 32260 6802
rect 32404 6724 32456 6730
rect 32404 6666 32456 6672
rect 32416 6458 32444 6666
rect 32404 6452 32456 6458
rect 32404 6394 32456 6400
rect 33336 3466 33364 12854
rect 33796 12306 33824 12922
rect 33784 12300 33836 12306
rect 33784 12242 33836 12248
rect 33508 12096 33560 12102
rect 33508 12038 33560 12044
rect 33520 11762 33548 12038
rect 33508 11756 33560 11762
rect 33508 11698 33560 11704
rect 33416 11552 33468 11558
rect 33416 11494 33468 11500
rect 33428 10674 33456 11494
rect 33416 10668 33468 10674
rect 33416 10610 33468 10616
rect 34072 3602 34100 22442
rect 34164 21894 34192 22646
rect 35636 22642 35664 23122
rect 35624 22636 35676 22642
rect 35624 22578 35676 22584
rect 34796 22432 34848 22438
rect 34796 22374 34848 22380
rect 35440 22432 35492 22438
rect 35440 22374 35492 22380
rect 34152 21888 34204 21894
rect 34152 21830 34204 21836
rect 34164 21622 34192 21830
rect 34152 21616 34204 21622
rect 34152 21558 34204 21564
rect 34808 20534 34836 22374
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 35452 22030 35480 22374
rect 36096 22098 36124 23462
rect 36360 22976 36412 22982
rect 36360 22918 36412 22924
rect 36372 22710 36400 22918
rect 36360 22704 36412 22710
rect 36360 22646 36412 22652
rect 36372 22098 36400 22646
rect 36084 22092 36136 22098
rect 36084 22034 36136 22040
rect 36360 22092 36412 22098
rect 36360 22034 36412 22040
rect 35256 22024 35308 22030
rect 35256 21966 35308 21972
rect 35440 22024 35492 22030
rect 35440 21966 35492 21972
rect 35268 21690 35296 21966
rect 35624 21956 35676 21962
rect 35624 21898 35676 21904
rect 35532 21888 35584 21894
rect 35532 21830 35584 21836
rect 35256 21684 35308 21690
rect 35256 21626 35308 21632
rect 35268 21298 35296 21626
rect 35544 21554 35572 21830
rect 35532 21548 35584 21554
rect 35532 21490 35584 21496
rect 35268 21270 35388 21298
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 35360 20942 35388 21270
rect 35544 21146 35572 21490
rect 35636 21486 35664 21898
rect 35624 21480 35676 21486
rect 35624 21422 35676 21428
rect 35636 21146 35664 21422
rect 35992 21344 36044 21350
rect 35992 21286 36044 21292
rect 35532 21140 35584 21146
rect 35532 21082 35584 21088
rect 35624 21140 35676 21146
rect 35624 21082 35676 21088
rect 35348 20936 35400 20942
rect 35348 20878 35400 20884
rect 34888 20800 34940 20806
rect 34888 20742 34940 20748
rect 34796 20528 34848 20534
rect 34796 20470 34848 20476
rect 34900 20262 34928 20742
rect 35348 20528 35400 20534
rect 35348 20470 35400 20476
rect 34888 20256 34940 20262
rect 34888 20198 34940 20204
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35360 20058 35388 20470
rect 35900 20460 35952 20466
rect 35900 20402 35952 20408
rect 35912 20058 35940 20402
rect 36004 20262 36032 21286
rect 36096 20346 36124 22034
rect 36096 20318 36308 20346
rect 35992 20256 36044 20262
rect 35992 20198 36044 20204
rect 36176 20256 36228 20262
rect 36176 20198 36228 20204
rect 35348 20052 35400 20058
rect 35348 19994 35400 20000
rect 35900 20052 35952 20058
rect 35900 19994 35952 20000
rect 35440 19848 35492 19854
rect 35440 19790 35492 19796
rect 34704 19508 34756 19514
rect 34704 19450 34756 19456
rect 34428 19372 34480 19378
rect 34428 19314 34480 19320
rect 34440 18358 34468 19314
rect 34428 18352 34480 18358
rect 34428 18294 34480 18300
rect 34716 18154 34744 19450
rect 34796 19168 34848 19174
rect 34796 19110 34848 19116
rect 34808 18834 34836 19110
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34796 18828 34848 18834
rect 34796 18770 34848 18776
rect 35452 18766 35480 19790
rect 35440 18760 35492 18766
rect 35440 18702 35492 18708
rect 34796 18420 34848 18426
rect 34796 18362 34848 18368
rect 34704 18148 34756 18154
rect 34704 18090 34756 18096
rect 34808 17610 34836 18362
rect 35348 18148 35400 18154
rect 35348 18090 35400 18096
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35360 17882 35388 18090
rect 35348 17876 35400 17882
rect 35348 17818 35400 17824
rect 34796 17604 34848 17610
rect 34796 17546 34848 17552
rect 34704 17264 34756 17270
rect 34704 17206 34756 17212
rect 34152 16448 34204 16454
rect 34152 16390 34204 16396
rect 34164 15502 34192 16390
rect 34244 16108 34296 16114
rect 34244 16050 34296 16056
rect 34256 15706 34284 16050
rect 34244 15700 34296 15706
rect 34244 15642 34296 15648
rect 34152 15496 34204 15502
rect 34152 15438 34204 15444
rect 34164 14550 34192 15438
rect 34152 14544 34204 14550
rect 34152 14486 34204 14492
rect 34164 14006 34192 14486
rect 34152 14000 34204 14006
rect 34152 13942 34204 13948
rect 34612 12844 34664 12850
rect 34612 12786 34664 12792
rect 34624 11558 34652 12786
rect 34716 12442 34744 17206
rect 35360 17202 35388 17818
rect 35452 17338 35480 18702
rect 36188 18154 36216 20198
rect 36176 18148 36228 18154
rect 36176 18090 36228 18096
rect 36084 18080 36136 18086
rect 36084 18022 36136 18028
rect 35440 17332 35492 17338
rect 35440 17274 35492 17280
rect 35348 17196 35400 17202
rect 35348 17138 35400 17144
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 36096 16590 36124 18022
rect 36280 17660 36308 20318
rect 36464 18766 36492 23598
rect 36648 23526 36676 23666
rect 36740 23662 36768 24006
rect 36728 23656 36780 23662
rect 36728 23598 36780 23604
rect 36636 23520 36688 23526
rect 36636 23462 36688 23468
rect 36740 23118 36768 23598
rect 36728 23112 36780 23118
rect 36728 23054 36780 23060
rect 36740 22642 36768 23054
rect 36728 22636 36780 22642
rect 36728 22578 36780 22584
rect 36820 22568 36872 22574
rect 36820 22510 36872 22516
rect 36832 22098 36860 22510
rect 36820 22092 36872 22098
rect 37108 22094 37136 27882
rect 37292 25922 37320 29174
rect 37372 28552 37424 28558
rect 37372 28494 37424 28500
rect 37384 26926 37412 28494
rect 37476 28490 37504 30670
rect 37752 30258 37780 31214
rect 37936 30666 37964 31350
rect 37924 30660 37976 30666
rect 37924 30602 37976 30608
rect 37832 30592 37884 30598
rect 37832 30534 37884 30540
rect 37740 30252 37792 30258
rect 37740 30194 37792 30200
rect 37844 29646 37872 30534
rect 38028 29646 38056 31690
rect 38384 31340 38436 31346
rect 38384 31282 38436 31288
rect 38292 30252 38344 30258
rect 38292 30194 38344 30200
rect 37832 29640 37884 29646
rect 37832 29582 37884 29588
rect 38016 29640 38068 29646
rect 38016 29582 38068 29588
rect 37464 28484 37516 28490
rect 37464 28426 37516 28432
rect 37476 27946 37504 28426
rect 37556 28416 37608 28422
rect 37556 28358 37608 28364
rect 37568 28150 37596 28358
rect 37556 28144 37608 28150
rect 37556 28086 37608 28092
rect 37464 27940 37516 27946
rect 37464 27882 37516 27888
rect 37372 26920 37424 26926
rect 37372 26862 37424 26868
rect 37200 25894 37320 25922
rect 37200 25838 37228 25894
rect 37188 25832 37240 25838
rect 37188 25774 37240 25780
rect 37740 24812 37792 24818
rect 37740 24754 37792 24760
rect 37752 23730 37780 24754
rect 37844 24614 37872 29582
rect 38028 29238 38056 29582
rect 38016 29232 38068 29238
rect 38016 29174 38068 29180
rect 38304 29170 38332 30194
rect 38396 30190 38424 31282
rect 38384 30184 38436 30190
rect 38436 30144 38608 30172
rect 38384 30126 38436 30132
rect 38292 29164 38344 29170
rect 38292 29106 38344 29112
rect 37924 29028 37976 29034
rect 37924 28970 37976 28976
rect 38292 29028 38344 29034
rect 38292 28970 38344 28976
rect 38384 29028 38436 29034
rect 38384 28970 38436 28976
rect 37832 24608 37884 24614
rect 37832 24550 37884 24556
rect 37648 23724 37700 23730
rect 37648 23666 37700 23672
rect 37740 23724 37792 23730
rect 37740 23666 37792 23672
rect 37660 23322 37688 23666
rect 37648 23316 37700 23322
rect 37648 23258 37700 23264
rect 37740 23112 37792 23118
rect 37740 23054 37792 23060
rect 37372 22432 37424 22438
rect 37372 22374 37424 22380
rect 37384 22098 37412 22374
rect 37752 22234 37780 23054
rect 37740 22228 37792 22234
rect 37740 22170 37792 22176
rect 37936 22098 37964 28970
rect 38304 28762 38332 28970
rect 38292 28756 38344 28762
rect 38292 28698 38344 28704
rect 38396 27674 38424 28970
rect 38476 28960 38528 28966
rect 38476 28902 38528 28908
rect 38488 28558 38516 28902
rect 38580 28642 38608 30144
rect 38672 29510 38700 35022
rect 38936 34944 38988 34950
rect 38936 34886 38988 34892
rect 38752 34672 38804 34678
rect 38752 34614 38804 34620
rect 38764 34066 38792 34614
rect 38752 34060 38804 34066
rect 38752 34002 38804 34008
rect 38948 33998 38976 34886
rect 39040 34134 39068 35022
rect 39120 34604 39172 34610
rect 39120 34546 39172 34552
rect 39028 34128 39080 34134
rect 39028 34070 39080 34076
rect 39132 33998 39160 34546
rect 39224 34202 39252 35022
rect 39672 34400 39724 34406
rect 39672 34342 39724 34348
rect 39212 34196 39264 34202
rect 39212 34138 39264 34144
rect 39684 34066 39712 34342
rect 40316 34196 40368 34202
rect 40316 34138 40368 34144
rect 39948 34128 40000 34134
rect 40000 34088 40080 34116
rect 39948 34070 40000 34076
rect 39212 34060 39264 34066
rect 39212 34002 39264 34008
rect 39672 34060 39724 34066
rect 39672 34002 39724 34008
rect 38936 33992 38988 33998
rect 38936 33934 38988 33940
rect 39120 33992 39172 33998
rect 39120 33934 39172 33940
rect 38936 32904 38988 32910
rect 38936 32846 38988 32852
rect 39120 32904 39172 32910
rect 39120 32846 39172 32852
rect 38948 31754 38976 32846
rect 39132 32026 39160 32846
rect 39120 32020 39172 32026
rect 39120 31962 39172 31968
rect 39224 31754 39252 34002
rect 40052 32434 40080 34088
rect 40224 32904 40276 32910
rect 40224 32846 40276 32852
rect 40132 32768 40184 32774
rect 40132 32710 40184 32716
rect 39856 32428 39908 32434
rect 39856 32370 39908 32376
rect 40040 32428 40092 32434
rect 40040 32370 40092 32376
rect 39396 32224 39448 32230
rect 39396 32166 39448 32172
rect 39408 31822 39436 32166
rect 39396 31816 39448 31822
rect 39396 31758 39448 31764
rect 38948 31726 39160 31754
rect 39132 31142 39160 31726
rect 39212 31748 39264 31754
rect 39212 31690 39264 31696
rect 39224 31346 39252 31690
rect 39408 31414 39436 31758
rect 39396 31408 39448 31414
rect 39396 31350 39448 31356
rect 39212 31340 39264 31346
rect 39212 31282 39264 31288
rect 39120 31136 39172 31142
rect 39120 31078 39172 31084
rect 39132 30326 39160 31078
rect 39120 30320 39172 30326
rect 39120 30262 39172 30268
rect 38844 30252 38896 30258
rect 38844 30194 38896 30200
rect 38856 30054 38884 30194
rect 39212 30184 39264 30190
rect 39212 30126 39264 30132
rect 39488 30184 39540 30190
rect 39488 30126 39540 30132
rect 38844 30048 38896 30054
rect 38844 29990 38896 29996
rect 38936 30048 38988 30054
rect 38936 29990 38988 29996
rect 38856 29510 38884 29990
rect 38948 29646 38976 29990
rect 38936 29640 38988 29646
rect 38936 29582 38988 29588
rect 39120 29640 39172 29646
rect 39120 29582 39172 29588
rect 38660 29504 38712 29510
rect 38660 29446 38712 29452
rect 38844 29504 38896 29510
rect 38844 29446 38896 29452
rect 38660 29164 38712 29170
rect 38660 29106 38712 29112
rect 38672 28762 38700 29106
rect 39132 28966 39160 29582
rect 39224 29102 39252 30126
rect 39500 29646 39528 30126
rect 39488 29640 39540 29646
rect 39488 29582 39540 29588
rect 39212 29096 39264 29102
rect 39212 29038 39264 29044
rect 39120 28960 39172 28966
rect 39120 28902 39172 28908
rect 38660 28756 38712 28762
rect 38660 28698 38712 28704
rect 38580 28614 38700 28642
rect 38476 28552 38528 28558
rect 38672 28536 38700 28614
rect 39120 28552 39172 28558
rect 38476 28494 38528 28500
rect 38660 28530 38712 28536
rect 39120 28494 39172 28500
rect 38660 28472 38712 28478
rect 39028 27872 39080 27878
rect 39028 27814 39080 27820
rect 38384 27668 38436 27674
rect 38384 27610 38436 27616
rect 38016 27464 38068 27470
rect 38016 27406 38068 27412
rect 38028 27130 38056 27406
rect 38016 27124 38068 27130
rect 38016 27066 38068 27072
rect 38028 26450 38056 27066
rect 38396 26518 38424 27610
rect 38568 26988 38620 26994
rect 38568 26930 38620 26936
rect 38384 26512 38436 26518
rect 38384 26454 38436 26460
rect 38016 26444 38068 26450
rect 38016 26386 38068 26392
rect 38028 25906 38056 26386
rect 38580 26314 38608 26930
rect 38844 26920 38896 26926
rect 38844 26862 38896 26868
rect 38856 26382 38884 26862
rect 38844 26376 38896 26382
rect 38844 26318 38896 26324
rect 38568 26308 38620 26314
rect 38568 26250 38620 26256
rect 38016 25900 38068 25906
rect 38016 25842 38068 25848
rect 38384 25832 38436 25838
rect 38384 25774 38436 25780
rect 38292 25696 38344 25702
rect 38292 25638 38344 25644
rect 38108 24744 38160 24750
rect 38108 24686 38160 24692
rect 38120 24410 38148 24686
rect 38108 24404 38160 24410
rect 38108 24346 38160 24352
rect 37108 22066 37228 22094
rect 36820 22034 36872 22040
rect 36832 21554 36860 22034
rect 36820 21548 36872 21554
rect 36820 21490 36872 21496
rect 36912 21548 36964 21554
rect 36912 21490 36964 21496
rect 36924 21146 36952 21490
rect 36912 21140 36964 21146
rect 36912 21082 36964 21088
rect 36544 20936 36596 20942
rect 36544 20878 36596 20884
rect 36556 20466 36584 20878
rect 36544 20460 36596 20466
rect 36544 20402 36596 20408
rect 36452 18760 36504 18766
rect 36452 18702 36504 18708
rect 36360 18284 36412 18290
rect 36360 18226 36412 18232
rect 36372 17882 36400 18226
rect 36360 17876 36412 17882
rect 36360 17818 36412 17824
rect 36464 17814 36492 18702
rect 36544 18624 36596 18630
rect 36544 18566 36596 18572
rect 36556 18358 36584 18566
rect 36544 18352 36596 18358
rect 36544 18294 36596 18300
rect 36452 17808 36504 17814
rect 36452 17750 36504 17756
rect 36360 17672 36412 17678
rect 36188 17632 36360 17660
rect 36084 16584 36136 16590
rect 36084 16526 36136 16532
rect 36096 16250 36124 16526
rect 36188 16454 36216 17632
rect 36360 17614 36412 17620
rect 36464 17270 36492 17750
rect 36452 17264 36504 17270
rect 36452 17206 36504 17212
rect 36176 16448 36228 16454
rect 36176 16390 36228 16396
rect 36452 16448 36504 16454
rect 36452 16390 36504 16396
rect 36084 16244 36136 16250
rect 36084 16186 36136 16192
rect 36176 16108 36228 16114
rect 36176 16050 36228 16056
rect 35440 15904 35492 15910
rect 35440 15846 35492 15852
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 35452 15570 35480 15846
rect 36188 15638 36216 16050
rect 36360 15904 36412 15910
rect 36360 15846 36412 15852
rect 36176 15632 36228 15638
rect 36176 15574 36228 15580
rect 36372 15570 36400 15846
rect 36464 15570 36492 16390
rect 36820 15700 36872 15706
rect 36820 15642 36872 15648
rect 35440 15564 35492 15570
rect 35440 15506 35492 15512
rect 36360 15564 36412 15570
rect 36360 15506 36412 15512
rect 36452 15564 36504 15570
rect 36452 15506 36504 15512
rect 36176 15360 36228 15366
rect 36176 15302 36228 15308
rect 36188 15026 36216 15302
rect 36372 15026 36400 15506
rect 36832 15366 36860 15642
rect 36820 15360 36872 15366
rect 36820 15302 36872 15308
rect 36832 15026 36860 15302
rect 36176 15020 36228 15026
rect 36176 14962 36228 14968
rect 36360 15020 36412 15026
rect 36360 14962 36412 14968
rect 36820 15020 36872 15026
rect 36820 14962 36872 14968
rect 36912 15020 36964 15026
rect 36912 14962 36964 14968
rect 35440 14884 35492 14890
rect 35440 14826 35492 14832
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35452 14618 35480 14826
rect 35440 14612 35492 14618
rect 35440 14554 35492 14560
rect 34980 14408 35032 14414
rect 34980 14350 35032 14356
rect 34992 14074 35020 14350
rect 34980 14068 35032 14074
rect 34980 14010 35032 14016
rect 34992 13802 35020 14010
rect 36188 14006 36216 14962
rect 36360 14544 36412 14550
rect 36360 14486 36412 14492
rect 36176 14000 36228 14006
rect 36176 13942 36228 13948
rect 34980 13796 35032 13802
rect 34980 13738 35032 13744
rect 35808 13796 35860 13802
rect 35808 13738 35860 13744
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35820 13326 35848 13738
rect 36372 13734 36400 14486
rect 36636 14476 36688 14482
rect 36636 14418 36688 14424
rect 36452 14408 36504 14414
rect 36452 14350 36504 14356
rect 36360 13728 36412 13734
rect 36360 13670 36412 13676
rect 35808 13320 35860 13326
rect 35808 13262 35860 13268
rect 36176 13252 36228 13258
rect 36176 13194 36228 13200
rect 34796 12776 34848 12782
rect 34796 12718 34848 12724
rect 34704 12436 34756 12442
rect 34704 12378 34756 12384
rect 34704 12164 34756 12170
rect 34704 12106 34756 12112
rect 34716 11762 34744 12106
rect 34808 11898 34836 12718
rect 35820 12714 35940 12730
rect 35808 12708 35940 12714
rect 35860 12702 35940 12708
rect 35808 12650 35860 12656
rect 35440 12640 35492 12646
rect 35440 12582 35492 12588
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35452 12238 35480 12582
rect 35912 12442 35940 12702
rect 36188 12646 36216 13194
rect 36372 12646 36400 13670
rect 36464 13394 36492 14350
rect 36452 13388 36504 13394
rect 36452 13330 36504 13336
rect 36464 12782 36492 13330
rect 36648 12850 36676 14418
rect 36728 13320 36780 13326
rect 36728 13262 36780 13268
rect 36740 12986 36768 13262
rect 36832 13190 36860 14962
rect 36924 13530 36952 14962
rect 36912 13524 36964 13530
rect 36912 13466 36964 13472
rect 36820 13184 36872 13190
rect 36820 13126 36872 13132
rect 36728 12980 36780 12986
rect 36728 12922 36780 12928
rect 36636 12844 36688 12850
rect 36636 12786 36688 12792
rect 36452 12776 36504 12782
rect 36452 12718 36504 12724
rect 36176 12640 36228 12646
rect 36176 12582 36228 12588
rect 36360 12640 36412 12646
rect 36360 12582 36412 12588
rect 35900 12436 35952 12442
rect 35900 12378 35952 12384
rect 36360 12436 36412 12442
rect 36360 12378 36412 12384
rect 35992 12300 36044 12306
rect 35992 12242 36044 12248
rect 35348 12232 35400 12238
rect 35348 12174 35400 12180
rect 35440 12232 35492 12238
rect 35440 12174 35492 12180
rect 34796 11892 34848 11898
rect 34796 11834 34848 11840
rect 34704 11756 34756 11762
rect 34704 11698 34756 11704
rect 34612 11552 34664 11558
rect 34612 11494 34664 11500
rect 34624 11354 34652 11494
rect 34612 11348 34664 11354
rect 34612 11290 34664 11296
rect 34716 11218 34744 11698
rect 35360 11626 35388 12174
rect 35452 11830 35480 12174
rect 35532 12096 35584 12102
rect 35532 12038 35584 12044
rect 35440 11824 35492 11830
rect 35440 11766 35492 11772
rect 35544 11762 35572 12038
rect 36004 11762 36032 12242
rect 36372 12238 36400 12378
rect 36360 12232 36412 12238
rect 36360 12174 36412 12180
rect 36648 11762 36676 12786
rect 36924 11898 36952 13466
rect 37200 13462 37228 22066
rect 37372 22092 37424 22098
rect 37372 22034 37424 22040
rect 37924 22092 37976 22098
rect 37924 22034 37976 22040
rect 37384 20942 37412 22034
rect 37936 21554 37964 22034
rect 38304 22030 38332 25638
rect 38396 25430 38424 25774
rect 38580 25770 38608 26250
rect 38856 25906 38884 26318
rect 39040 25906 39068 27814
rect 39132 27674 39160 28494
rect 39224 28150 39252 29038
rect 39212 28144 39264 28150
rect 39212 28086 39264 28092
rect 39868 28014 39896 32370
rect 40040 31884 40092 31890
rect 40040 31826 40092 31832
rect 40052 29714 40080 31826
rect 40144 31822 40172 32710
rect 40236 32570 40264 32846
rect 40224 32564 40276 32570
rect 40224 32506 40276 32512
rect 40328 32434 40356 34138
rect 40408 33992 40460 33998
rect 40408 33934 40460 33940
rect 40420 33114 40448 33934
rect 40408 33108 40460 33114
rect 40408 33050 40460 33056
rect 41328 32904 41380 32910
rect 41328 32846 41380 32852
rect 40316 32428 40368 32434
rect 40316 32370 40368 32376
rect 41340 32026 41368 32846
rect 41328 32020 41380 32026
rect 41328 31962 41380 31968
rect 40132 31816 40184 31822
rect 40132 31758 40184 31764
rect 41236 30592 41288 30598
rect 41236 30534 41288 30540
rect 40132 30388 40184 30394
rect 40132 30330 40184 30336
rect 40040 29708 40092 29714
rect 40040 29650 40092 29656
rect 40052 28150 40080 29650
rect 40144 28626 40172 30330
rect 40684 30252 40736 30258
rect 40684 30194 40736 30200
rect 40776 30252 40828 30258
rect 40776 30194 40828 30200
rect 40592 30184 40644 30190
rect 40592 30126 40644 30132
rect 40224 30116 40276 30122
rect 40224 30058 40276 30064
rect 40236 29238 40264 30058
rect 40500 29504 40552 29510
rect 40500 29446 40552 29452
rect 40224 29232 40276 29238
rect 40276 29180 40448 29186
rect 40224 29174 40448 29180
rect 40236 29158 40448 29174
rect 40224 29028 40276 29034
rect 40224 28970 40276 28976
rect 40132 28620 40184 28626
rect 40132 28562 40184 28568
rect 40236 28558 40264 28970
rect 40316 28688 40368 28694
rect 40316 28630 40368 28636
rect 40224 28552 40276 28558
rect 40224 28494 40276 28500
rect 40040 28144 40092 28150
rect 40040 28086 40092 28092
rect 40132 28076 40184 28082
rect 40132 28018 40184 28024
rect 39856 28008 39908 28014
rect 39856 27950 39908 27956
rect 39120 27668 39172 27674
rect 39120 27610 39172 27616
rect 39672 27328 39724 27334
rect 39672 27270 39724 27276
rect 39684 26926 39712 27270
rect 39672 26920 39724 26926
rect 39672 26862 39724 26868
rect 39684 26450 39712 26862
rect 39672 26444 39724 26450
rect 39672 26386 39724 26392
rect 40144 25974 40172 28018
rect 40328 27690 40356 28630
rect 40420 28558 40448 29158
rect 40408 28552 40460 28558
rect 40408 28494 40460 28500
rect 40512 28490 40540 29446
rect 40604 29170 40632 30126
rect 40696 29238 40724 30194
rect 40788 29646 40816 30194
rect 40776 29640 40828 29646
rect 40776 29582 40828 29588
rect 40684 29232 40736 29238
rect 40684 29174 40736 29180
rect 40592 29164 40644 29170
rect 40592 29106 40644 29112
rect 40696 29034 40724 29174
rect 40788 29170 40816 29582
rect 40776 29164 40828 29170
rect 40776 29106 40828 29112
rect 40684 29028 40736 29034
rect 40684 28970 40736 28976
rect 40500 28484 40552 28490
rect 40500 28426 40552 28432
rect 40684 28144 40736 28150
rect 40684 28086 40736 28092
rect 40236 27662 40356 27690
rect 40696 27674 40724 28086
rect 40684 27668 40736 27674
rect 40236 27470 40264 27662
rect 40684 27610 40736 27616
rect 40316 27600 40368 27606
rect 40316 27542 40368 27548
rect 40224 27464 40276 27470
rect 40224 27406 40276 27412
rect 40236 27062 40264 27406
rect 40224 27056 40276 27062
rect 40224 26998 40276 27004
rect 40236 26450 40264 26998
rect 40224 26444 40276 26450
rect 40224 26386 40276 26392
rect 40224 26308 40276 26314
rect 40224 26250 40276 26256
rect 40132 25968 40184 25974
rect 40132 25910 40184 25916
rect 38844 25900 38896 25906
rect 38844 25842 38896 25848
rect 39028 25900 39080 25906
rect 39028 25842 39080 25848
rect 38568 25764 38620 25770
rect 38568 25706 38620 25712
rect 38660 25764 38712 25770
rect 38660 25706 38712 25712
rect 38384 25424 38436 25430
rect 38384 25366 38436 25372
rect 38580 24750 38608 25706
rect 38672 24818 38700 25706
rect 39040 25276 39068 25842
rect 40144 25294 40172 25910
rect 40236 25838 40264 26250
rect 40328 25906 40356 27542
rect 41248 27402 41276 30534
rect 41340 30258 41368 31962
rect 42616 31340 42668 31346
rect 42616 31282 42668 31288
rect 42628 30938 42656 31282
rect 42892 31272 42944 31278
rect 42892 31214 42944 31220
rect 42616 30932 42668 30938
rect 42616 30874 42668 30880
rect 42904 30870 42932 31214
rect 42892 30864 42944 30870
rect 42892 30806 42944 30812
rect 42800 30592 42852 30598
rect 42800 30534 42852 30540
rect 43536 30592 43588 30598
rect 43536 30534 43588 30540
rect 41328 30252 41380 30258
rect 41328 30194 41380 30200
rect 42812 29170 42840 30534
rect 43352 30252 43404 30258
rect 43352 30194 43404 30200
rect 43364 30122 43392 30194
rect 43444 30184 43496 30190
rect 43444 30126 43496 30132
rect 43168 30116 43220 30122
rect 43168 30058 43220 30064
rect 43352 30116 43404 30122
rect 43352 30058 43404 30064
rect 42984 29708 43036 29714
rect 42984 29650 43036 29656
rect 42892 29640 42944 29646
rect 42892 29582 42944 29588
rect 42800 29164 42852 29170
rect 42800 29106 42852 29112
rect 42064 28620 42116 28626
rect 42064 28562 42116 28568
rect 41788 28416 41840 28422
rect 41788 28358 41840 28364
rect 41420 27940 41472 27946
rect 41420 27882 41472 27888
rect 41236 27396 41288 27402
rect 41236 27338 41288 27344
rect 41432 26994 41460 27882
rect 41800 27470 41828 28358
rect 42076 28082 42104 28562
rect 42800 28552 42852 28558
rect 42800 28494 42852 28500
rect 42812 28218 42840 28494
rect 42800 28212 42852 28218
rect 42800 28154 42852 28160
rect 42064 28076 42116 28082
rect 42064 28018 42116 28024
rect 42076 27878 42104 28018
rect 42800 28008 42852 28014
rect 42800 27950 42852 27956
rect 42064 27872 42116 27878
rect 42064 27814 42116 27820
rect 41788 27464 41840 27470
rect 41788 27406 41840 27412
rect 41512 27396 41564 27402
rect 41512 27338 41564 27344
rect 41420 26988 41472 26994
rect 41420 26930 41472 26936
rect 40500 26784 40552 26790
rect 40500 26726 40552 26732
rect 40512 26042 40540 26726
rect 40868 26376 40920 26382
rect 40868 26318 40920 26324
rect 40500 26036 40552 26042
rect 40500 25978 40552 25984
rect 40316 25900 40368 25906
rect 40316 25842 40368 25848
rect 40224 25832 40276 25838
rect 40224 25774 40276 25780
rect 40132 25288 40184 25294
rect 39040 25248 39344 25276
rect 38660 24812 38712 24818
rect 38660 24754 38712 24760
rect 38844 24812 38896 24818
rect 38844 24754 38896 24760
rect 38568 24744 38620 24750
rect 38568 24686 38620 24692
rect 38660 24608 38712 24614
rect 38660 24550 38712 24556
rect 38672 23050 38700 24550
rect 38856 23866 38884 24754
rect 39212 24608 39264 24614
rect 39212 24550 39264 24556
rect 38936 24200 38988 24206
rect 38936 24142 38988 24148
rect 38844 23860 38896 23866
rect 38844 23802 38896 23808
rect 38660 23044 38712 23050
rect 38660 22986 38712 22992
rect 38948 22642 38976 24142
rect 39224 24138 39252 24550
rect 39120 24132 39172 24138
rect 39120 24074 39172 24080
rect 39212 24132 39264 24138
rect 39212 24074 39264 24080
rect 39028 23860 39080 23866
rect 39028 23802 39080 23808
rect 39040 23594 39068 23802
rect 39132 23730 39160 24074
rect 39120 23724 39172 23730
rect 39120 23666 39172 23672
rect 39028 23588 39080 23594
rect 39028 23530 39080 23536
rect 38936 22636 38988 22642
rect 38936 22578 38988 22584
rect 39028 22636 39080 22642
rect 39028 22578 39080 22584
rect 39040 22234 39068 22578
rect 39028 22228 39080 22234
rect 39028 22170 39080 22176
rect 38292 22024 38344 22030
rect 38292 21966 38344 21972
rect 39212 22024 39264 22030
rect 39212 21966 39264 21972
rect 38304 21690 38332 21966
rect 38292 21684 38344 21690
rect 38292 21626 38344 21632
rect 37924 21548 37976 21554
rect 37924 21490 37976 21496
rect 39224 21418 39252 21966
rect 39212 21412 39264 21418
rect 39212 21354 39264 21360
rect 37556 21344 37608 21350
rect 37556 21286 37608 21292
rect 37372 20936 37424 20942
rect 37372 20878 37424 20884
rect 37568 16794 37596 21286
rect 37740 20392 37792 20398
rect 37740 20334 37792 20340
rect 37752 19310 37780 20334
rect 39212 19848 39264 19854
rect 39212 19790 39264 19796
rect 37740 19304 37792 19310
rect 37740 19246 37792 19252
rect 37752 18766 37780 19246
rect 39224 18970 39252 19790
rect 39212 18964 39264 18970
rect 39212 18906 39264 18912
rect 37740 18760 37792 18766
rect 37740 18702 37792 18708
rect 37752 18358 37780 18702
rect 37740 18352 37792 18358
rect 37740 18294 37792 18300
rect 37752 17746 37780 18294
rect 37740 17740 37792 17746
rect 37740 17682 37792 17688
rect 37556 16788 37608 16794
rect 37556 16730 37608 16736
rect 37280 16652 37332 16658
rect 37280 16594 37332 16600
rect 37292 16182 37320 16594
rect 37568 16250 37596 16730
rect 37556 16244 37608 16250
rect 37556 16186 37608 16192
rect 37280 16176 37332 16182
rect 37280 16118 37332 16124
rect 37740 16108 37792 16114
rect 37740 16050 37792 16056
rect 37556 15564 37608 15570
rect 37556 15506 37608 15512
rect 37568 14958 37596 15506
rect 37752 15162 37780 16050
rect 38476 15496 38528 15502
rect 38476 15438 38528 15444
rect 37740 15156 37792 15162
rect 37740 15098 37792 15104
rect 37556 14952 37608 14958
rect 37556 14894 37608 14900
rect 37648 14272 37700 14278
rect 37648 14214 37700 14220
rect 37188 13456 37240 13462
rect 37188 13398 37240 13404
rect 37660 13394 37688 14214
rect 38488 13394 38516 15438
rect 37648 13388 37700 13394
rect 37648 13330 37700 13336
rect 38476 13388 38528 13394
rect 38476 13330 38528 13336
rect 37832 13320 37884 13326
rect 37832 13262 37884 13268
rect 37372 13184 37424 13190
rect 37372 13126 37424 13132
rect 37004 12980 37056 12986
rect 37004 12922 37056 12928
rect 37016 12306 37044 12922
rect 37384 12918 37412 13126
rect 37372 12912 37424 12918
rect 37372 12854 37424 12860
rect 37556 12708 37608 12714
rect 37556 12650 37608 12656
rect 37464 12640 37516 12646
rect 37464 12582 37516 12588
rect 37004 12300 37056 12306
rect 37004 12242 37056 12248
rect 37476 12238 37504 12582
rect 37464 12232 37516 12238
rect 37464 12174 37516 12180
rect 36912 11892 36964 11898
rect 36912 11834 36964 11840
rect 35532 11756 35584 11762
rect 35532 11698 35584 11704
rect 35992 11756 36044 11762
rect 35992 11698 36044 11704
rect 36268 11756 36320 11762
rect 36268 11698 36320 11704
rect 36636 11756 36688 11762
rect 36636 11698 36688 11704
rect 35348 11620 35400 11626
rect 35348 11562 35400 11568
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 35544 11354 35572 11698
rect 36280 11354 36308 11698
rect 35532 11348 35584 11354
rect 35532 11290 35584 11296
rect 36268 11348 36320 11354
rect 36268 11290 36320 11296
rect 34704 11212 34756 11218
rect 34704 11154 34756 11160
rect 34716 10810 34744 11154
rect 37476 11082 37504 12174
rect 37568 11898 37596 12650
rect 37844 12442 37872 13262
rect 37832 12436 37884 12442
rect 37832 12378 37884 12384
rect 39316 12306 39344 25248
rect 40132 25230 40184 25236
rect 40880 25226 40908 26318
rect 40868 25220 40920 25226
rect 40868 25162 40920 25168
rect 39488 25152 39540 25158
rect 39488 25094 39540 25100
rect 39500 23730 39528 25094
rect 40880 24206 40908 25162
rect 41432 25158 41460 26930
rect 41420 25152 41472 25158
rect 41420 25094 41472 25100
rect 40868 24200 40920 24206
rect 40868 24142 40920 24148
rect 39488 23724 39540 23730
rect 39488 23666 39540 23672
rect 39396 23656 39448 23662
rect 39396 23598 39448 23604
rect 39500 23610 39528 23666
rect 39408 22094 39436 23598
rect 39500 23582 39620 23610
rect 39408 22066 39528 22094
rect 39500 22030 39528 22066
rect 39488 22024 39540 22030
rect 39488 21966 39540 21972
rect 39304 12300 39356 12306
rect 39304 12242 39356 12248
rect 37556 11892 37608 11898
rect 37556 11834 37608 11840
rect 37648 11756 37700 11762
rect 37648 11698 37700 11704
rect 37660 11286 37688 11698
rect 37648 11280 37700 11286
rect 37648 11222 37700 11228
rect 37464 11076 37516 11082
rect 37464 11018 37516 11024
rect 34704 10804 34756 10810
rect 34704 10746 34756 10752
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 39592 9178 39620 23582
rect 40408 23520 40460 23526
rect 40408 23462 40460 23468
rect 40420 23186 40448 23462
rect 39856 23180 39908 23186
rect 39856 23122 39908 23128
rect 40408 23180 40460 23186
rect 40408 23122 40460 23128
rect 39868 19360 39896 23122
rect 40316 22432 40368 22438
rect 40316 22374 40368 22380
rect 40328 22030 40356 22374
rect 40316 22024 40368 22030
rect 40316 21966 40368 21972
rect 40960 21888 41012 21894
rect 40960 21830 41012 21836
rect 40592 20596 40644 20602
rect 40592 20538 40644 20544
rect 39948 20460 40000 20466
rect 39948 20402 40000 20408
rect 39960 19786 39988 20402
rect 40132 20392 40184 20398
rect 40132 20334 40184 20340
rect 40144 19854 40172 20334
rect 40132 19848 40184 19854
rect 40132 19790 40184 19796
rect 40500 19848 40552 19854
rect 40604 19836 40632 20538
rect 40776 20324 40828 20330
rect 40776 20266 40828 20272
rect 40788 19854 40816 20266
rect 40552 19808 40632 19836
rect 40500 19790 40552 19796
rect 39948 19780 40000 19786
rect 39948 19722 40000 19728
rect 40132 19712 40184 19718
rect 40132 19654 40184 19660
rect 39948 19372 40000 19378
rect 39868 19332 39948 19360
rect 39868 15502 39896 19332
rect 39948 19314 40000 19320
rect 40144 19258 40172 19654
rect 40224 19508 40276 19514
rect 40224 19450 40276 19456
rect 40236 19310 40264 19450
rect 40408 19440 40460 19446
rect 40408 19382 40460 19388
rect 39960 19242 40172 19258
rect 40224 19304 40276 19310
rect 40224 19246 40276 19252
rect 39948 19236 40172 19242
rect 40000 19230 40172 19236
rect 39948 19178 40000 19184
rect 39960 18970 39988 19178
rect 39948 18964 40000 18970
rect 39948 18906 40000 18912
rect 40236 18834 40264 19246
rect 40316 18896 40368 18902
rect 40316 18838 40368 18844
rect 40224 18828 40276 18834
rect 40224 18770 40276 18776
rect 40040 18760 40092 18766
rect 40040 18702 40092 18708
rect 40052 18358 40080 18702
rect 40224 18692 40276 18698
rect 40224 18634 40276 18640
rect 40236 18358 40264 18634
rect 40040 18352 40092 18358
rect 40040 18294 40092 18300
rect 40224 18352 40276 18358
rect 40224 18294 40276 18300
rect 40052 17882 40080 18294
rect 40040 17876 40092 17882
rect 40040 17818 40092 17824
rect 40328 17678 40356 18838
rect 40420 18426 40448 19382
rect 40604 19378 40632 19808
rect 40776 19848 40828 19854
rect 40776 19790 40828 19796
rect 40788 19530 40816 19790
rect 40788 19502 40908 19530
rect 40592 19372 40644 19378
rect 40592 19314 40644 19320
rect 40604 18952 40632 19314
rect 40776 19304 40828 19310
rect 40776 19246 40828 19252
rect 40788 18970 40816 19246
rect 40880 19174 40908 19502
rect 40972 19378 41000 21830
rect 41524 20534 41552 27338
rect 42076 26926 42104 27814
rect 42812 27334 42840 27950
rect 42800 27328 42852 27334
rect 42800 27270 42852 27276
rect 42064 26920 42116 26926
rect 42064 26862 42116 26868
rect 41788 25424 41840 25430
rect 41788 25366 41840 25372
rect 41800 24818 41828 25366
rect 42340 25288 42392 25294
rect 42340 25230 42392 25236
rect 42064 25220 42116 25226
rect 42064 25162 42116 25168
rect 41972 25152 42024 25158
rect 41972 25094 42024 25100
rect 41984 24954 42012 25094
rect 41972 24948 42024 24954
rect 41972 24890 42024 24896
rect 41788 24812 41840 24818
rect 41788 24754 41840 24760
rect 41604 24608 41656 24614
rect 41604 24550 41656 24556
rect 41616 24138 41644 24550
rect 42076 24410 42104 25162
rect 42064 24404 42116 24410
rect 42064 24346 42116 24352
rect 42352 24138 42380 25230
rect 42708 24608 42760 24614
rect 42708 24550 42760 24556
rect 42720 24206 42748 24550
rect 42708 24200 42760 24206
rect 42708 24142 42760 24148
rect 41604 24132 41656 24138
rect 41604 24074 41656 24080
rect 42340 24132 42392 24138
rect 42340 24074 42392 24080
rect 42352 23322 42380 24074
rect 42340 23316 42392 23322
rect 42340 23258 42392 23264
rect 41788 22636 41840 22642
rect 41788 22578 41840 22584
rect 41696 22568 41748 22574
rect 41696 22510 41748 22516
rect 41708 21962 41736 22510
rect 41800 22234 41828 22578
rect 42432 22432 42484 22438
rect 42432 22374 42484 22380
rect 41788 22228 41840 22234
rect 41788 22170 41840 22176
rect 42444 22030 42472 22374
rect 42720 22030 42748 24142
rect 42812 24070 42840 27270
rect 42904 26994 42932 29582
rect 42996 27878 43024 29650
rect 43180 29102 43208 30058
rect 43260 30048 43312 30054
rect 43260 29990 43312 29996
rect 43272 29102 43300 29990
rect 43456 29646 43484 30126
rect 43548 29714 43576 30534
rect 43536 29708 43588 29714
rect 43536 29650 43588 29656
rect 43444 29640 43496 29646
rect 43496 29588 43576 29594
rect 43444 29582 43576 29588
rect 43456 29566 43576 29582
rect 43548 29238 43576 29566
rect 43536 29232 43588 29238
rect 43536 29174 43588 29180
rect 43168 29096 43220 29102
rect 43168 29038 43220 29044
rect 43260 29096 43312 29102
rect 43260 29038 43312 29044
rect 43180 28218 43208 29038
rect 43168 28212 43220 28218
rect 43168 28154 43220 28160
rect 42984 27872 43036 27878
rect 42984 27814 43036 27820
rect 42892 26988 42944 26994
rect 42892 26930 42944 26936
rect 42904 25294 42932 26930
rect 42984 26920 43036 26926
rect 42984 26862 43036 26868
rect 42892 25288 42944 25294
rect 42892 25230 42944 25236
rect 42904 24750 42932 25230
rect 42892 24744 42944 24750
rect 42892 24686 42944 24692
rect 42996 24562 43024 26862
rect 43076 25832 43128 25838
rect 43076 25774 43128 25780
rect 43088 25498 43116 25774
rect 43076 25492 43128 25498
rect 43076 25434 43128 25440
rect 43180 25378 43208 28154
rect 43272 28082 43300 29038
rect 43352 29028 43404 29034
rect 43352 28970 43404 28976
rect 43364 28626 43392 28970
rect 43352 28620 43404 28626
rect 43352 28562 43404 28568
rect 43260 28076 43312 28082
rect 43260 28018 43312 28024
rect 43364 27470 43392 28562
rect 43548 28422 43576 29174
rect 43536 28416 43588 28422
rect 43536 28358 43588 28364
rect 43548 28014 43576 28358
rect 43536 28008 43588 28014
rect 43536 27950 43588 27956
rect 43352 27464 43404 27470
rect 43352 27406 43404 27412
rect 43548 25498 43576 27950
rect 43536 25492 43588 25498
rect 43536 25434 43588 25440
rect 43352 25424 43404 25430
rect 43180 25372 43352 25378
rect 43180 25366 43404 25372
rect 43180 25350 43392 25366
rect 43076 25152 43128 25158
rect 43076 25094 43128 25100
rect 43088 24750 43116 25094
rect 43168 24812 43220 24818
rect 43168 24754 43220 24760
rect 43076 24744 43128 24750
rect 43076 24686 43128 24692
rect 42904 24534 43024 24562
rect 42800 24064 42852 24070
rect 42800 24006 42852 24012
rect 42800 23520 42852 23526
rect 42800 23462 42852 23468
rect 42812 22778 42840 23462
rect 42904 22778 42932 24534
rect 43180 24274 43208 24754
rect 43272 24750 43300 25350
rect 43444 25288 43496 25294
rect 43444 25230 43496 25236
rect 43456 25158 43484 25230
rect 43444 25152 43496 25158
rect 43444 25094 43496 25100
rect 43456 24970 43484 25094
rect 43456 24942 43576 24970
rect 43548 24886 43576 24942
rect 43536 24880 43588 24886
rect 43536 24822 43588 24828
rect 43444 24812 43496 24818
rect 43444 24754 43496 24760
rect 43260 24744 43312 24750
rect 43260 24686 43312 24692
rect 43352 24744 43404 24750
rect 43352 24686 43404 24692
rect 43168 24268 43220 24274
rect 43168 24210 43220 24216
rect 43272 23730 43300 24686
rect 43364 24206 43392 24686
rect 43456 24614 43484 24754
rect 43444 24608 43496 24614
rect 43444 24550 43496 24556
rect 43548 24410 43576 24822
rect 43536 24404 43588 24410
rect 43536 24346 43588 24352
rect 43352 24200 43404 24206
rect 43352 24142 43404 24148
rect 43640 23866 43668 47126
rect 46294 47016 46350 47025
rect 46294 46951 46350 46960
rect 45928 46504 45980 46510
rect 45928 46446 45980 46452
rect 45836 46436 45888 46442
rect 45836 46378 45888 46384
rect 45558 46336 45614 46345
rect 45558 46271 45614 46280
rect 45572 40458 45600 46271
rect 45848 45490 45876 46378
rect 45940 46170 45968 46446
rect 45928 46164 45980 46170
rect 45928 46106 45980 46112
rect 46020 45960 46072 45966
rect 46020 45902 46072 45908
rect 45836 45484 45888 45490
rect 45836 45426 45888 45432
rect 46032 44878 46060 45902
rect 46308 45422 46336 46951
rect 46400 46510 46428 49200
rect 46754 49056 46810 49065
rect 46754 48991 46810 49000
rect 46768 47122 46796 48991
rect 46756 47116 46808 47122
rect 46756 47058 46808 47064
rect 47216 47048 47268 47054
rect 47216 46990 47268 46996
rect 47032 46980 47084 46986
rect 47032 46922 47084 46928
rect 46388 46504 46440 46510
rect 46388 46446 46440 46452
rect 46664 46368 46716 46374
rect 46664 46310 46716 46316
rect 46676 46034 46704 46310
rect 46664 46028 46716 46034
rect 46664 45970 46716 45976
rect 47044 45558 47072 46922
rect 46940 45552 46992 45558
rect 46940 45494 46992 45500
rect 47032 45552 47084 45558
rect 47032 45494 47084 45500
rect 46296 45416 46348 45422
rect 46296 45358 46348 45364
rect 46846 44976 46902 44985
rect 46846 44911 46848 44920
rect 46900 44911 46902 44920
rect 46848 44882 46900 44888
rect 46020 44872 46072 44878
rect 46020 44814 46072 44820
rect 46388 44872 46440 44878
rect 46388 44814 46440 44820
rect 45560 40452 45612 40458
rect 45560 40394 45612 40400
rect 46400 39982 46428 44814
rect 46952 44470 46980 45494
rect 46940 44464 46992 44470
rect 46940 44406 46992 44412
rect 46480 42016 46532 42022
rect 46480 41958 46532 41964
rect 46492 41682 46520 41958
rect 46480 41676 46532 41682
rect 46480 41618 46532 41624
rect 46952 41138 46980 44406
rect 47228 44402 47256 46990
rect 47216 44396 47268 44402
rect 47216 44338 47268 44344
rect 47032 43104 47084 43110
rect 47032 43046 47084 43052
rect 47044 42770 47072 43046
rect 47032 42764 47084 42770
rect 47032 42706 47084 42712
rect 47124 41540 47176 41546
rect 47124 41482 47176 41488
rect 47136 41274 47164 41482
rect 47124 41268 47176 41274
rect 47124 41210 47176 41216
rect 46940 41132 46992 41138
rect 46940 41074 46992 41080
rect 46480 40928 46532 40934
rect 46480 40870 46532 40876
rect 46492 40594 46520 40870
rect 46480 40588 46532 40594
rect 46480 40530 46532 40536
rect 46388 39976 46440 39982
rect 46388 39918 46440 39924
rect 46846 39536 46902 39545
rect 46846 39471 46848 39480
rect 46900 39471 46902 39480
rect 46848 39442 46900 39448
rect 46478 38176 46534 38185
rect 46478 38111 46534 38120
rect 46492 37262 46520 38111
rect 46952 37874 46980 41074
rect 47124 40452 47176 40458
rect 47124 40394 47176 40400
rect 47136 40050 47164 40394
rect 47124 40044 47176 40050
rect 47124 39986 47176 39992
rect 46940 37868 46992 37874
rect 46940 37810 46992 37816
rect 46480 37256 46532 37262
rect 46480 37198 46532 37204
rect 46848 36236 46900 36242
rect 46848 36178 46900 36184
rect 46860 36145 46888 36178
rect 46846 36136 46902 36145
rect 46846 36071 46902 36080
rect 47124 35692 47176 35698
rect 47124 35634 47176 35640
rect 46940 33516 46992 33522
rect 46940 33458 46992 33464
rect 46952 33386 46980 33458
rect 46940 33380 46992 33386
rect 46940 33322 46992 33328
rect 46756 33040 46808 33046
rect 46756 32982 46808 32988
rect 46480 32904 46532 32910
rect 46480 32846 46532 32852
rect 45560 32768 45612 32774
rect 45560 32710 45612 32716
rect 45572 32502 45600 32710
rect 46492 32502 46520 32846
rect 45560 32496 45612 32502
rect 45560 32438 45612 32444
rect 46480 32496 46532 32502
rect 46480 32438 46532 32444
rect 44640 32428 44692 32434
rect 44640 32370 44692 32376
rect 44456 31476 44508 31482
rect 44456 31418 44508 31424
rect 44088 30864 44140 30870
rect 44088 30806 44140 30812
rect 43720 30592 43772 30598
rect 43720 30534 43772 30540
rect 43732 29170 43760 30534
rect 43904 30048 43956 30054
rect 43904 29990 43956 29996
rect 43916 29646 43944 29990
rect 43904 29640 43956 29646
rect 43904 29582 43956 29588
rect 43720 29164 43772 29170
rect 43720 29106 43772 29112
rect 43732 28558 43760 29106
rect 43904 29096 43956 29102
rect 43904 29038 43956 29044
rect 43916 28558 43944 29038
rect 43720 28552 43772 28558
rect 43720 28494 43772 28500
rect 43904 28552 43956 28558
rect 43904 28494 43956 28500
rect 43732 28082 43760 28494
rect 43812 28484 43864 28490
rect 43812 28426 43864 28432
rect 43824 28218 43852 28426
rect 43812 28212 43864 28218
rect 43812 28154 43864 28160
rect 43720 28076 43772 28082
rect 43720 28018 43772 28024
rect 43916 27878 43944 28494
rect 43996 28416 44048 28422
rect 43996 28358 44048 28364
rect 43904 27872 43956 27878
rect 43904 27814 43956 27820
rect 43916 27674 43944 27814
rect 43904 27668 43956 27674
rect 43904 27610 43956 27616
rect 44008 27402 44036 28358
rect 44100 28082 44128 30806
rect 44468 30734 44496 31418
rect 44456 30728 44508 30734
rect 44456 30670 44508 30676
rect 44180 30660 44232 30666
rect 44180 30602 44232 30608
rect 44548 30660 44600 30666
rect 44548 30602 44600 30608
rect 44192 30394 44220 30602
rect 44180 30388 44232 30394
rect 44180 30330 44232 30336
rect 44560 30326 44588 30602
rect 44548 30320 44600 30326
rect 44548 30262 44600 30268
rect 44180 30252 44232 30258
rect 44180 30194 44232 30200
rect 44192 29578 44220 30194
rect 44652 29782 44680 32370
rect 45376 32360 45428 32366
rect 45376 32302 45428 32308
rect 45388 31482 45416 32302
rect 46020 32224 46072 32230
rect 46020 32166 46072 32172
rect 46032 31890 46060 32166
rect 46020 31884 46072 31890
rect 46020 31826 46072 31832
rect 45836 31816 45888 31822
rect 45836 31758 45888 31764
rect 45376 31476 45428 31482
rect 45376 31418 45428 31424
rect 44732 31340 44784 31346
rect 44732 31282 44784 31288
rect 44744 29850 44772 31282
rect 44916 31136 44968 31142
rect 44916 31078 44968 31084
rect 44928 30734 44956 31078
rect 45848 30938 45876 31758
rect 45836 30932 45888 30938
rect 45836 30874 45888 30880
rect 44916 30728 44968 30734
rect 44916 30670 44968 30676
rect 45848 30666 45876 30874
rect 45836 30660 45888 30666
rect 45836 30602 45888 30608
rect 46480 30048 46532 30054
rect 46480 29990 46532 29996
rect 44732 29844 44784 29850
rect 44732 29786 44784 29792
rect 44640 29776 44692 29782
rect 44640 29718 44692 29724
rect 44180 29572 44232 29578
rect 44180 29514 44232 29520
rect 44652 29034 44680 29718
rect 46492 29714 46520 29990
rect 46480 29708 46532 29714
rect 46480 29650 46532 29656
rect 44640 29028 44692 29034
rect 44640 28970 44692 28976
rect 46204 29028 46256 29034
rect 46204 28970 46256 28976
rect 44088 28076 44140 28082
rect 44088 28018 44140 28024
rect 44732 28076 44784 28082
rect 44732 28018 44784 28024
rect 44100 27538 44128 28018
rect 44364 27940 44416 27946
rect 44364 27882 44416 27888
rect 44088 27532 44140 27538
rect 44088 27474 44140 27480
rect 43996 27396 44048 27402
rect 43996 27338 44048 27344
rect 44100 27010 44128 27474
rect 44376 27470 44404 27882
rect 44744 27674 44772 28018
rect 44732 27668 44784 27674
rect 44732 27610 44784 27616
rect 44364 27464 44416 27470
rect 44364 27406 44416 27412
rect 44008 26994 44128 27010
rect 43996 26988 44128 26994
rect 44048 26982 44128 26988
rect 44180 26988 44232 26994
rect 43996 26930 44048 26936
rect 44180 26930 44232 26936
rect 44192 26586 44220 26930
rect 44180 26580 44232 26586
rect 44180 26522 44232 26528
rect 43996 26376 44048 26382
rect 43996 26318 44048 26324
rect 44008 26042 44036 26318
rect 43996 26036 44048 26042
rect 43996 25978 44048 25984
rect 43996 25832 44048 25838
rect 43996 25774 44048 25780
rect 44008 24274 44036 25774
rect 44180 24608 44232 24614
rect 44180 24550 44232 24556
rect 43996 24268 44048 24274
rect 43996 24210 44048 24216
rect 44192 24206 44220 24550
rect 44180 24200 44232 24206
rect 44180 24142 44232 24148
rect 44272 24064 44324 24070
rect 44272 24006 44324 24012
rect 43628 23860 43680 23866
rect 43628 23802 43680 23808
rect 44284 23730 44312 24006
rect 43260 23724 43312 23730
rect 43260 23666 43312 23672
rect 44272 23724 44324 23730
rect 44272 23666 44324 23672
rect 42984 23520 43036 23526
rect 42984 23462 43036 23468
rect 42800 22772 42852 22778
rect 42800 22714 42852 22720
rect 42892 22772 42944 22778
rect 42892 22714 42944 22720
rect 42800 22636 42852 22642
rect 42800 22578 42852 22584
rect 41880 22024 41932 22030
rect 41880 21966 41932 21972
rect 42432 22024 42484 22030
rect 42432 21966 42484 21972
rect 42708 22024 42760 22030
rect 42708 21966 42760 21972
rect 41696 21956 41748 21962
rect 41696 21898 41748 21904
rect 41512 20528 41564 20534
rect 41512 20470 41564 20476
rect 41696 20528 41748 20534
rect 41696 20470 41748 20476
rect 41328 20392 41380 20398
rect 41328 20334 41380 20340
rect 41340 19854 41368 20334
rect 41708 19854 41736 20470
rect 41892 20466 41920 21966
rect 42720 21010 42748 21966
rect 42812 21690 42840 22578
rect 42892 22500 42944 22506
rect 42892 22442 42944 22448
rect 42904 22234 42932 22442
rect 42892 22228 42944 22234
rect 42892 22170 42944 22176
rect 42800 21684 42852 21690
rect 42800 21626 42852 21632
rect 42892 21480 42944 21486
rect 42892 21422 42944 21428
rect 42800 21344 42852 21350
rect 42800 21286 42852 21292
rect 42708 21004 42760 21010
rect 42708 20946 42760 20952
rect 41880 20460 41932 20466
rect 41880 20402 41932 20408
rect 41788 19916 41840 19922
rect 41788 19858 41840 19864
rect 41328 19848 41380 19854
rect 41328 19790 41380 19796
rect 41696 19848 41748 19854
rect 41696 19790 41748 19796
rect 41340 19530 41368 19790
rect 41156 19502 41368 19530
rect 40960 19372 41012 19378
rect 41012 19332 41092 19360
rect 40960 19314 41012 19320
rect 40868 19168 40920 19174
rect 40868 19110 40920 19116
rect 40776 18964 40828 18970
rect 40604 18924 40724 18952
rect 40590 18728 40646 18737
rect 40590 18663 40592 18672
rect 40644 18663 40646 18672
rect 40592 18634 40644 18640
rect 40408 18420 40460 18426
rect 40408 18362 40460 18368
rect 40696 18086 40724 18924
rect 40776 18906 40828 18912
rect 40684 18080 40736 18086
rect 40684 18022 40736 18028
rect 40316 17672 40368 17678
rect 40316 17614 40368 17620
rect 40132 17536 40184 17542
rect 40132 17478 40184 17484
rect 40144 16998 40172 17478
rect 40132 16992 40184 16998
rect 40132 16934 40184 16940
rect 40040 16652 40092 16658
rect 40040 16594 40092 16600
rect 39948 16448 40000 16454
rect 40052 16402 40080 16594
rect 40144 16590 40172 16934
rect 40224 16788 40276 16794
rect 40224 16730 40276 16736
rect 40132 16584 40184 16590
rect 40132 16526 40184 16532
rect 40000 16396 40080 16402
rect 39948 16390 40080 16396
rect 39960 16374 40080 16390
rect 39960 16046 39988 16374
rect 39948 16040 40000 16046
rect 40000 15988 40080 15994
rect 39948 15982 40080 15988
rect 39960 15966 40080 15982
rect 40052 15502 40080 15966
rect 40144 15502 40172 16526
rect 39856 15496 39908 15502
rect 39856 15438 39908 15444
rect 40040 15496 40092 15502
rect 40040 15438 40092 15444
rect 40132 15496 40184 15502
rect 40132 15438 40184 15444
rect 40236 14414 40264 16730
rect 40328 16250 40356 17614
rect 40408 17196 40460 17202
rect 40408 17138 40460 17144
rect 40316 16244 40368 16250
rect 40316 16186 40368 16192
rect 40316 16108 40368 16114
rect 40316 16050 40368 16056
rect 40328 15366 40356 16050
rect 40420 15910 40448 17138
rect 40696 16522 40724 18022
rect 40960 17604 41012 17610
rect 40960 17546 41012 17552
rect 40972 17202 41000 17546
rect 40960 17196 41012 17202
rect 40960 17138 41012 17144
rect 40684 16516 40736 16522
rect 40684 16458 40736 16464
rect 40408 15904 40460 15910
rect 40408 15846 40460 15852
rect 40408 15632 40460 15638
rect 40408 15574 40460 15580
rect 40316 15360 40368 15366
rect 40316 15302 40368 15308
rect 40420 14958 40448 15574
rect 40408 14952 40460 14958
rect 40408 14894 40460 14900
rect 40224 14408 40276 14414
rect 40224 14350 40276 14356
rect 40236 12850 40264 14350
rect 40500 14340 40552 14346
rect 40500 14282 40552 14288
rect 40512 14074 40540 14282
rect 40696 14278 40724 16458
rect 41064 16182 41092 19332
rect 41156 18290 41184 19502
rect 41800 19378 41828 19858
rect 41788 19372 41840 19378
rect 41788 19314 41840 19320
rect 41236 19168 41288 19174
rect 41236 19110 41288 19116
rect 41604 19168 41656 19174
rect 41604 19110 41656 19116
rect 41248 18766 41276 19110
rect 41236 18760 41288 18766
rect 41236 18702 41288 18708
rect 41420 18760 41472 18766
rect 41420 18702 41472 18708
rect 41144 18284 41196 18290
rect 41144 18226 41196 18232
rect 41328 18080 41380 18086
rect 41328 18022 41380 18028
rect 41340 17678 41368 18022
rect 41328 17672 41380 17678
rect 41328 17614 41380 17620
rect 41144 17536 41196 17542
rect 41144 17478 41196 17484
rect 41052 16176 41104 16182
rect 41052 16118 41104 16124
rect 40960 15904 41012 15910
rect 40960 15846 41012 15852
rect 40972 14958 41000 15846
rect 40960 14952 41012 14958
rect 40960 14894 41012 14900
rect 40868 14816 40920 14822
rect 40868 14758 40920 14764
rect 40684 14272 40736 14278
rect 40684 14214 40736 14220
rect 40500 14068 40552 14074
rect 40500 14010 40552 14016
rect 40696 13938 40724 14214
rect 40880 14006 40908 14758
rect 40972 14618 41000 14894
rect 41156 14890 41184 17478
rect 41432 17202 41460 18702
rect 41616 18358 41644 19110
rect 41800 18970 41828 19314
rect 41788 18964 41840 18970
rect 41788 18906 41840 18912
rect 41892 18737 41920 20402
rect 41878 18728 41934 18737
rect 41878 18663 41880 18672
rect 41932 18663 41934 18672
rect 41880 18634 41932 18640
rect 41892 18603 41920 18634
rect 41604 18352 41656 18358
rect 41604 18294 41656 18300
rect 41616 17610 41644 18294
rect 41604 17604 41656 17610
rect 41604 17546 41656 17552
rect 41512 17536 41564 17542
rect 41512 17478 41564 17484
rect 41420 17196 41472 17202
rect 41420 17138 41472 17144
rect 41432 16998 41460 17138
rect 41420 16992 41472 16998
rect 41420 16934 41472 16940
rect 41524 16658 41552 17478
rect 41788 17060 41840 17066
rect 41788 17002 41840 17008
rect 41512 16652 41564 16658
rect 41512 16594 41564 16600
rect 41800 16590 41828 17002
rect 42340 16652 42392 16658
rect 42340 16594 42392 16600
rect 41788 16584 41840 16590
rect 41788 16526 41840 16532
rect 42248 16584 42300 16590
rect 42248 16526 42300 16532
rect 42260 15978 42288 16526
rect 42352 16250 42380 16594
rect 42812 16454 42840 21286
rect 42904 18902 42932 21422
rect 42892 18896 42944 18902
rect 42892 18838 42944 18844
rect 42892 18760 42944 18766
rect 42892 18702 42944 18708
rect 42800 16448 42852 16454
rect 42800 16390 42852 16396
rect 42340 16244 42392 16250
rect 42340 16186 42392 16192
rect 42248 15972 42300 15978
rect 42248 15914 42300 15920
rect 42260 15502 42288 15914
rect 42248 15496 42300 15502
rect 42248 15438 42300 15444
rect 42352 15434 42380 16186
rect 42904 16114 42932 18702
rect 42996 17202 43024 23462
rect 43260 23248 43312 23254
rect 43260 23190 43312 23196
rect 43168 23180 43220 23186
rect 43168 23122 43220 23128
rect 43076 23044 43128 23050
rect 43076 22986 43128 22992
rect 43088 22030 43116 22986
rect 43180 22234 43208 23122
rect 43272 22438 43300 23190
rect 43444 23112 43496 23118
rect 43444 23054 43496 23060
rect 43456 22506 43484 23054
rect 44180 22704 44232 22710
rect 44180 22646 44232 22652
rect 43904 22636 43956 22642
rect 43904 22578 43956 22584
rect 43444 22500 43496 22506
rect 43444 22442 43496 22448
rect 43260 22432 43312 22438
rect 43260 22374 43312 22380
rect 43168 22228 43220 22234
rect 43168 22170 43220 22176
rect 43180 22098 43208 22170
rect 43168 22092 43220 22098
rect 43168 22034 43220 22040
rect 43076 22024 43128 22030
rect 43076 21966 43128 21972
rect 43088 21486 43116 21966
rect 43076 21480 43128 21486
rect 43076 21422 43128 21428
rect 43272 21350 43300 22374
rect 43352 22228 43404 22234
rect 43352 22170 43404 22176
rect 43364 21962 43392 22170
rect 43456 22166 43484 22442
rect 43916 22234 43944 22578
rect 44192 22234 44220 22646
rect 44272 22432 44324 22438
rect 44272 22374 44324 22380
rect 44284 22234 44312 22374
rect 43904 22228 43956 22234
rect 43904 22170 43956 22176
rect 44180 22228 44232 22234
rect 44180 22170 44232 22176
rect 44272 22228 44324 22234
rect 44272 22170 44324 22176
rect 43444 22160 43496 22166
rect 43444 22102 43496 22108
rect 44376 22094 44404 27406
rect 45284 26784 45336 26790
rect 45284 26726 45336 26732
rect 45192 25900 45244 25906
rect 45192 25842 45244 25848
rect 44456 25832 44508 25838
rect 44456 25774 44508 25780
rect 44468 25498 44496 25774
rect 45204 25498 45232 25842
rect 45296 25838 45324 26726
rect 45284 25832 45336 25838
rect 45284 25774 45336 25780
rect 44456 25492 44508 25498
rect 44456 25434 44508 25440
rect 45192 25492 45244 25498
rect 45192 25434 45244 25440
rect 45560 25220 45612 25226
rect 45560 25162 45612 25168
rect 45572 24954 45600 25162
rect 45560 24948 45612 24954
rect 45560 24890 45612 24896
rect 44548 24812 44600 24818
rect 44548 24754 44600 24760
rect 44560 23866 44588 24754
rect 45560 24608 45612 24614
rect 45560 24550 45612 24556
rect 45572 23905 45600 24550
rect 45558 23896 45614 23905
rect 44548 23860 44600 23866
rect 45558 23831 45614 23840
rect 44548 23802 44600 23808
rect 44192 22066 44404 22094
rect 43352 21956 43404 21962
rect 43352 21898 43404 21904
rect 43364 21690 43392 21898
rect 43628 21888 43680 21894
rect 43628 21830 43680 21836
rect 43352 21684 43404 21690
rect 43352 21626 43404 21632
rect 43640 21554 43668 21830
rect 43628 21548 43680 21554
rect 43628 21490 43680 21496
rect 43996 21412 44048 21418
rect 43996 21354 44048 21360
rect 43260 21344 43312 21350
rect 43260 21286 43312 21292
rect 43720 20868 43772 20874
rect 43720 20810 43772 20816
rect 43732 20602 43760 20810
rect 43720 20596 43772 20602
rect 43720 20538 43772 20544
rect 43904 20392 43956 20398
rect 43904 20334 43956 20340
rect 43916 19514 43944 20334
rect 44008 19922 44036 21354
rect 44192 20466 44220 22066
rect 44640 21548 44692 21554
rect 44640 21490 44692 21496
rect 44456 21412 44508 21418
rect 44456 21354 44508 21360
rect 44468 20806 44496 21354
rect 44456 20800 44508 20806
rect 44456 20742 44508 20748
rect 44088 20460 44140 20466
rect 44088 20402 44140 20408
rect 44180 20460 44232 20466
rect 44180 20402 44232 20408
rect 44100 20058 44128 20402
rect 44468 20398 44496 20742
rect 44456 20392 44508 20398
rect 44456 20334 44508 20340
rect 44088 20052 44140 20058
rect 44088 19994 44140 20000
rect 43996 19916 44048 19922
rect 43996 19858 44048 19864
rect 43904 19508 43956 19514
rect 43904 19450 43956 19456
rect 44008 19446 44036 19858
rect 44364 19848 44416 19854
rect 44364 19790 44416 19796
rect 44272 19780 44324 19786
rect 44272 19722 44324 19728
rect 43996 19440 44048 19446
rect 43996 19382 44048 19388
rect 44284 19378 44312 19722
rect 44376 19378 44404 19790
rect 43444 19372 43496 19378
rect 43444 19314 43496 19320
rect 44272 19372 44324 19378
rect 44272 19314 44324 19320
rect 44364 19372 44416 19378
rect 44364 19314 44416 19320
rect 43456 18630 43484 19314
rect 44180 19168 44232 19174
rect 44180 19110 44232 19116
rect 43444 18624 43496 18630
rect 43444 18566 43496 18572
rect 43904 18624 43956 18630
rect 43904 18566 43956 18572
rect 43916 18290 43944 18566
rect 43904 18284 43956 18290
rect 43904 18226 43956 18232
rect 43916 18086 43944 18226
rect 43904 18080 43956 18086
rect 43904 18022 43956 18028
rect 43720 17672 43772 17678
rect 43720 17614 43772 17620
rect 43352 17536 43404 17542
rect 43352 17478 43404 17484
rect 42984 17196 43036 17202
rect 42984 17138 43036 17144
rect 42892 16108 42944 16114
rect 42892 16050 42944 16056
rect 42340 15428 42392 15434
rect 42340 15370 42392 15376
rect 41144 14884 41196 14890
rect 41144 14826 41196 14832
rect 40960 14612 41012 14618
rect 40960 14554 41012 14560
rect 40868 14000 40920 14006
rect 40868 13942 40920 13948
rect 40972 13938 41000 14554
rect 40684 13932 40736 13938
rect 40684 13874 40736 13880
rect 40960 13932 41012 13938
rect 40960 13874 41012 13880
rect 42352 12986 42380 15370
rect 42904 15026 42932 16050
rect 42996 15570 43024 17138
rect 43364 16998 43392 17478
rect 43732 17134 43760 17614
rect 43444 17128 43496 17134
rect 43444 17070 43496 17076
rect 43720 17128 43772 17134
rect 43720 17070 43772 17076
rect 43352 16992 43404 16998
rect 43352 16934 43404 16940
rect 43456 16794 43484 17070
rect 43444 16788 43496 16794
rect 43444 16730 43496 16736
rect 43076 16584 43128 16590
rect 43076 16526 43128 16532
rect 43260 16584 43312 16590
rect 43260 16526 43312 16532
rect 43088 16250 43116 16526
rect 43076 16244 43128 16250
rect 43076 16186 43128 16192
rect 43272 15706 43300 16526
rect 43260 15700 43312 15706
rect 43260 15642 43312 15648
rect 42984 15564 43036 15570
rect 42984 15506 43036 15512
rect 42892 15020 42944 15026
rect 42892 14962 42944 14968
rect 42996 13938 43024 15506
rect 43260 15496 43312 15502
rect 43260 15438 43312 15444
rect 43352 15496 43404 15502
rect 43352 15438 43404 15444
rect 43272 15094 43300 15438
rect 43260 15088 43312 15094
rect 43260 15030 43312 15036
rect 43364 14958 43392 15438
rect 44192 15434 44220 19110
rect 44284 18834 44312 19314
rect 44376 18834 44404 19314
rect 44272 18828 44324 18834
rect 44272 18770 44324 18776
rect 44364 18828 44416 18834
rect 44364 18770 44416 18776
rect 44376 18426 44404 18770
rect 44364 18420 44416 18426
rect 44364 18362 44416 18368
rect 44272 18352 44324 18358
rect 44468 18306 44496 20334
rect 44652 19378 44680 21490
rect 46216 20466 46244 28970
rect 46480 28960 46532 28966
rect 46480 28902 46532 28908
rect 46492 28626 46520 28902
rect 46480 28620 46532 28626
rect 46480 28562 46532 28568
rect 46480 27872 46532 27878
rect 46480 27814 46532 27820
rect 46492 26450 46520 27814
rect 46768 26994 46796 32982
rect 46846 27976 46902 27985
rect 46846 27911 46902 27920
rect 46860 27538 46888 27911
rect 46848 27532 46900 27538
rect 46848 27474 46900 27480
rect 46756 26988 46808 26994
rect 46756 26930 46808 26936
rect 46664 26784 46716 26790
rect 46664 26726 46716 26732
rect 46676 26450 46704 26726
rect 46846 26616 46902 26625
rect 46846 26551 46902 26560
rect 46480 26444 46532 26450
rect 46480 26386 46532 26392
rect 46664 26444 46716 26450
rect 46664 26386 46716 26392
rect 46754 25936 46810 25945
rect 46754 25871 46810 25880
rect 46768 25838 46796 25871
rect 46756 25832 46808 25838
rect 46756 25774 46808 25780
rect 46860 25362 46888 26551
rect 46848 25356 46900 25362
rect 46848 25298 46900 25304
rect 46480 24200 46532 24206
rect 46480 24142 46532 24148
rect 46492 23730 46520 24142
rect 46480 23724 46532 23730
rect 46480 23666 46532 23672
rect 46846 22536 46902 22545
rect 46846 22471 46902 22480
rect 46860 22098 46888 22471
rect 46848 22092 46900 22098
rect 46848 22034 46900 22040
rect 46388 21548 46440 21554
rect 46388 21490 46440 21496
rect 45652 20460 45704 20466
rect 45652 20402 45704 20408
rect 46204 20460 46256 20466
rect 46204 20402 46256 20408
rect 44640 19372 44692 19378
rect 44640 19314 44692 19320
rect 44548 19304 44600 19310
rect 44548 19246 44600 19252
rect 44560 18902 44588 19246
rect 44548 18896 44600 18902
rect 44548 18838 44600 18844
rect 44560 18698 44588 18838
rect 44652 18766 44680 19314
rect 45468 18896 45520 18902
rect 45468 18838 45520 18844
rect 44640 18760 44692 18766
rect 44640 18702 44692 18708
rect 45376 18760 45428 18766
rect 45376 18702 45428 18708
rect 44548 18692 44600 18698
rect 44548 18634 44600 18640
rect 44272 18294 44324 18300
rect 44284 17610 44312 18294
rect 44376 18278 44496 18306
rect 44376 17814 44404 18278
rect 44560 17882 44588 18634
rect 45192 18624 45244 18630
rect 45192 18566 45244 18572
rect 45204 18358 45232 18566
rect 45192 18352 45244 18358
rect 45192 18294 45244 18300
rect 44640 18080 44692 18086
rect 44640 18022 44692 18028
rect 44548 17876 44600 17882
rect 44548 17818 44600 17824
rect 44364 17808 44416 17814
rect 44364 17750 44416 17756
rect 44456 17740 44508 17746
rect 44456 17682 44508 17688
rect 44272 17604 44324 17610
rect 44272 17546 44324 17552
rect 44284 17338 44312 17546
rect 44272 17332 44324 17338
rect 44272 17274 44324 17280
rect 44468 17202 44496 17682
rect 44652 17678 44680 18022
rect 45388 17882 45416 18702
rect 45480 18426 45508 18838
rect 45664 18698 45692 20402
rect 45560 18692 45612 18698
rect 45560 18634 45612 18640
rect 45652 18692 45704 18698
rect 45652 18634 45704 18640
rect 45468 18420 45520 18426
rect 45468 18362 45520 18368
rect 45468 18284 45520 18290
rect 45468 18226 45520 18232
rect 45376 17876 45428 17882
rect 45376 17818 45428 17824
rect 45480 17678 45508 18226
rect 44640 17672 44692 17678
rect 44640 17614 44692 17620
rect 45468 17672 45520 17678
rect 45468 17614 45520 17620
rect 44548 17536 44600 17542
rect 44548 17478 44600 17484
rect 44560 17202 44588 17478
rect 44456 17196 44508 17202
rect 44456 17138 44508 17144
rect 44548 17196 44600 17202
rect 44548 17138 44600 17144
rect 44468 16182 44496 17138
rect 44456 16176 44508 16182
rect 44456 16118 44508 16124
rect 44468 16046 44496 16118
rect 44456 16040 44508 16046
rect 44456 15982 44508 15988
rect 44456 15496 44508 15502
rect 44376 15456 44456 15484
rect 44180 15428 44232 15434
rect 44180 15370 44232 15376
rect 43536 15360 43588 15366
rect 43536 15302 43588 15308
rect 43548 15026 43576 15302
rect 43536 15020 43588 15026
rect 43536 14962 43588 14968
rect 44376 14958 44404 15456
rect 44560 15484 44588 17138
rect 45284 17128 45336 17134
rect 45284 17070 45336 17076
rect 45192 16584 45244 16590
rect 45192 16526 45244 16532
rect 45204 16114 45232 16526
rect 45296 16250 45324 17070
rect 45480 16794 45508 17614
rect 45468 16788 45520 16794
rect 45468 16730 45520 16736
rect 45468 16584 45520 16590
rect 45468 16526 45520 16532
rect 45284 16244 45336 16250
rect 45284 16186 45336 16192
rect 45192 16108 45244 16114
rect 45192 16050 45244 16056
rect 44640 15904 44692 15910
rect 44640 15846 44692 15852
rect 44652 15706 44680 15846
rect 44640 15700 44692 15706
rect 44640 15642 44692 15648
rect 45296 15502 45324 16186
rect 45376 16040 45428 16046
rect 45376 15982 45428 15988
rect 45388 15706 45416 15982
rect 45376 15700 45428 15706
rect 45376 15642 45428 15648
rect 44508 15456 44588 15484
rect 45284 15496 45336 15502
rect 44456 15438 44508 15444
rect 45284 15438 45336 15444
rect 45480 15434 45508 16526
rect 45572 16114 45600 18634
rect 46112 16652 46164 16658
rect 46112 16594 46164 16600
rect 45560 16108 45612 16114
rect 45560 16050 45612 16056
rect 45572 15570 45600 16050
rect 45560 15564 45612 15570
rect 45560 15506 45612 15512
rect 45008 15428 45060 15434
rect 45008 15370 45060 15376
rect 45468 15428 45520 15434
rect 45468 15370 45520 15376
rect 45020 15026 45048 15370
rect 45008 15020 45060 15026
rect 45008 14962 45060 14968
rect 43352 14952 43404 14958
rect 43352 14894 43404 14900
rect 44272 14952 44324 14958
rect 44272 14894 44324 14900
rect 44364 14952 44416 14958
rect 44364 14894 44416 14900
rect 43720 14816 43772 14822
rect 43720 14758 43772 14764
rect 43732 14346 43760 14758
rect 43720 14340 43772 14346
rect 43720 14282 43772 14288
rect 44284 14278 44312 14894
rect 44376 14822 44404 14894
rect 45480 14890 45508 15370
rect 45468 14884 45520 14890
rect 45468 14826 45520 14832
rect 44364 14816 44416 14822
rect 44364 14758 44416 14764
rect 44376 14618 44404 14758
rect 44364 14612 44416 14618
rect 44364 14554 44416 14560
rect 46124 14414 46152 16594
rect 46112 14408 46164 14414
rect 46112 14350 46164 14356
rect 44272 14272 44324 14278
rect 44272 14214 44324 14220
rect 42984 13932 43036 13938
rect 42984 13874 43036 13880
rect 42340 12980 42392 12986
rect 42340 12922 42392 12928
rect 40224 12844 40276 12850
rect 40224 12786 40276 12792
rect 39580 9172 39632 9178
rect 39580 9114 39632 9120
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 43260 7200 43312 7206
rect 43260 7142 43312 7148
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 43272 6866 43300 7142
rect 43260 6860 43312 6866
rect 43260 6802 43312 6808
rect 46112 6792 46164 6798
rect 46112 6734 46164 6740
rect 43076 6724 43128 6730
rect 43076 6666 43128 6672
rect 43088 6458 43116 6666
rect 43076 6452 43128 6458
rect 43076 6394 43128 6400
rect 43076 6316 43128 6322
rect 43076 6258 43128 6264
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 43088 4622 43116 6258
rect 46124 5778 46152 6734
rect 46112 5772 46164 5778
rect 46112 5714 46164 5720
rect 45652 5704 45704 5710
rect 45652 5646 45704 5652
rect 46216 5658 46244 20402
rect 46296 20256 46348 20262
rect 46296 20198 46348 20204
rect 46308 19990 46336 20198
rect 46296 19984 46348 19990
rect 46296 19926 46348 19932
rect 46296 6656 46348 6662
rect 46296 6598 46348 6604
rect 46308 5778 46336 6598
rect 46400 6322 46428 21490
rect 46664 21344 46716 21350
rect 46664 21286 46716 21292
rect 46676 21010 46704 21286
rect 46664 21004 46716 21010
rect 46664 20946 46716 20952
rect 46480 20256 46532 20262
rect 46480 20198 46532 20204
rect 46492 19922 46520 20198
rect 46480 19916 46532 19922
rect 46480 19858 46532 19864
rect 46480 18692 46532 18698
rect 46480 18634 46532 18640
rect 46492 16114 46520 18634
rect 46846 17776 46902 17785
rect 46846 17711 46848 17720
rect 46900 17711 46902 17720
rect 46848 17682 46900 17688
rect 46664 16516 46716 16522
rect 46664 16458 46716 16464
rect 46676 16250 46704 16458
rect 46664 16244 46716 16250
rect 46664 16186 46716 16192
rect 46480 16108 46532 16114
rect 46480 16050 46532 16056
rect 46846 15056 46902 15065
rect 46846 14991 46902 15000
rect 46860 14482 46888 14991
rect 46848 14476 46900 14482
rect 46848 14418 46900 14424
rect 46846 13696 46902 13705
rect 46846 13631 46902 13640
rect 46754 13560 46810 13569
rect 46754 13495 46810 13504
rect 46768 12850 46796 13495
rect 46860 13394 46888 13631
rect 46848 13388 46900 13394
rect 46848 13330 46900 13336
rect 46756 12844 46808 12850
rect 46756 12786 46808 12792
rect 46664 12640 46716 12646
rect 46664 12582 46716 12588
rect 46676 12306 46704 12582
rect 46664 12300 46716 12306
rect 46664 12242 46716 12248
rect 46846 6896 46902 6905
rect 46846 6831 46848 6840
rect 46900 6831 46902 6840
rect 46848 6802 46900 6808
rect 46388 6316 46440 6322
rect 46388 6258 46440 6264
rect 46952 6202 46980 33322
rect 47032 33312 47084 33318
rect 47032 33254 47084 33260
rect 47044 32978 47072 33254
rect 47136 33046 47164 35634
rect 47124 33040 47176 33046
rect 47124 32982 47176 32988
rect 47032 32972 47084 32978
rect 47032 32914 47084 32920
rect 47320 32502 47348 49286
rect 48290 49200 48402 49800
rect 48934 49200 49046 49800
rect 49578 49200 49690 49800
rect 47768 46980 47820 46986
rect 47768 46922 47820 46928
rect 47400 46572 47452 46578
rect 47400 46514 47452 46520
rect 47412 45830 47440 46514
rect 47400 45824 47452 45830
rect 47400 45766 47452 45772
rect 47412 45490 47440 45766
rect 47400 45484 47452 45490
rect 47400 45426 47452 45432
rect 47412 44305 47440 45426
rect 47398 44296 47454 44305
rect 47398 44231 47454 44240
rect 47676 43308 47728 43314
rect 47676 43250 47728 43256
rect 47400 40044 47452 40050
rect 47400 39986 47452 39992
rect 47308 32496 47360 32502
rect 47308 32438 47360 32444
rect 47308 29164 47360 29170
rect 47308 29106 47360 29112
rect 47124 28960 47176 28966
rect 47124 28902 47176 28908
rect 47136 28626 47164 28902
rect 47124 28620 47176 28626
rect 47124 28562 47176 28568
rect 47124 26988 47176 26994
rect 47124 26930 47176 26936
rect 47032 25832 47084 25838
rect 47032 25774 47084 25780
rect 47044 24818 47072 25774
rect 47032 24812 47084 24818
rect 47032 24754 47084 24760
rect 47136 23798 47164 26930
rect 47216 25832 47268 25838
rect 47216 25774 47268 25780
rect 47228 24818 47256 25774
rect 47216 24812 47268 24818
rect 47216 24754 47268 24760
rect 47216 24676 47268 24682
rect 47216 24618 47268 24624
rect 47124 23792 47176 23798
rect 47124 23734 47176 23740
rect 47032 21344 47084 21350
rect 47032 21286 47084 21292
rect 47044 21078 47072 21286
rect 47032 21072 47084 21078
rect 47032 21014 47084 21020
rect 47228 19378 47256 24618
rect 47320 22094 47348 29106
rect 47412 26994 47440 39986
rect 47584 38956 47636 38962
rect 47584 38898 47636 38904
rect 47492 27328 47544 27334
rect 47492 27270 47544 27276
rect 47400 26988 47452 26994
rect 47400 26930 47452 26936
rect 47504 24750 47532 27270
rect 47492 24744 47544 24750
rect 47492 24686 47544 24692
rect 47320 22066 47532 22094
rect 47308 20800 47360 20806
rect 47308 20742 47360 20748
rect 47216 19372 47268 19378
rect 47216 19314 47268 19320
rect 47124 19168 47176 19174
rect 47124 19110 47176 19116
rect 47136 18834 47164 19110
rect 47124 18828 47176 18834
rect 47124 18770 47176 18776
rect 47216 17196 47268 17202
rect 47216 17138 47268 17144
rect 47032 12640 47084 12646
rect 47032 12582 47084 12588
rect 47044 12374 47072 12582
rect 47032 12368 47084 12374
rect 47032 12310 47084 12316
rect 47228 6322 47256 17138
rect 47320 6798 47348 20742
rect 47400 16448 47452 16454
rect 47400 16390 47452 16396
rect 47412 16182 47440 16390
rect 47400 16176 47452 16182
rect 47400 16118 47452 16124
rect 47504 15026 47532 22066
rect 47596 21554 47624 38898
rect 47688 27334 47716 43250
rect 47780 32570 47808 46922
rect 48332 46034 48360 49200
rect 48976 47054 49004 49200
rect 48964 47048 49016 47054
rect 48964 46990 49016 46996
rect 48320 46028 48372 46034
rect 48320 45970 48372 45976
rect 48320 45280 48372 45286
rect 48320 45222 48372 45228
rect 48332 44946 48360 45222
rect 48320 44940 48372 44946
rect 48320 44882 48372 44888
rect 47860 44804 47912 44810
rect 47860 44746 47912 44752
rect 47872 44538 47900 44746
rect 47860 44532 47912 44538
rect 47860 44474 47912 44480
rect 47860 43104 47912 43110
rect 47860 43046 47912 43052
rect 47872 42634 47900 43046
rect 48226 42936 48282 42945
rect 48226 42871 48282 42880
rect 48240 42770 48268 42871
rect 48228 42764 48280 42770
rect 48228 42706 48280 42712
rect 47860 42628 47912 42634
rect 47860 42570 47912 42576
rect 48228 41676 48280 41682
rect 48228 41618 48280 41624
rect 48240 41585 48268 41618
rect 48226 41576 48282 41585
rect 48226 41511 48282 41520
rect 48320 40452 48372 40458
rect 48320 40394 48372 40400
rect 48332 40225 48360 40394
rect 48318 40216 48374 40225
rect 48318 40151 48374 40160
rect 48320 39840 48372 39846
rect 48320 39782 48372 39788
rect 48332 39506 48360 39782
rect 48320 39500 48372 39506
rect 48320 39442 48372 39448
rect 47860 39364 47912 39370
rect 47860 39306 47912 39312
rect 47872 39098 47900 39306
rect 47860 39092 47912 39098
rect 47860 39034 47912 39040
rect 48320 38344 48372 38350
rect 48320 38286 48372 38292
rect 48044 37868 48096 37874
rect 48044 37810 48096 37816
rect 47950 37496 48006 37505
rect 47950 37431 48006 37440
rect 47768 32564 47820 32570
rect 47768 32506 47820 32512
rect 47964 31890 47992 37431
rect 47952 31884 48004 31890
rect 47952 31826 48004 31832
rect 48056 31754 48084 37810
rect 48136 37664 48188 37670
rect 48136 37606 48188 37612
rect 48148 37330 48176 37606
rect 48136 37324 48188 37330
rect 48136 37266 48188 37272
rect 48332 37262 48360 38286
rect 48320 37256 48372 37262
rect 48320 37198 48372 37204
rect 48320 36576 48372 36582
rect 48320 36518 48372 36524
rect 48332 36242 48360 36518
rect 48320 36236 48372 36242
rect 48320 36178 48372 36184
rect 48136 36100 48188 36106
rect 48136 36042 48188 36048
rect 48148 35834 48176 36042
rect 48136 35828 48188 35834
rect 48136 35770 48188 35776
rect 48320 32836 48372 32842
rect 48320 32778 48372 32784
rect 48332 32745 48360 32778
rect 48318 32736 48374 32745
rect 48318 32671 48374 32680
rect 47964 31726 48084 31754
rect 47766 30288 47822 30297
rect 47766 30223 47768 30232
rect 47820 30223 47822 30232
rect 47768 30194 47820 30200
rect 47780 28082 47808 30194
rect 47860 30048 47912 30054
rect 47860 29990 47912 29996
rect 47872 29714 47900 29990
rect 47860 29708 47912 29714
rect 47860 29650 47912 29656
rect 47768 28076 47820 28082
rect 47768 28018 47820 28024
rect 47780 27849 47808 28018
rect 47766 27840 47822 27849
rect 47766 27775 47822 27784
rect 47676 27328 47728 27334
rect 47676 27270 47728 27276
rect 47964 27146 47992 31726
rect 48320 29572 48372 29578
rect 48320 29514 48372 29520
rect 48332 29345 48360 29514
rect 48318 29336 48374 29345
rect 48318 29271 48374 29280
rect 48320 29028 48372 29034
rect 48320 28970 48372 28976
rect 48226 28656 48282 28665
rect 48226 28591 48228 28600
rect 48280 28591 48282 28600
rect 48228 28562 48280 28568
rect 48136 27872 48188 27878
rect 48136 27814 48188 27820
rect 48148 27538 48176 27814
rect 48332 27538 48360 28970
rect 48136 27532 48188 27538
rect 48136 27474 48188 27480
rect 48320 27532 48372 27538
rect 48320 27474 48372 27480
rect 47688 27118 47992 27146
rect 47584 21548 47636 21554
rect 47584 21490 47636 21496
rect 47584 19372 47636 19378
rect 47584 19314 47636 19320
rect 47596 17082 47624 19314
rect 47688 17202 47716 27118
rect 47768 26988 47820 26994
rect 47768 26930 47820 26936
rect 47780 21554 47808 26930
rect 48136 26784 48188 26790
rect 48136 26726 48188 26732
rect 47952 26444 48004 26450
rect 47952 26386 48004 26392
rect 47860 24132 47912 24138
rect 47860 24074 47912 24080
rect 47872 23866 47900 24074
rect 47860 23860 47912 23866
rect 47860 23802 47912 23808
rect 47860 21956 47912 21962
rect 47860 21898 47912 21904
rect 47872 21690 47900 21898
rect 47860 21684 47912 21690
rect 47860 21626 47912 21632
rect 47768 21548 47820 21554
rect 47768 21490 47820 21496
rect 47780 20806 47808 21490
rect 47768 20800 47820 20806
rect 47768 20742 47820 20748
rect 47768 19168 47820 19174
rect 47768 19110 47820 19116
rect 47780 18902 47808 19110
rect 47768 18896 47820 18902
rect 47768 18838 47820 18844
rect 47860 17604 47912 17610
rect 47860 17546 47912 17552
rect 47872 17338 47900 17546
rect 47860 17332 47912 17338
rect 47860 17274 47912 17280
rect 47676 17196 47728 17202
rect 47676 17138 47728 17144
rect 47596 17054 47808 17082
rect 47492 15020 47544 15026
rect 47492 14962 47544 14968
rect 47504 12850 47532 14962
rect 47492 12844 47544 12850
rect 47492 12786 47544 12792
rect 47676 12844 47728 12850
rect 47676 12786 47728 12792
rect 47688 6798 47716 12786
rect 47308 6792 47360 6798
rect 47308 6734 47360 6740
rect 47676 6792 47728 6798
rect 47676 6734 47728 6740
rect 47320 6390 47348 6734
rect 47584 6656 47636 6662
rect 47584 6598 47636 6604
rect 47308 6384 47360 6390
rect 47308 6326 47360 6332
rect 47216 6316 47268 6322
rect 47216 6258 47268 6264
rect 46860 6174 46980 6202
rect 47308 6248 47360 6254
rect 47308 6190 47360 6196
rect 46860 5846 46888 6174
rect 46940 6112 46992 6118
rect 46940 6054 46992 6060
rect 47032 6112 47084 6118
rect 47032 6054 47084 6060
rect 46848 5840 46900 5846
rect 46848 5782 46900 5788
rect 46296 5772 46348 5778
rect 46296 5714 46348 5720
rect 45560 5568 45612 5574
rect 45560 5510 45612 5516
rect 44732 5024 44784 5030
rect 44732 4966 44784 4972
rect 39028 4616 39080 4622
rect 39028 4558 39080 4564
rect 43076 4616 43128 4622
rect 43076 4558 43128 4564
rect 44364 4616 44416 4622
rect 44364 4558 44416 4564
rect 44548 4616 44600 4622
rect 44548 4558 44600 4564
rect 39040 4146 39068 4558
rect 38384 4140 38436 4146
rect 38384 4082 38436 4088
rect 39028 4140 39080 4146
rect 39028 4082 39080 4088
rect 41972 4140 42024 4146
rect 41972 4082 42024 4088
rect 38200 4072 38252 4078
rect 38200 4014 38252 4020
rect 38108 4004 38160 4010
rect 38108 3946 38160 3952
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34060 3596 34112 3602
rect 34060 3538 34112 3544
rect 38120 3534 38148 3946
rect 38212 3670 38240 4014
rect 38396 4010 38424 4082
rect 40500 4072 40552 4078
rect 40500 4014 40552 4020
rect 38384 4004 38436 4010
rect 38384 3946 38436 3952
rect 38200 3664 38252 3670
rect 38200 3606 38252 3612
rect 38108 3528 38160 3534
rect 38108 3470 38160 3476
rect 33324 3460 33376 3466
rect 33324 3402 33376 3408
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 38396 2446 38424 3946
rect 38936 3936 38988 3942
rect 38936 3878 38988 3884
rect 38752 3528 38804 3534
rect 38752 3470 38804 3476
rect 38764 3058 38792 3470
rect 38948 3126 38976 3878
rect 38936 3120 38988 3126
rect 38936 3062 38988 3068
rect 38752 3052 38804 3058
rect 38752 2994 38804 3000
rect 39304 2984 39356 2990
rect 39304 2926 39356 2932
rect 38384 2440 38436 2446
rect 38384 2382 38436 2388
rect 38660 2372 38712 2378
rect 38660 2314 38712 2320
rect 38672 800 38700 2314
rect 39316 800 39344 2926
rect 40512 2258 40540 4014
rect 40776 3936 40828 3942
rect 40776 3878 40828 3884
rect 40788 3602 40816 3878
rect 40776 3596 40828 3602
rect 40776 3538 40828 3544
rect 41236 3596 41288 3602
rect 41236 3538 41288 3544
rect 40592 3528 40644 3534
rect 40592 3470 40644 3476
rect 40604 3058 40632 3470
rect 40592 3052 40644 3058
rect 40592 2994 40644 3000
rect 40512 2230 40632 2258
rect 40604 800 40632 2230
rect 41248 800 41276 3538
rect 41984 3534 42012 4082
rect 43088 3738 43116 4558
rect 44180 4072 44232 4078
rect 44180 4014 44232 4020
rect 44088 4004 44140 4010
rect 44088 3946 44140 3952
rect 44100 3738 44128 3946
rect 43076 3732 43128 3738
rect 43076 3674 43128 3680
rect 44088 3732 44140 3738
rect 44088 3674 44140 3680
rect 41972 3528 42024 3534
rect 41972 3470 42024 3476
rect 43812 3460 43864 3466
rect 43812 3402 43864 3408
rect 42800 3392 42852 3398
rect 42800 3334 42852 3340
rect 42812 3126 42840 3334
rect 42800 3120 42852 3126
rect 42800 3062 42852 3068
rect 41880 2848 41932 2854
rect 41880 2790 41932 2796
rect 41892 800 41920 2790
rect 43824 800 43852 3402
rect 44192 2106 44220 4014
rect 44376 3058 44404 4558
rect 44560 3602 44588 4558
rect 44548 3596 44600 3602
rect 44548 3538 44600 3544
rect 44364 3052 44416 3058
rect 44364 2994 44416 3000
rect 44744 2514 44772 4966
rect 45100 4480 45152 4486
rect 45100 4422 45152 4428
rect 45376 4480 45428 4486
rect 45376 4422 45428 4428
rect 45112 3126 45140 4422
rect 45284 3664 45336 3670
rect 45284 3606 45336 3612
rect 45100 3120 45152 3126
rect 45100 3062 45152 3068
rect 44732 2508 44784 2514
rect 44732 2450 44784 2456
rect 44180 2100 44232 2106
rect 44180 2042 44232 2048
rect 45296 1986 45324 3606
rect 45388 3602 45416 4422
rect 45376 3596 45428 3602
rect 45376 3538 45428 3544
rect 45572 2378 45600 5510
rect 45664 3466 45692 5646
rect 46216 5630 46336 5658
rect 45744 4072 45796 4078
rect 45744 4014 45796 4020
rect 45652 3460 45704 3466
rect 45652 3402 45704 3408
rect 45560 2372 45612 2378
rect 45560 2314 45612 2320
rect 45112 1958 45324 1986
rect 45112 800 45140 1958
rect 45756 800 45784 4014
rect 46308 3058 46336 5630
rect 46846 5536 46902 5545
rect 46846 5471 46902 5480
rect 46860 4690 46888 5471
rect 46848 4684 46900 4690
rect 46848 4626 46900 4632
rect 46756 4616 46808 4622
rect 46756 4558 46808 4564
rect 46768 4146 46796 4558
rect 46756 4140 46808 4146
rect 46756 4082 46808 4088
rect 46296 3052 46348 3058
rect 46296 2994 46348 3000
rect 46756 2984 46808 2990
rect 46756 2926 46808 2932
rect 46768 1465 46796 2926
rect 46952 2378 46980 6054
rect 47044 5302 47072 6054
rect 47124 5772 47176 5778
rect 47124 5714 47176 5720
rect 47032 5296 47084 5302
rect 47032 5238 47084 5244
rect 47136 2774 47164 5714
rect 47216 5160 47268 5166
rect 47216 5102 47268 5108
rect 47228 4146 47256 5102
rect 47216 4140 47268 4146
rect 47216 4082 47268 4088
rect 47320 3738 47348 6190
rect 47596 4010 47624 6598
rect 47780 6322 47808 17054
rect 47860 13252 47912 13258
rect 47860 13194 47912 13200
rect 47872 12986 47900 13194
rect 47860 12980 47912 12986
rect 47860 12922 47912 12928
rect 47964 12345 47992 26386
rect 48148 25362 48176 26726
rect 48320 25696 48372 25702
rect 48320 25638 48372 25644
rect 48332 25362 48360 25638
rect 48136 25356 48188 25362
rect 48136 25298 48188 25304
rect 48320 25356 48372 25362
rect 48320 25298 48372 25304
rect 48228 24812 48280 24818
rect 48228 24754 48280 24760
rect 48044 24676 48096 24682
rect 48044 24618 48096 24624
rect 48056 23322 48084 24618
rect 48240 24585 48268 24754
rect 48226 24576 48282 24585
rect 48226 24511 48282 24520
rect 48136 24268 48188 24274
rect 48136 24210 48188 24216
rect 48044 23316 48096 23322
rect 48044 23258 48096 23264
rect 48148 17105 48176 24210
rect 48320 22432 48372 22438
rect 48320 22374 48372 22380
rect 48332 22098 48360 22374
rect 48320 22092 48372 22098
rect 48320 22034 48372 22040
rect 48226 21856 48282 21865
rect 48226 21791 48282 21800
rect 48240 21010 48268 21791
rect 48228 21004 48280 21010
rect 48228 20946 48280 20952
rect 48226 20496 48282 20505
rect 48226 20431 48282 20440
rect 48240 19922 48268 20431
rect 48228 19916 48280 19922
rect 48228 19858 48280 19864
rect 48226 19136 48282 19145
rect 48226 19071 48282 19080
rect 48240 18834 48268 19071
rect 48228 18828 48280 18834
rect 48228 18770 48280 18776
rect 48320 18080 48372 18086
rect 48320 18022 48372 18028
rect 48332 17746 48360 18022
rect 48320 17740 48372 17746
rect 48320 17682 48372 17688
rect 48134 17096 48190 17105
rect 48134 17031 48190 17040
rect 48320 15496 48372 15502
rect 48320 15438 48372 15444
rect 48136 14816 48188 14822
rect 48136 14758 48188 14764
rect 48148 14482 48176 14758
rect 48332 14482 48360 15438
rect 48136 14476 48188 14482
rect 48136 14418 48188 14424
rect 48320 14476 48372 14482
rect 48320 14418 48372 14424
rect 48320 13864 48372 13870
rect 48320 13806 48372 13812
rect 48332 13394 48360 13806
rect 48320 13388 48372 13394
rect 48320 13330 48372 13336
rect 48226 13016 48282 13025
rect 48226 12951 48282 12960
rect 47950 12336 48006 12345
rect 48240 12306 48268 12951
rect 47950 12271 48006 12280
rect 48228 12300 48280 12306
rect 48228 12242 48280 12248
rect 48226 8936 48282 8945
rect 48226 8871 48228 8880
rect 48280 8871 48282 8880
rect 48228 8842 48280 8848
rect 48228 8492 48280 8498
rect 48228 8434 48280 8440
rect 48240 8265 48268 8434
rect 48226 8256 48282 8265
rect 48226 8191 48282 8200
rect 47952 6792 48004 6798
rect 47952 6734 48004 6740
rect 47768 6316 47820 6322
rect 47768 6258 47820 6264
rect 47780 4758 47808 6258
rect 47768 4752 47820 4758
rect 47768 4694 47820 4700
rect 47860 4072 47912 4078
rect 47860 4014 47912 4020
rect 47584 4004 47636 4010
rect 47584 3946 47636 3952
rect 47308 3732 47360 3738
rect 47308 3674 47360 3680
rect 47872 3194 47900 4014
rect 47964 3942 47992 6734
rect 48136 6112 48188 6118
rect 48136 6054 48188 6060
rect 48148 4690 48176 6054
rect 48412 5092 48464 5098
rect 48412 5034 48464 5040
rect 48320 5024 48372 5030
rect 48320 4966 48372 4972
rect 48332 4690 48360 4966
rect 48136 4684 48188 4690
rect 48136 4626 48188 4632
rect 48320 4684 48372 4690
rect 48320 4626 48372 4632
rect 47952 3936 48004 3942
rect 47952 3878 48004 3884
rect 48320 3528 48372 3534
rect 48318 3496 48320 3505
rect 48372 3496 48374 3505
rect 48318 3431 48374 3440
rect 47860 3188 47912 3194
rect 47860 3130 47912 3136
rect 47044 2746 47164 2774
rect 46940 2372 46992 2378
rect 46940 2314 46992 2320
rect 46846 2136 46902 2145
rect 46846 2071 46848 2080
rect 46900 2071 46902 2080
rect 46848 2042 46900 2048
rect 46754 1456 46810 1465
rect 46754 1391 46810 1400
rect 47044 800 47072 2746
rect 47676 2508 47728 2514
rect 47676 2450 47728 2456
rect 47688 800 47716 2450
rect 22756 734 22968 762
rect 23818 200 23930 800
rect 24462 200 24574 800
rect 25750 200 25862 800
rect 26394 200 26506 800
rect 27682 200 27794 800
rect 28326 200 28438 800
rect 28970 200 29082 800
rect 30258 200 30370 800
rect 30902 200 31014 800
rect 32190 200 32302 800
rect 32834 200 32946 800
rect 34122 200 34234 800
rect 34766 200 34878 800
rect 35410 200 35522 800
rect 36698 200 36810 800
rect 37342 200 37454 800
rect 38630 200 38742 800
rect 39274 200 39386 800
rect 40562 200 40674 800
rect 41206 200 41318 800
rect 41850 200 41962 800
rect 43138 200 43250 800
rect 43782 200 43894 800
rect 45070 200 45182 800
rect 45714 200 45826 800
rect 47002 200 47114 800
rect 47646 200 47758 800
rect 48424 105 48452 5034
rect 48964 2576 49016 2582
rect 48964 2518 49016 2524
rect 48976 800 49004 2518
rect 48934 200 49046 800
rect 49578 200 49690 800
rect 48410 96 48466 105
rect 48410 31 48466 40
<< via2 >>
rect 2870 48320 2926 48376
rect 2778 47640 2834 47696
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4066 46280 4122 46336
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 3146 45600 3202 45656
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 2778 43560 2834 43616
rect 1674 38800 1730 38856
rect 1674 36760 1730 36816
rect 1582 34040 1638 34096
rect 1582 32000 1638 32056
rect 1582 25236 1584 25256
rect 1584 25236 1636 25256
rect 1636 25236 1638 25256
rect 1582 25200 1638 25236
rect 1582 21800 1638 21856
rect 3054 41540 3110 41576
rect 3054 41520 3056 41540
rect 3056 41520 3108 41540
rect 3108 41520 3110 41540
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 3238 40840 3294 40896
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4066 32680 4122 32736
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 2778 20440 2834 20496
rect 2778 18400 2834 18456
rect 1582 14356 1584 14376
rect 1584 14356 1636 14376
rect 1636 14356 1638 14376
rect 1582 14320 1638 14356
rect 1582 10240 1638 10296
rect 1582 7520 1638 7576
rect 1582 6860 1638 6896
rect 1582 6840 1584 6860
rect 1584 6840 1636 6860
rect 1636 6840 1638 6860
rect 2870 17076 2872 17096
rect 2872 17076 2924 17096
rect 2924 17076 2926 17096
rect 2870 17040 2926 17076
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 3330 23840 3386 23896
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 2778 11636 2780 11656
rect 2780 11636 2832 11656
rect 2832 11636 2834 11656
rect 2778 11600 2834 11636
rect 2962 9560 3018 9616
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 3422 15036 3424 15056
rect 3424 15036 3476 15056
rect 3476 15036 3478 15056
rect 3422 15000 3478 15036
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 1582 5480 1638 5536
rect 2778 4800 2834 4856
rect 1582 3476 1584 3496
rect 1584 3476 1636 3496
rect 1636 3476 1638 3496
rect 1582 3440 1638 3476
rect 1582 2760 1638 2816
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 2870 1400 2926 1456
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 16670 20304 16726 20360
rect 17038 20460 17094 20496
rect 17038 20440 17040 20460
rect 17040 20440 17092 20460
rect 17092 20440 17094 20460
rect 17958 20304 18014 20360
rect 18142 20460 18198 20496
rect 18142 20440 18144 20460
rect 18144 20440 18196 20460
rect 18196 20440 18198 20460
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 25962 31592 26018 31648
rect 22098 19216 22154 19272
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 2778 720 2834 776
rect 25594 26152 25650 26208
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 27158 22072 27214 22128
rect 27434 22072 27490 22128
rect 27710 19216 27766 19272
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34334 30252 34390 30288
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34334 30232 34336 30252
rect 34336 30232 34388 30252
rect 34388 30232 34390 30252
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 35438 30252 35494 30288
rect 35438 30232 35440 30252
rect 35440 30232 35492 30252
rect 35492 30232 35494 30252
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 46294 46960 46350 47016
rect 45558 46280 45614 46336
rect 46754 49000 46810 49056
rect 46846 44940 46902 44976
rect 46846 44920 46848 44940
rect 46848 44920 46900 44940
rect 46900 44920 46902 44940
rect 46846 39500 46902 39536
rect 46846 39480 46848 39500
rect 46848 39480 46900 39500
rect 46900 39480 46902 39500
rect 46478 38120 46534 38176
rect 46846 36080 46902 36136
rect 40590 18692 40646 18728
rect 40590 18672 40592 18692
rect 40592 18672 40644 18692
rect 40644 18672 40646 18692
rect 41878 18692 41934 18728
rect 41878 18672 41880 18692
rect 41880 18672 41932 18692
rect 41932 18672 41934 18692
rect 45558 23840 45614 23896
rect 46846 27920 46902 27976
rect 46846 26560 46902 26616
rect 46754 25880 46810 25936
rect 46846 22480 46902 22536
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 46846 17740 46902 17776
rect 46846 17720 46848 17740
rect 46848 17720 46900 17740
rect 46900 17720 46902 17740
rect 46846 15000 46902 15056
rect 46846 13640 46902 13696
rect 46754 13504 46810 13560
rect 46846 6860 46902 6896
rect 46846 6840 46848 6860
rect 46848 6840 46900 6860
rect 46900 6840 46902 6860
rect 47398 44240 47454 44296
rect 48226 42880 48282 42936
rect 48226 41520 48282 41576
rect 48318 40160 48374 40216
rect 47950 37440 48006 37496
rect 48318 32680 48374 32736
rect 47766 30252 47822 30288
rect 47766 30232 47768 30252
rect 47768 30232 47820 30252
rect 47820 30232 47822 30252
rect 47766 27784 47822 27840
rect 48318 29280 48374 29336
rect 48226 28620 48282 28656
rect 48226 28600 48228 28620
rect 48228 28600 48280 28620
rect 48280 28600 48282 28620
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 46846 5480 46902 5536
rect 48226 24520 48282 24576
rect 48226 21800 48282 21856
rect 48226 20440 48282 20496
rect 48226 19080 48282 19136
rect 48134 17040 48190 17096
rect 48226 12960 48282 13016
rect 47950 12280 48006 12336
rect 48226 8900 48282 8936
rect 48226 8880 48228 8900
rect 48228 8880 48280 8900
rect 48280 8880 48282 8900
rect 48226 8200 48282 8256
rect 48318 3476 48320 3496
rect 48320 3476 48372 3496
rect 48372 3476 48374 3496
rect 48318 3440 48374 3476
rect 46846 2100 46902 2136
rect 46846 2080 46848 2100
rect 46848 2080 46900 2100
rect 46900 2080 46902 2100
rect 46754 1400 46810 1456
rect 48410 40 48466 96
<< metal3 >>
rect 200 49588 800 49828
rect 46749 49058 46815 49061
rect 49200 49058 49800 49148
rect 46749 49056 49800 49058
rect 46749 49000 46754 49056
rect 46810 49000 49800 49056
rect 46749 48998 49800 49000
rect 46749 48995 46815 48998
rect 49200 48908 49800 48998
rect 200 48378 800 48468
rect 2865 48378 2931 48381
rect 200 48376 2931 48378
rect 200 48320 2870 48376
rect 2926 48320 2931 48376
rect 200 48318 2931 48320
rect 200 48228 800 48318
rect 2865 48315 2931 48318
rect 49200 48228 49800 48468
rect 200 47698 800 47788
rect 2773 47698 2839 47701
rect 200 47696 2839 47698
rect 200 47640 2778 47696
rect 2834 47640 2839 47696
rect 200 47638 2839 47640
rect 200 47548 800 47638
rect 2773 47635 2839 47638
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 46289 47018 46355 47021
rect 49200 47018 49800 47108
rect 46289 47016 49800 47018
rect 46289 46960 46294 47016
rect 46350 46960 49800 47016
rect 46289 46958 49800 46960
rect 46289 46955 46355 46958
rect 49200 46868 49800 46958
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 200 46338 800 46428
rect 4061 46338 4127 46341
rect 200 46336 4127 46338
rect 200 46280 4066 46336
rect 4122 46280 4127 46336
rect 200 46278 4127 46280
rect 200 46188 800 46278
rect 4061 46275 4127 46278
rect 45553 46338 45619 46341
rect 49200 46338 49800 46428
rect 45553 46336 49800 46338
rect 45553 46280 45558 46336
rect 45614 46280 49800 46336
rect 45553 46278 49800 46280
rect 45553 46275 45619 46278
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 49200 46188 49800 46278
rect 200 45658 800 45748
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 3141 45658 3207 45661
rect 200 45656 3207 45658
rect 200 45600 3146 45656
rect 3202 45600 3207 45656
rect 200 45598 3207 45600
rect 200 45508 800 45598
rect 3141 45595 3207 45598
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 46841 44978 46907 44981
rect 49200 44978 49800 45068
rect 46841 44976 49800 44978
rect 46841 44920 46846 44976
rect 46902 44920 49800 44976
rect 46841 44918 49800 44920
rect 46841 44915 46907 44918
rect 49200 44828 49800 44918
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 200 44148 800 44388
rect 47393 44298 47459 44301
rect 47894 44298 47900 44300
rect 47393 44296 47900 44298
rect 47393 44240 47398 44296
rect 47454 44240 47900 44296
rect 47393 44238 47900 44240
rect 47393 44235 47459 44238
rect 47894 44236 47900 44238
rect 47964 44236 47970 44300
rect 49200 44148 49800 44388
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 200 43618 800 43708
rect 2773 43618 2839 43621
rect 200 43616 2839 43618
rect 200 43560 2778 43616
rect 2834 43560 2839 43616
rect 200 43558 2839 43560
rect 200 43468 800 43558
rect 2773 43555 2839 43558
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 200 42788 800 43028
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 48221 42938 48287 42941
rect 49200 42938 49800 43028
rect 48221 42936 49800 42938
rect 48221 42880 48226 42936
rect 48282 42880 49800 42936
rect 48221 42878 49800 42880
rect 48221 42875 48287 42878
rect 49200 42788 49800 42878
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 49200 42108 49800 42348
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 200 41578 800 41668
rect 3049 41578 3115 41581
rect 200 41576 3115 41578
rect 200 41520 3054 41576
rect 3110 41520 3115 41576
rect 200 41518 3115 41520
rect 200 41428 800 41518
rect 3049 41515 3115 41518
rect 48221 41578 48287 41581
rect 49200 41578 49800 41668
rect 48221 41576 49800 41578
rect 48221 41520 48226 41576
rect 48282 41520 49800 41576
rect 48221 41518 49800 41520
rect 48221 41515 48287 41518
rect 49200 41428 49800 41518
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 200 40898 800 40988
rect 3233 40898 3299 40901
rect 200 40896 3299 40898
rect 200 40840 3238 40896
rect 3294 40840 3299 40896
rect 200 40838 3299 40840
rect 200 40748 800 40838
rect 3233 40835 3299 40838
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 48313 40218 48379 40221
rect 49200 40218 49800 40308
rect 48313 40216 49800 40218
rect 48313 40160 48318 40216
rect 48374 40160 49800 40216
rect 48313 40158 49800 40160
rect 48313 40155 48379 40158
rect 49200 40068 49800 40158
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 200 39388 800 39628
rect 46841 39538 46907 39541
rect 49200 39538 49800 39628
rect 46841 39536 49800 39538
rect 46841 39480 46846 39536
rect 46902 39480 49800 39536
rect 46841 39478 49800 39480
rect 46841 39475 46907 39478
rect 49200 39388 49800 39478
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 200 38858 800 38948
rect 1669 38858 1735 38861
rect 200 38856 1735 38858
rect 200 38800 1674 38856
rect 1730 38800 1735 38856
rect 200 38798 1735 38800
rect 200 38708 800 38798
rect 1669 38795 1735 38798
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 46473 38178 46539 38181
rect 49200 38178 49800 38268
rect 46473 38176 49800 38178
rect 46473 38120 46478 38176
rect 46534 38120 49800 38176
rect 46473 38118 49800 38120
rect 46473 38115 46539 38118
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 49200 38028 49800 38118
rect 200 37348 800 37588
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 47945 37498 48011 37501
rect 49200 37498 49800 37588
rect 47945 37496 49800 37498
rect 47945 37440 47950 37496
rect 48006 37440 49800 37496
rect 47945 37438 49800 37440
rect 47945 37435 48011 37438
rect 49200 37348 49800 37438
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 200 36818 800 36908
rect 1669 36818 1735 36821
rect 200 36816 1735 36818
rect 200 36760 1674 36816
rect 1730 36760 1735 36816
rect 200 36758 1735 36760
rect 200 36668 800 36758
rect 1669 36755 1735 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 200 35988 800 36228
rect 46841 36138 46907 36141
rect 49200 36138 49800 36228
rect 46841 36136 49800 36138
rect 46841 36080 46846 36136
rect 46902 36080 49800 36136
rect 46841 36078 49800 36080
rect 46841 36075 46907 36078
rect 49200 35988 49800 36078
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 49200 35308 49800 35548
rect 200 34628 800 34868
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 49200 34628 49800 34868
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 200 34098 800 34188
rect 1577 34098 1643 34101
rect 200 34096 1643 34098
rect 200 34040 1582 34096
rect 1638 34040 1643 34096
rect 200 34038 1643 34040
rect 200 33948 800 34038
rect 1577 34035 1643 34038
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 49200 33268 49800 33508
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 200 32738 800 32828
rect 4061 32738 4127 32741
rect 200 32736 4127 32738
rect 200 32680 4066 32736
rect 4122 32680 4127 32736
rect 200 32678 4127 32680
rect 200 32588 800 32678
rect 4061 32675 4127 32678
rect 48313 32738 48379 32741
rect 49200 32738 49800 32828
rect 48313 32736 49800 32738
rect 48313 32680 48318 32736
rect 48374 32680 49800 32736
rect 48313 32678 49800 32680
rect 48313 32675 48379 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 49200 32588 49800 32678
rect 200 32058 800 32148
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 1577 32058 1643 32061
rect 200 32056 1643 32058
rect 200 32000 1582 32056
rect 1638 32000 1643 32056
rect 200 31998 1643 32000
rect 200 31908 800 31998
rect 1577 31995 1643 31998
rect 25814 31588 25820 31652
rect 25884 31650 25890 31652
rect 25957 31650 26023 31653
rect 25884 31648 26023 31650
rect 25884 31592 25962 31648
rect 26018 31592 26023 31648
rect 25884 31590 26023 31592
rect 25884 31588 25890 31590
rect 25957 31587 26023 31590
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 49200 31228 49800 31468
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 200 30548 800 30788
rect 49200 30548 49800 30788
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 34329 30290 34395 30293
rect 35433 30290 35499 30293
rect 34329 30288 35499 30290
rect 34329 30232 34334 30288
rect 34390 30232 35438 30288
rect 35494 30232 35499 30288
rect 34329 30230 35499 30232
rect 34329 30227 34395 30230
rect 35433 30227 35499 30230
rect 47761 30290 47827 30293
rect 47894 30290 47900 30292
rect 47761 30288 47900 30290
rect 47761 30232 47766 30288
rect 47822 30232 47900 30288
rect 47761 30230 47900 30232
rect 47761 30227 47827 30230
rect 47894 30228 47900 30230
rect 47964 30228 47970 30292
rect 200 29868 800 30108
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 200 29188 800 29428
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 48313 29338 48379 29341
rect 49200 29338 49800 29428
rect 48313 29336 49800 29338
rect 48313 29280 48318 29336
rect 48374 29280 49800 29336
rect 48313 29278 49800 29280
rect 48313 29275 48379 29278
rect 49200 29188 49800 29278
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 48221 28658 48287 28661
rect 49200 28658 49800 28748
rect 48221 28656 49800 28658
rect 48221 28600 48226 28656
rect 48282 28600 49800 28656
rect 48221 28598 49800 28600
rect 48221 28595 48287 28598
rect 49200 28508 49800 28598
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 200 27828 800 28068
rect 46841 27978 46907 27981
rect 49200 27978 49800 28068
rect 46841 27976 49800 27978
rect 46841 27920 46846 27976
rect 46902 27920 49800 27976
rect 46841 27918 49800 27920
rect 46841 27915 46907 27918
rect 47761 27842 47827 27845
rect 47894 27842 47900 27844
rect 47761 27840 47900 27842
rect 47761 27784 47766 27840
rect 47822 27784 47900 27840
rect 47761 27782 47900 27784
rect 47761 27779 47827 27782
rect 47894 27780 47900 27782
rect 47964 27780 47970 27844
rect 49200 27828 49800 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 200 27148 800 27388
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 46841 26618 46907 26621
rect 49200 26618 49800 26708
rect 46841 26616 49800 26618
rect 46841 26560 46846 26616
rect 46902 26560 49800 26616
rect 46841 26558 49800 26560
rect 46841 26555 46907 26558
rect 49200 26468 49800 26558
rect 25589 26210 25655 26213
rect 25814 26210 25820 26212
rect 25589 26208 25820 26210
rect 25589 26152 25594 26208
rect 25650 26152 25820 26208
rect 25589 26150 25820 26152
rect 25589 26147 25655 26150
rect 25814 26148 25820 26150
rect 25884 26148 25890 26212
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 200 25788 800 26028
rect 46749 25938 46815 25941
rect 49200 25938 49800 26028
rect 46749 25936 49800 25938
rect 46749 25880 46754 25936
rect 46810 25880 49800 25936
rect 46749 25878 49800 25880
rect 46749 25875 46815 25878
rect 49200 25788 49800 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 200 25258 800 25348
rect 1577 25258 1643 25261
rect 200 25256 1643 25258
rect 200 25200 1582 25256
rect 1638 25200 1643 25256
rect 200 25198 1643 25200
rect 200 25108 800 25198
rect 1577 25195 1643 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 48221 24578 48287 24581
rect 49200 24578 49800 24668
rect 48221 24576 49800 24578
rect 48221 24520 48226 24576
rect 48282 24520 49800 24576
rect 48221 24518 49800 24520
rect 48221 24515 48287 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 49200 24428 49800 24518
rect 200 23898 800 23988
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 3325 23898 3391 23901
rect 200 23896 3391 23898
rect 200 23840 3330 23896
rect 3386 23840 3391 23896
rect 200 23838 3391 23840
rect 200 23748 800 23838
rect 3325 23835 3391 23838
rect 45553 23898 45619 23901
rect 49200 23898 49800 23988
rect 45553 23896 49800 23898
rect 45553 23840 45558 23896
rect 45614 23840 49800 23896
rect 45553 23838 49800 23840
rect 45553 23835 45619 23838
rect 49200 23748 49800 23838
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 200 23068 800 23308
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 46841 22538 46907 22541
rect 49200 22538 49800 22628
rect 46841 22536 49800 22538
rect 46841 22480 46846 22536
rect 46902 22480 49800 22536
rect 46841 22478 49800 22480
rect 46841 22475 46907 22478
rect 49200 22388 49800 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 27153 22130 27219 22133
rect 27429 22130 27495 22133
rect 27153 22128 27495 22130
rect 27153 22072 27158 22128
rect 27214 22072 27434 22128
rect 27490 22072 27495 22128
rect 27153 22070 27495 22072
rect 27153 22067 27219 22070
rect 27429 22067 27495 22070
rect 200 21858 800 21948
rect 1577 21858 1643 21861
rect 200 21856 1643 21858
rect 200 21800 1582 21856
rect 1638 21800 1643 21856
rect 200 21798 1643 21800
rect 200 21708 800 21798
rect 1577 21795 1643 21798
rect 48221 21858 48287 21861
rect 49200 21858 49800 21948
rect 48221 21856 49800 21858
rect 48221 21800 48226 21856
rect 48282 21800 49800 21856
rect 48221 21798 49800 21800
rect 48221 21795 48287 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 49200 21708 49800 21798
rect 200 21028 800 21268
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 200 20498 800 20588
rect 2773 20498 2839 20501
rect 200 20496 2839 20498
rect 200 20440 2778 20496
rect 2834 20440 2839 20496
rect 200 20438 2839 20440
rect 200 20348 800 20438
rect 2773 20435 2839 20438
rect 17033 20498 17099 20501
rect 18137 20498 18203 20501
rect 17033 20496 18203 20498
rect 17033 20440 17038 20496
rect 17094 20440 18142 20496
rect 18198 20440 18203 20496
rect 17033 20438 18203 20440
rect 17033 20435 17099 20438
rect 18137 20435 18203 20438
rect 48221 20498 48287 20501
rect 49200 20498 49800 20588
rect 48221 20496 49800 20498
rect 48221 20440 48226 20496
rect 48282 20440 49800 20496
rect 48221 20438 49800 20440
rect 48221 20435 48287 20438
rect 16665 20362 16731 20365
rect 17953 20362 18019 20365
rect 16665 20360 18019 20362
rect 16665 20304 16670 20360
rect 16726 20304 17958 20360
rect 18014 20304 18019 20360
rect 49200 20348 49800 20438
rect 16665 20302 18019 20304
rect 16665 20299 16731 20302
rect 17953 20299 18019 20302
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 49200 19668 49800 19908
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 22093 19274 22159 19277
rect 27705 19274 27771 19277
rect 22093 19272 27771 19274
rect 200 18988 800 19228
rect 22093 19216 22098 19272
rect 22154 19216 27710 19272
rect 27766 19216 27771 19272
rect 22093 19214 27771 19216
rect 22093 19211 22159 19214
rect 27705 19211 27771 19214
rect 48221 19138 48287 19141
rect 49200 19138 49800 19228
rect 48221 19136 49800 19138
rect 48221 19080 48226 19136
rect 48282 19080 49800 19136
rect 48221 19078 49800 19080
rect 48221 19075 48287 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 49200 18988 49800 19078
rect 40585 18730 40651 18733
rect 41873 18730 41939 18733
rect 40585 18728 41939 18730
rect 40585 18672 40590 18728
rect 40646 18672 41878 18728
rect 41934 18672 41939 18728
rect 40585 18670 41939 18672
rect 40585 18667 40651 18670
rect 41873 18667 41939 18670
rect 200 18458 800 18548
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 2773 18458 2839 18461
rect 200 18456 2839 18458
rect 200 18400 2778 18456
rect 2834 18400 2839 18456
rect 200 18398 2839 18400
rect 200 18308 800 18398
rect 2773 18395 2839 18398
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 46841 17778 46907 17781
rect 49200 17778 49800 17868
rect 46841 17776 49800 17778
rect 46841 17720 46846 17776
rect 46902 17720 49800 17776
rect 46841 17718 49800 17720
rect 46841 17715 46907 17718
rect 49200 17628 49800 17718
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 200 17098 800 17188
rect 2865 17098 2931 17101
rect 200 17096 2931 17098
rect 200 17040 2870 17096
rect 2926 17040 2931 17096
rect 200 17038 2931 17040
rect 200 16948 800 17038
rect 2865 17035 2931 17038
rect 48129 17098 48195 17101
rect 49200 17098 49800 17188
rect 48129 17096 49800 17098
rect 48129 17040 48134 17096
rect 48190 17040 49800 17096
rect 48129 17038 49800 17040
rect 48129 17035 48195 17038
rect 49200 16948 49800 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 200 16268 800 16508
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 49200 15588 49800 15828
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 200 15058 800 15148
rect 3417 15058 3483 15061
rect 200 15056 3483 15058
rect 200 15000 3422 15056
rect 3478 15000 3483 15056
rect 200 14998 3483 15000
rect 200 14908 800 14998
rect 3417 14995 3483 14998
rect 46841 15058 46907 15061
rect 49200 15058 49800 15148
rect 46841 15056 49800 15058
rect 46841 15000 46846 15056
rect 46902 15000 49800 15056
rect 46841 14998 49800 15000
rect 46841 14995 46907 14998
rect 49200 14908 49800 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 200 14378 800 14468
rect 1577 14378 1643 14381
rect 200 14376 1643 14378
rect 200 14320 1582 14376
rect 1638 14320 1643 14376
rect 200 14318 1643 14320
rect 200 14228 800 14318
rect 1577 14315 1643 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 200 13548 800 13788
rect 46841 13698 46907 13701
rect 49200 13698 49800 13788
rect 46841 13696 49800 13698
rect 46841 13640 46846 13696
rect 46902 13640 49800 13696
rect 46841 13638 49800 13640
rect 46841 13635 46907 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 46749 13562 46815 13565
rect 47894 13562 47900 13564
rect 46749 13560 47900 13562
rect 46749 13504 46754 13560
rect 46810 13504 47900 13560
rect 46749 13502 47900 13504
rect 46749 13499 46815 13502
rect 47894 13500 47900 13502
rect 47964 13500 47970 13564
rect 49200 13548 49800 13638
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 48221 13018 48287 13021
rect 49200 13018 49800 13108
rect 48221 13016 49800 13018
rect 48221 12960 48226 13016
rect 48282 12960 49800 13016
rect 48221 12958 49800 12960
rect 48221 12955 48287 12958
rect 49200 12868 49800 12958
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 200 12188 800 12428
rect 47945 12338 48011 12341
rect 49200 12338 49800 12428
rect 47945 12336 49800 12338
rect 47945 12280 47950 12336
rect 48006 12280 49800 12336
rect 47945 12278 49800 12280
rect 47945 12275 48011 12278
rect 49200 12188 49800 12278
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 200 11658 800 11748
rect 2773 11658 2839 11661
rect 200 11656 2839 11658
rect 200 11600 2778 11656
rect 2834 11600 2839 11656
rect 200 11598 2839 11600
rect 200 11508 800 11598
rect 2773 11595 2839 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 49200 10828 49800 11068
rect 200 10298 800 10388
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 1577 10298 1643 10301
rect 200 10296 1643 10298
rect 200 10240 1582 10296
rect 1638 10240 1643 10296
rect 200 10238 1643 10240
rect 200 10148 800 10238
rect 1577 10235 1643 10238
rect 49200 10148 49800 10388
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 200 9618 800 9708
rect 2957 9618 3023 9621
rect 200 9616 3023 9618
rect 200 9560 2962 9616
rect 3018 9560 3023 9616
rect 200 9558 3023 9560
rect 200 9468 800 9558
rect 2957 9555 3023 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 48221 8938 48287 8941
rect 49200 8938 49800 9028
rect 48221 8936 49800 8938
rect 48221 8880 48226 8936
rect 48282 8880 49800 8936
rect 48221 8878 49800 8880
rect 48221 8875 48287 8878
rect 49200 8788 49800 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 200 8108 800 8348
rect 48221 8258 48287 8261
rect 49200 8258 49800 8348
rect 48221 8256 49800 8258
rect 48221 8200 48226 8256
rect 48282 8200 49800 8256
rect 48221 8198 49800 8200
rect 48221 8195 48287 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 49200 8108 49800 8198
rect 200 7578 800 7668
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 1577 7578 1643 7581
rect 200 7576 1643 7578
rect 200 7520 1582 7576
rect 1638 7520 1643 7576
rect 200 7518 1643 7520
rect 200 7428 800 7518
rect 1577 7515 1643 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 200 6898 800 6988
rect 1577 6898 1643 6901
rect 200 6896 1643 6898
rect 200 6840 1582 6896
rect 1638 6840 1643 6896
rect 200 6838 1643 6840
rect 200 6748 800 6838
rect 1577 6835 1643 6838
rect 46841 6898 46907 6901
rect 49200 6898 49800 6988
rect 46841 6896 49800 6898
rect 46841 6840 46846 6896
rect 46902 6840 49800 6896
rect 46841 6838 49800 6840
rect 46841 6835 46907 6838
rect 49200 6748 49800 6838
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 49200 6068 49800 6308
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 200 5538 800 5628
rect 1577 5538 1643 5541
rect 200 5536 1643 5538
rect 200 5480 1582 5536
rect 1638 5480 1643 5536
rect 200 5478 1643 5480
rect 200 5388 800 5478
rect 1577 5475 1643 5478
rect 46841 5538 46907 5541
rect 49200 5538 49800 5628
rect 46841 5536 49800 5538
rect 46841 5480 46846 5536
rect 46902 5480 49800 5536
rect 46841 5478 49800 5480
rect 46841 5475 46907 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 49200 5388 49800 5478
rect 200 4858 800 4948
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 2773 4858 2839 4861
rect 200 4856 2839 4858
rect 200 4800 2778 4856
rect 2834 4800 2839 4856
rect 200 4798 2839 4800
rect 200 4708 800 4798
rect 2773 4795 2839 4798
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 49200 4028 49800 4268
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 200 3498 800 3588
rect 1577 3498 1643 3501
rect 200 3496 1643 3498
rect 200 3440 1582 3496
rect 1638 3440 1643 3496
rect 200 3438 1643 3440
rect 200 3348 800 3438
rect 1577 3435 1643 3438
rect 48313 3498 48379 3501
rect 49200 3498 49800 3588
rect 48313 3496 49800 3498
rect 48313 3440 48318 3496
rect 48374 3440 49800 3496
rect 48313 3438 49800 3440
rect 48313 3435 48379 3438
rect 49200 3348 49800 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 200 2818 800 2908
rect 1577 2818 1643 2821
rect 200 2816 1643 2818
rect 200 2760 1582 2816
rect 1638 2760 1643 2816
rect 200 2758 1643 2760
rect 200 2668 800 2758
rect 1577 2755 1643 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 46841 2138 46907 2141
rect 49200 2138 49800 2228
rect 46841 2136 49800 2138
rect 46841 2080 46846 2136
rect 46902 2080 49800 2136
rect 46841 2078 49800 2080
rect 46841 2075 46907 2078
rect 49200 1988 49800 2078
rect 200 1458 800 1548
rect 2865 1458 2931 1461
rect 200 1456 2931 1458
rect 200 1400 2870 1456
rect 2926 1400 2931 1456
rect 200 1398 2931 1400
rect 200 1308 800 1398
rect 2865 1395 2931 1398
rect 46749 1458 46815 1461
rect 49200 1458 49800 1548
rect 46749 1456 49800 1458
rect 46749 1400 46754 1456
rect 46810 1400 49800 1456
rect 46749 1398 49800 1400
rect 46749 1395 46815 1398
rect 49200 1308 49800 1398
rect 200 778 800 868
rect 2773 778 2839 781
rect 200 776 2839 778
rect 200 720 2778 776
rect 2834 720 2839 776
rect 200 718 2839 720
rect 200 628 800 718
rect 2773 715 2839 718
rect 48405 98 48471 101
rect 49200 98 49800 188
rect 48405 96 49800 98
rect 48405 40 48410 96
rect 48466 40 49800 96
rect 48405 38 49800 40
rect 48405 35 48471 38
rect 49200 -52 49800 38
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 47900 44236 47964 44300
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 25820 31588 25884 31652
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 47900 30228 47964 30292
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 47900 27780 47964 27844
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 25820 26148 25884 26212
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 47900 13500 47964 13564
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 46816 19888 47376
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 47899 44300 47965 44301
rect 47899 44236 47900 44300
rect 47964 44236 47965 44300
rect 47899 44235 47965 44236
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 25819 31652 25885 31653
rect 25819 31588 25820 31652
rect 25884 31588 25885 31652
rect 25819 31587 25885 31588
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 25822 26213 25882 31587
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 47902 30293 47962 44235
rect 47899 30292 47965 30293
rect 47899 30228 47900 30292
rect 47964 30228 47965 30292
rect 47899 30227 47965 30228
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 47899 27844 47965 27845
rect 47899 27780 47900 27844
rect 47964 27780 47965 27844
rect 47899 27779 47965 27780
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 25819 26212 25885 26213
rect 25819 26148 25820 26212
rect 25884 26148 25885 26212
rect 25819 26147 25885 26148
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 47902 13565 47962 27779
rect 47899 13564 47965 13565
rect 47899 13500 47900 13564
rect 47964 13500 47965 13564
rect 47899 13499 47965 13500
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1667941163
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1667941163
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1667941163
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1667941163
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1667941163
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1667941163
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147
timestamp 1667941163
transform 1 0 14628 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_159 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 15732 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1667941163
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1667941163
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1667941163
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1667941163
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1667941163
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_261
timestamp 1667941163
transform 1 0 25116 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_266
timestamp 1667941163
transform 1 0 25576 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1667941163
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1667941163
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1667941163
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_315
timestamp 1667941163
transform 1 0 30084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_327
timestamp 1667941163
transform 1 0 31188 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1667941163
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1667941163
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1667941163
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1667941163
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1667941163
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_405
timestamp 1667941163
transform 1 0 38364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_413 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 39100 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1667941163
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1667941163
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1667941163
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1667941163
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_449
timestamp 1667941163
transform 1 0 42412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_474
timestamp 1667941163
transform 1 0 44712 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_477
timestamp 1667941163
transform 1 0 44988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_502
timestamp 1667941163
transform 1 0 47288 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_505
timestamp 1667941163
transform 1 0 47564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_510
timestamp 1667941163
transform 1 0 48024 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7
timestamp 1667941163
transform 1 0 1748 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_29
timestamp 1667941163
transform 1 0 3772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1667941163
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_63
timestamp 1667941163
transform 1 0 6900 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_90
timestamp 1667941163
transform 1 0 9384 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1667941163
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1667941163
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_119
timestamp 1667941163
transform 1 0 12052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_126
timestamp 1667941163
transform 1 0 12696 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_130
timestamp 1667941163
transform 1 0 13064 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_152
timestamp 1667941163
transform 1 0 15088 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1667941163
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_192
timestamp 1667941163
transform 1 0 18768 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_200
timestamp 1667941163
transform 1 0 19504 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1667941163
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1667941163
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_249
timestamp 1667941163
transform 1 0 24012 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1667941163
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_304
timestamp 1667941163
transform 1 0 29072 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_316
timestamp 1667941163
transform 1 0 30176 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_328
timestamp 1667941163
transform 1 0 31280 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1667941163
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1667941163
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1667941163
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1667941163
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1667941163
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_430
timestamp 1667941163
transform 1 0 40664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_437
timestamp 1667941163
transform 1 0 41308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_444
timestamp 1667941163
transform 1 0 41952 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_449
timestamp 1667941163
transform 1 0 42412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_472
timestamp 1667941163
transform 1 0 44528 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1667941163
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1667941163
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_505
timestamp 1667941163
transform 1 0 47564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_510
timestamp 1667941163
transform 1 0 48024 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1667941163
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_34
timestamp 1667941163
transform 1 0 4232 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_41
timestamp 1667941163
transform 1 0 4876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_48
timestamp 1667941163
transform 1 0 5520 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_73
timestamp 1667941163
transform 1 0 7820 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1667941163
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_101
timestamp 1667941163
transform 1 0 10396 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_123
timestamp 1667941163
transform 1 0 12420 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_134
timestamp 1667941163
transform 1 0 13432 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1667941163
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_165
timestamp 1667941163
transform 1 0 16284 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_169
timestamp 1667941163
transform 1 0 16652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_173
timestamp 1667941163
transform 1 0 17020 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_180
timestamp 1667941163
transform 1 0 17664 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_188
timestamp 1667941163
transform 1 0 18400 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1667941163
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_202
timestamp 1667941163
transform 1 0 19688 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_212
timestamp 1667941163
transform 1 0 20608 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_224
timestamp 1667941163
transform 1 0 21712 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_236
timestamp 1667941163
transform 1 0 22816 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1667941163
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_264
timestamp 1667941163
transform 1 0 25392 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_289
timestamp 1667941163
transform 1 0 27692 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_296
timestamp 1667941163
transform 1 0 28336 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1667941163
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1667941163
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1667941163
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1667941163
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1667941163
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1667941163
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_401
timestamp 1667941163
transform 1 0 37996 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_405
timestamp 1667941163
transform 1 0 38364 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_412
timestamp 1667941163
transform 1 0 39008 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_421
timestamp 1667941163
transform 1 0 39836 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_450
timestamp 1667941163
transform 1 0 42504 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_457
timestamp 1667941163
transform 1 0 43148 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_471
timestamp 1667941163
transform 1 0 44436 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1667941163
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_477
timestamp 1667941163
transform 1 0 44988 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_500
timestamp 1667941163
transform 1 0 47104 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_508
timestamp 1667941163
transform 1 0 47840 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_514
timestamp 1667941163
transform 1 0 48392 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_11
timestamp 1667941163
transform 1 0 2116 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_22
timestamp 1667941163
transform 1 0 3128 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_30
timestamp 1667941163
transform 1 0 3864 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_35
timestamp 1667941163
transform 1 0 4324 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_41
timestamp 1667941163
transform 1 0 4876 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_45
timestamp 1667941163
transform 1 0 5244 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1667941163
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_63
timestamp 1667941163
transform 1 0 6900 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_69
timestamp 1667941163
transform 1 0 7452 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_73
timestamp 1667941163
transform 1 0 7820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_85
timestamp 1667941163
transform 1 0 8924 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_97
timestamp 1667941163
transform 1 0 10028 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_101
timestamp 1667941163
transform 1 0 10396 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1667941163
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1667941163
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_121
timestamp 1667941163
transform 1 0 12236 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_125
timestamp 1667941163
transform 1 0 12604 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_134
timestamp 1667941163
transform 1 0 13432 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_146
timestamp 1667941163
transform 1 0 14536 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_158
timestamp 1667941163
transform 1 0 15640 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1667941163
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_181
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_189
timestamp 1667941163
transform 1 0 18492 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1667941163
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_205
timestamp 1667941163
transform 1 0 19964 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_209
timestamp 1667941163
transform 1 0 20332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_221
timestamp 1667941163
transform 1 0 21436 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1667941163
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1667941163
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_261
timestamp 1667941163
transform 1 0 25116 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_266
timestamp 1667941163
transform 1 0 25576 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1667941163
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1667941163
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_286
timestamp 1667941163
transform 1 0 27416 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_298
timestamp 1667941163
transform 1 0 28520 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_310
timestamp 1667941163
transform 1 0 29624 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_322
timestamp 1667941163
transform 1 0 30728 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp 1667941163
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1667941163
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1667941163
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1667941163
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_408
timestamp 1667941163
transform 1 0 38640 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_433
timestamp 1667941163
transform 1 0 40940 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_440
timestamp 1667941163
transform 1 0 41584 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_449
timestamp 1667941163
transform 1 0 42412 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_472
timestamp 1667941163
transform 1 0 44528 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1667941163
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1667941163
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_505
timestamp 1667941163
transform 1 0 47564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_510
timestamp 1667941163
transform 1 0 48024 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_9
timestamp 1667941163
transform 1 0 1932 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_16
timestamp 1667941163
transform 1 0 2576 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_23
timestamp 1667941163
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1667941163
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_34
timestamp 1667941163
transform 1 0 4232 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_41
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_48
timestamp 1667941163
transform 1 0 5520 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_60
timestamp 1667941163
transform 1 0 6624 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_72
timestamp 1667941163
transform 1 0 7728 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1667941163
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1667941163
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1667941163
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1667941163
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1667941163
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1667941163
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1667941163
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1667941163
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1667941163
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1667941163
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1667941163
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1667941163
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1667941163
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1667941163
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1667941163
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1667941163
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1667941163
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1667941163
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1667941163
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1667941163
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1667941163
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1667941163
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1667941163
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1667941163
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1667941163
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_401
timestamp 1667941163
transform 1 0 37996 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_409
timestamp 1667941163
transform 1 0 38732 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_415
timestamp 1667941163
transform 1 0 39284 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1667941163
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1667941163
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1667941163
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_445
timestamp 1667941163
transform 1 0 42044 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_453
timestamp 1667941163
transform 1 0 42780 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_459
timestamp 1667941163
transform 1 0 43332 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_466
timestamp 1667941163
transform 1 0 43976 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_473
timestamp 1667941163
transform 1 0 44620 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_477
timestamp 1667941163
transform 1 0 44988 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_482
timestamp 1667941163
transform 1 0 45448 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_489
timestamp 1667941163
transform 1 0 46092 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_514
timestamp 1667941163
transform 1 0 48392 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_32
timestamp 1667941163
transform 1 0 4048 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1667941163
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1667941163
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1667941163
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1667941163
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1667941163
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1667941163
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1667941163
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1667941163
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1667941163
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1667941163
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1667941163
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1667941163
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1667941163
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1667941163
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1667941163
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1667941163
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1667941163
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1667941163
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1667941163
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1667941163
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1667941163
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1667941163
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1667941163
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1667941163
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1667941163
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1667941163
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1667941163
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1667941163
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1667941163
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1667941163
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1667941163
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1667941163
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1667941163
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1667941163
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1667941163
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_473
timestamp 1667941163
transform 1 0 44620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_477
timestamp 1667941163
transform 1 0 44988 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_502
timestamp 1667941163
transform 1 0 47288 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_505
timestamp 1667941163
transform 1 0 47564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_510
timestamp 1667941163
transform 1 0 48024 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1667941163
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_34
timestamp 1667941163
transform 1 0 4232 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_46
timestamp 1667941163
transform 1 0 5336 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_58
timestamp 1667941163
transform 1 0 6440 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_70
timestamp 1667941163
transform 1 0 7544 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1667941163
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1667941163
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1667941163
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1667941163
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1667941163
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1667941163
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1667941163
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1667941163
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1667941163
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1667941163
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1667941163
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1667941163
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1667941163
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1667941163
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1667941163
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1667941163
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1667941163
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1667941163
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1667941163
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1667941163
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1667941163
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1667941163
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1667941163
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1667941163
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1667941163
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1667941163
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1667941163
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1667941163
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1667941163
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1667941163
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1667941163
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1667941163
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1667941163
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1667941163
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_477
timestamp 1667941163
transform 1 0 44988 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_481
timestamp 1667941163
transform 1 0 45356 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_485
timestamp 1667941163
transform 1 0 45724 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_510
timestamp 1667941163
transform 1 0 48024 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_9
timestamp 1667941163
transform 1 0 1932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_16
timestamp 1667941163
transform 1 0 2576 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_23
timestamp 1667941163
transform 1 0 3220 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_35
timestamp 1667941163
transform 1 0 4324 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_47
timestamp 1667941163
transform 1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1667941163
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1667941163
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1667941163
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1667941163
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1667941163
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1667941163
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1667941163
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1667941163
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1667941163
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1667941163
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1667941163
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1667941163
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1667941163
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1667941163
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1667941163
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1667941163
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1667941163
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1667941163
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1667941163
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1667941163
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1667941163
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1667941163
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1667941163
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1667941163
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1667941163
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_342
timestamp 1667941163
transform 1 0 32568 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_354
timestamp 1667941163
transform 1 0 33672 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_366
timestamp 1667941163
transform 1 0 34776 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_378
timestamp 1667941163
transform 1 0 35880 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_390
timestamp 1667941163
transform 1 0 36984 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1667941163
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1667941163
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1667941163
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1667941163
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_449
timestamp 1667941163
transform 1 0 42412 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_458
timestamp 1667941163
transform 1 0 43240 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_470
timestamp 1667941163
transform 1 0 44344 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_482
timestamp 1667941163
transform 1 0 45448 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_490
timestamp 1667941163
transform 1 0 46184 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_495
timestamp 1667941163
transform 1 0 46644 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_502
timestamp 1667941163
transform 1 0 47288 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_505
timestamp 1667941163
transform 1 0 47564 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_510
timestamp 1667941163
transform 1 0 48024 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1667941163
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1667941163
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1667941163
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1667941163
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1667941163
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1667941163
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1667941163
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1667941163
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1667941163
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1667941163
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1667941163
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1667941163
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1667941163
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1667941163
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1667941163
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1667941163
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1667941163
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1667941163
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1667941163
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1667941163
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1667941163
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1667941163
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1667941163
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1667941163
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1667941163
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_330
timestamp 1667941163
transform 1 0 31464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_355
timestamp 1667941163
transform 1 0 33764 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1667941163
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1667941163
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1667941163
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1667941163
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1667941163
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1667941163
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_445
timestamp 1667941163
transform 1 0 42044 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_474
timestamp 1667941163
transform 1 0 44712 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1667941163
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_489
timestamp 1667941163
transform 1 0 46092 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_493
timestamp 1667941163
transform 1 0 46460 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_500
timestamp 1667941163
transform 1 0 47104 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_507
timestamp 1667941163
transform 1 0 47748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_514
timestamp 1667941163
transform 1 0 48392 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_14
timestamp 1667941163
transform 1 0 2392 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_21
timestamp 1667941163
transform 1 0 3036 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_28
timestamp 1667941163
transform 1 0 3680 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_40
timestamp 1667941163
transform 1 0 4784 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1667941163
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1667941163
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1667941163
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1667941163
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1667941163
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1667941163
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1667941163
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1667941163
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1667941163
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1667941163
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1667941163
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1667941163
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1667941163
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1667941163
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1667941163
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1667941163
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1667941163
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1667941163
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1667941163
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1667941163
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1667941163
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1667941163
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1667941163
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1667941163
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1667941163
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1667941163
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1667941163
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1667941163
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1667941163
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1667941163
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1667941163
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1667941163
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_449
timestamp 1667941163
transform 1 0 42412 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_457
timestamp 1667941163
transform 1 0 43148 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1667941163
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1667941163
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1667941163
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1667941163
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1667941163
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_505
timestamp 1667941163
transform 1 0 47564 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_513
timestamp 1667941163
transform 1 0 48300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1667941163
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1667941163
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1667941163
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1667941163
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1667941163
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1667941163
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1667941163
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1667941163
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1667941163
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1667941163
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1667941163
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1667941163
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1667941163
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1667941163
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1667941163
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1667941163
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1667941163
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1667941163
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1667941163
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1667941163
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1667941163
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1667941163
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1667941163
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1667941163
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1667941163
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1667941163
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1667941163
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1667941163
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1667941163
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1667941163
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1667941163
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1667941163
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1667941163
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1667941163
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1667941163
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1667941163
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1667941163
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1667941163
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1667941163
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1667941163
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1667941163
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1667941163
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_513
timestamp 1667941163
transform 1 0 48300 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1667941163
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1667941163
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1667941163
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1667941163
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1667941163
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1667941163
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1667941163
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1667941163
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1667941163
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1667941163
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1667941163
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1667941163
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1667941163
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1667941163
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1667941163
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1667941163
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1667941163
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1667941163
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1667941163
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1667941163
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1667941163
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1667941163
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1667941163
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1667941163
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1667941163
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1667941163
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1667941163
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1667941163
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1667941163
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1667941163
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1667941163
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1667941163
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1667941163
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1667941163
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1667941163
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1667941163
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1667941163
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1667941163
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1667941163
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1667941163
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_505
timestamp 1667941163
transform 1 0 47564 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_514
timestamp 1667941163
transform 1 0 48392 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_14
timestamp 1667941163
transform 1 0 2392 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_21
timestamp 1667941163
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1667941163
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1667941163
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1667941163
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1667941163
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1667941163
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1667941163
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1667941163
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1667941163
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1667941163
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1667941163
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1667941163
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1667941163
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1667941163
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1667941163
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1667941163
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1667941163
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1667941163
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1667941163
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1667941163
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1667941163
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1667941163
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1667941163
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1667941163
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1667941163
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1667941163
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1667941163
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1667941163
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1667941163
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1667941163
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1667941163
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1667941163
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1667941163
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1667941163
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1667941163
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1667941163
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1667941163
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1667941163
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1667941163
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1667941163
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1667941163
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1667941163
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1667941163
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_501
timestamp 1667941163
transform 1 0 47196 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_507
timestamp 1667941163
transform 1 0 47748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_514
timestamp 1667941163
transform 1 0 48392 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_9
timestamp 1667941163
transform 1 0 1932 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_31
timestamp 1667941163
transform 1 0 3956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_43
timestamp 1667941163
transform 1 0 5060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1667941163
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1667941163
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1667941163
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1667941163
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1667941163
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1667941163
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1667941163
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1667941163
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1667941163
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1667941163
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1667941163
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1667941163
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1667941163
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1667941163
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1667941163
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_230
timestamp 1667941163
transform 1 0 22264 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_241
timestamp 1667941163
transform 1 0 23276 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_248
timestamp 1667941163
transform 1 0 23920 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_260
timestamp 1667941163
transform 1 0 25024 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_272
timestamp 1667941163
transform 1 0 26128 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1667941163
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1667941163
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1667941163
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1667941163
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1667941163
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1667941163
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1667941163
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1667941163
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1667941163
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1667941163
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1667941163
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1667941163
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1667941163
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1667941163
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1667941163
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_505
timestamp 1667941163
transform 1 0 47564 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_513
timestamp 1667941163
transform 1 0 48300 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1667941163
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1667941163
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1667941163
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1667941163
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1667941163
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1667941163
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1667941163
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1667941163
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1667941163
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1667941163
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1667941163
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1667941163
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1667941163
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_177
timestamp 1667941163
transform 1 0 17388 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_185
timestamp 1667941163
transform 1 0 18124 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1667941163
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_203
timestamp 1667941163
transform 1 0 19780 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_213
timestamp 1667941163
transform 1 0 20700 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_226
timestamp 1667941163
transform 1 0 21896 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_237
timestamp 1667941163
transform 1 0 22908 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_248
timestamp 1667941163
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_259
timestamp 1667941163
transform 1 0 24932 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_271
timestamp 1667941163
transform 1 0 26036 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_281
timestamp 1667941163
transform 1 0 26956 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_293
timestamp 1667941163
transform 1 0 28060 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_305
timestamp 1667941163
transform 1 0 29164 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1667941163
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1667941163
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1667941163
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1667941163
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1667941163
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1667941163
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1667941163
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1667941163
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1667941163
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1667941163
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1667941163
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1667941163
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1667941163
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1667941163
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1667941163
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1667941163
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1667941163
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1667941163
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_513
timestamp 1667941163
transform 1 0 48300 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_14
timestamp 1667941163
transform 1 0 2392 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_21
timestamp 1667941163
transform 1 0 3036 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_33
timestamp 1667941163
transform 1 0 4140 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_45
timestamp 1667941163
transform 1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1667941163
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1667941163
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1667941163
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1667941163
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1667941163
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1667941163
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1667941163
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1667941163
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1667941163
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1667941163
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1667941163
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_175
timestamp 1667941163
transform 1 0 17204 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_192
timestamp 1667941163
transform 1 0 18768 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_212
timestamp 1667941163
transform 1 0 20608 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_218
timestamp 1667941163
transform 1 0 21160 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1667941163
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_235
timestamp 1667941163
transform 1 0 22724 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_243
timestamp 1667941163
transform 1 0 23460 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_250
timestamp 1667941163
transform 1 0 24104 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_254
timestamp 1667941163
transform 1 0 24472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_271
timestamp 1667941163
transform 1 0 26036 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1667941163
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_299
timestamp 1667941163
transform 1 0 28612 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_307
timestamp 1667941163
transform 1 0 29348 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_315
timestamp 1667941163
transform 1 0 30084 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_327
timestamp 1667941163
transform 1 0 31188 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1667941163
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_345
timestamp 1667941163
transform 1 0 32844 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_364
timestamp 1667941163
transform 1 0 34592 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_376
timestamp 1667941163
transform 1 0 35696 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_388
timestamp 1667941163
transform 1 0 36800 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1667941163
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1667941163
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1667941163
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1667941163
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1667941163
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1667941163
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1667941163
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1667941163
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1667941163
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1667941163
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_505
timestamp 1667941163
transform 1 0 47564 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_513
timestamp 1667941163
transform 1 0 48300 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_9
timestamp 1667941163
transform 1 0 1932 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_13
timestamp 1667941163
transform 1 0 2300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_25
timestamp 1667941163
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1667941163
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1667941163
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1667941163
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1667941163
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1667941163
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1667941163
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1667941163
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1667941163
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1667941163
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1667941163
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_153
timestamp 1667941163
transform 1 0 15180 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_177
timestamp 1667941163
transform 1 0 17388 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_187
timestamp 1667941163
transform 1 0 18308 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1667941163
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_203
timestamp 1667941163
transform 1 0 19780 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_215
timestamp 1667941163
transform 1 0 20884 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_227
timestamp 1667941163
transform 1 0 21988 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_238
timestamp 1667941163
transform 1 0 23000 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1667941163
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_264
timestamp 1667941163
transform 1 0 25392 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_272
timestamp 1667941163
transform 1 0 26128 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_281
timestamp 1667941163
transform 1 0 26956 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_293
timestamp 1667941163
transform 1 0 28060 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_297
timestamp 1667941163
transform 1 0 28428 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 1667941163
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_327
timestamp 1667941163
transform 1 0 31188 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_331
timestamp 1667941163
transform 1 0 31556 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_348
timestamp 1667941163
transform 1 0 33120 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_360
timestamp 1667941163
transform 1 0 34224 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_370
timestamp 1667941163
transform 1 0 35144 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_386
timestamp 1667941163
transform 1 0 36616 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_393
timestamp 1667941163
transform 1 0 37260 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_405
timestamp 1667941163
transform 1 0 38364 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_417
timestamp 1667941163
transform 1 0 39468 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1667941163
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1667941163
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1667941163
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1667941163
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1667941163
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1667941163
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1667941163
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1667941163
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1667941163
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_513
timestamp 1667941163
transform 1 0 48300 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_9
timestamp 1667941163
transform 1 0 1932 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_31
timestamp 1667941163
transform 1 0 3956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_43
timestamp 1667941163
transform 1 0 5060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1667941163
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1667941163
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1667941163
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1667941163
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1667941163
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1667941163
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1667941163
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1667941163
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1667941163
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1667941163
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1667941163
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_174
timestamp 1667941163
transform 1 0 17112 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_186
timestamp 1667941163
transform 1 0 18216 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_200
timestamp 1667941163
transform 1 0 19504 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_208
timestamp 1667941163
transform 1 0 20240 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_216
timestamp 1667941163
transform 1 0 20976 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1667941163
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_234
timestamp 1667941163
transform 1 0 22632 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_246
timestamp 1667941163
transform 1 0 23736 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_258
timestamp 1667941163
transform 1 0 24840 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_268
timestamp 1667941163
transform 1 0 25760 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_297
timestamp 1667941163
transform 1 0 28428 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_302
timestamp 1667941163
transform 1 0 28888 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_314
timestamp 1667941163
transform 1 0 29992 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_320
timestamp 1667941163
transform 1 0 30544 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1667941163
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1667941163
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_345
timestamp 1667941163
transform 1 0 32844 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_353
timestamp 1667941163
transform 1 0 33580 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_361
timestamp 1667941163
transform 1 0 34316 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_368
timestamp 1667941163
transform 1 0 34960 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_376
timestamp 1667941163
transform 1 0 35696 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1667941163
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1667941163
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_398
timestamp 1667941163
transform 1 0 37720 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_410
timestamp 1667941163
transform 1 0 38824 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_422
timestamp 1667941163
transform 1 0 39928 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_434
timestamp 1667941163
transform 1 0 41032 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_446
timestamp 1667941163
transform 1 0 42136 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1667941163
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1667941163
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1667941163
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1667941163
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1667941163
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1667941163
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_505
timestamp 1667941163
transform 1 0 47564 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_513
timestamp 1667941163
transform 1 0 48300 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_11
timestamp 1667941163
transform 1 0 2116 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1667941163
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1667941163
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1667941163
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1667941163
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1667941163
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1667941163
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1667941163
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1667941163
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1667941163
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1667941163
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1667941163
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1667941163
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1667941163
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_165
timestamp 1667941163
transform 1 0 16284 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_180
timestamp 1667941163
transform 1 0 17664 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_187
timestamp 1667941163
transform 1 0 18308 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1667941163
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_201
timestamp 1667941163
transform 1 0 19596 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1667941163
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1667941163
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_233
timestamp 1667941163
transform 1 0 22540 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_237
timestamp 1667941163
transform 1 0 22908 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_247
timestamp 1667941163
transform 1 0 23828 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1667941163
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_261
timestamp 1667941163
transform 1 0 25116 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_268
timestamp 1667941163
transform 1 0 25760 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_278
timestamp 1667941163
transform 1 0 26680 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_290
timestamp 1667941163
transform 1 0 27784 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_296
timestamp 1667941163
transform 1 0 28336 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_305
timestamp 1667941163
transform 1 0 29164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_315
timestamp 1667941163
transform 1 0 30084 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_324
timestamp 1667941163
transform 1 0 30912 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_336
timestamp 1667941163
transform 1 0 32016 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_348
timestamp 1667941163
transform 1 0 33120 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_360
timestamp 1667941163
transform 1 0 34224 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_374
timestamp 1667941163
transform 1 0 35512 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_385
timestamp 1667941163
transform 1 0 36524 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_393
timestamp 1667941163
transform 1 0 37260 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_402
timestamp 1667941163
transform 1 0 38088 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_414
timestamp 1667941163
transform 1 0 39192 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1667941163
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1667941163
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1667941163
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1667941163
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1667941163
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1667941163
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1667941163
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_489
timestamp 1667941163
transform 1 0 46092 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_514
timestamp 1667941163
transform 1 0 48392 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1667941163
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1667941163
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1667941163
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1667941163
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1667941163
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1667941163
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1667941163
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1667941163
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1667941163
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1667941163
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1667941163
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1667941163
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1667941163
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1667941163
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1667941163
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_179
timestamp 1667941163
transform 1 0 17572 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_191
timestamp 1667941163
transform 1 0 18676 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_203
timestamp 1667941163
transform 1 0 19780 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_215
timestamp 1667941163
transform 1 0 20884 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1667941163
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_237
timestamp 1667941163
transform 1 0 22908 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1667941163
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_261
timestamp 1667941163
transform 1 0 25116 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1667941163
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_305
timestamp 1667941163
transform 1 0 29164 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_313
timestamp 1667941163
transform 1 0 29900 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_330
timestamp 1667941163
transform 1 0 31464 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_354
timestamp 1667941163
transform 1 0 33672 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_366
timestamp 1667941163
transform 1 0 34776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_370
timestamp 1667941163
transform 1 0 35144 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_379
timestamp 1667941163
transform 1 0 35972 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_388
timestamp 1667941163
transform 1 0 36800 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_413
timestamp 1667941163
transform 1 0 39100 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_425
timestamp 1667941163
transform 1 0 40204 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_437
timestamp 1667941163
transform 1 0 41308 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_445
timestamp 1667941163
transform 1 0 42044 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1667941163
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1667941163
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1667941163
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_485
timestamp 1667941163
transform 1 0 45724 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_491
timestamp 1667941163
transform 1 0 46276 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_495
timestamp 1667941163
transform 1 0 46644 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_502
timestamp 1667941163
transform 1 0 47288 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_505
timestamp 1667941163
transform 1 0 47564 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_510
timestamp 1667941163
transform 1 0 48024 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1667941163
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1667941163
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1667941163
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1667941163
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1667941163
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1667941163
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1667941163
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1667941163
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1667941163
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1667941163
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1667941163
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1667941163
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_153
timestamp 1667941163
transform 1 0 15180 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_161
timestamp 1667941163
transform 1 0 15916 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_180
timestamp 1667941163
transform 1 0 17664 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_192
timestamp 1667941163
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_203
timestamp 1667941163
transform 1 0 19780 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_208
timestamp 1667941163
transform 1 0 20240 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_224
timestamp 1667941163
transform 1 0 21712 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_232
timestamp 1667941163
transform 1 0 22448 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1667941163
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_265
timestamp 1667941163
transform 1 0 25484 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_279
timestamp 1667941163
transform 1 0 26772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_287
timestamp 1667941163
transform 1 0 27508 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_293
timestamp 1667941163
transform 1 0 28060 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_300
timestamp 1667941163
transform 1 0 28704 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_321
timestamp 1667941163
transform 1 0 30636 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_327
timestamp 1667941163
transform 1 0 31188 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_344
timestamp 1667941163
transform 1 0 32752 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_354
timestamp 1667941163
transform 1 0 33672 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_362
timestamp 1667941163
transform 1 0 34408 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_385
timestamp 1667941163
transform 1 0 36524 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_393
timestamp 1667941163
transform 1 0 37260 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1667941163
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1667941163
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1667941163
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1667941163
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1667941163
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1667941163
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1667941163
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1667941163
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1667941163
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_489
timestamp 1667941163
transform 1 0 46092 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_514
timestamp 1667941163
transform 1 0 48392 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_11
timestamp 1667941163
transform 1 0 2116 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_16
timestamp 1667941163
transform 1 0 2576 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_28
timestamp 1667941163
transform 1 0 3680 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_40
timestamp 1667941163
transform 1 0 4784 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1667941163
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1667941163
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1667941163
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1667941163
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1667941163
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_125
timestamp 1667941163
transform 1 0 12604 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_147
timestamp 1667941163
transform 1 0 14628 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_159
timestamp 1667941163
transform 1 0 15732 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1667941163
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1667941163
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_193
timestamp 1667941163
transform 1 0 18860 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_202
timestamp 1667941163
transform 1 0 19688 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1667941163
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_237
timestamp 1667941163
transform 1 0 22908 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_246
timestamp 1667941163
transform 1 0 23736 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_258
timestamp 1667941163
transform 1 0 24840 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_266
timestamp 1667941163
transform 1 0 25576 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 1667941163
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1667941163
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_305
timestamp 1667941163
transform 1 0 29164 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_319
timestamp 1667941163
transform 1 0 30452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_331
timestamp 1667941163
transform 1 0 31556 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1667941163
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_345
timestamp 1667941163
transform 1 0 32844 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_350
timestamp 1667941163
transform 1 0 33304 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_360
timestamp 1667941163
transform 1 0 34224 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_372
timestamp 1667941163
transform 1 0 35328 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_384
timestamp 1667941163
transform 1 0 36432 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_417
timestamp 1667941163
transform 1 0 39468 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_425
timestamp 1667941163
transform 1 0 40204 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_435
timestamp 1667941163
transform 1 0 41124 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1667941163
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1667941163
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1667941163
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1667941163
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1667941163
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1667941163
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1667941163
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_505
timestamp 1667941163
transform 1 0 47564 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_510
timestamp 1667941163
transform 1 0 48024 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1667941163
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_41
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_45
timestamp 1667941163
transform 1 0 5244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_57
timestamp 1667941163
transform 1 0 6348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_69
timestamp 1667941163
transform 1 0 7452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 1667941163
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1667941163
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1667941163
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1667941163
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_133
timestamp 1667941163
transform 1 0 13340 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1667941163
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_153
timestamp 1667941163
transform 1 0 15180 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_161
timestamp 1667941163
transform 1 0 15916 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_172
timestamp 1667941163
transform 1 0 16928 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_184
timestamp 1667941163
transform 1 0 18032 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_193
timestamp 1667941163
transform 1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_208
timestamp 1667941163
transform 1 0 20240 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_214
timestamp 1667941163
transform 1 0 20792 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1667941163
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1667941163
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1667941163
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1667941163
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_281
timestamp 1667941163
transform 1 0 26956 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_293
timestamp 1667941163
transform 1 0 28060 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_305
timestamp 1667941163
transform 1 0 29164 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_319
timestamp 1667941163
transform 1 0 30452 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_329
timestamp 1667941163
transform 1 0 31372 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_341
timestamp 1667941163
transform 1 0 32476 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_351
timestamp 1667941163
transform 1 0 33396 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_358
timestamp 1667941163
transform 1 0 34040 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_374
timestamp 1667941163
transform 1 0 35512 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_382
timestamp 1667941163
transform 1 0 36248 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_387
timestamp 1667941163
transform 1 0 36708 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_399
timestamp 1667941163
transform 1 0 37812 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_411
timestamp 1667941163
transform 1 0 38916 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1667941163
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_421
timestamp 1667941163
transform 1 0 39836 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_441
timestamp 1667941163
transform 1 0 41676 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_453
timestamp 1667941163
transform 1 0 42780 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_457
timestamp 1667941163
transform 1 0 43148 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_474
timestamp 1667941163
transform 1 0 44712 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1667941163
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_489
timestamp 1667941163
transform 1 0 46092 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_514
timestamp 1667941163
transform 1 0 48392 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_14
timestamp 1667941163
transform 1 0 2392 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_26
timestamp 1667941163
transform 1 0 3496 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_32
timestamp 1667941163
transform 1 0 4048 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1667941163
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1667941163
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1667941163
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1667941163
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1667941163
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1667941163
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1667941163
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_137
timestamp 1667941163
transform 1 0 13708 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_141
timestamp 1667941163
transform 1 0 14076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_145
timestamp 1667941163
transform 1 0 14444 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_157
timestamp 1667941163
transform 1 0 15548 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_165
timestamp 1667941163
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_177
timestamp 1667941163
transform 1 0 17388 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_194
timestamp 1667941163
transform 1 0 18952 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_202
timestamp 1667941163
transform 1 0 19688 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_207
timestamp 1667941163
transform 1 0 20148 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_216
timestamp 1667941163
transform 1 0 20976 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1667941163
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_265
timestamp 1667941163
transform 1 0 25484 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_269
timestamp 1667941163
transform 1 0 25852 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_276
timestamp 1667941163
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_293
timestamp 1667941163
transform 1 0 28060 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_299
timestamp 1667941163
transform 1 0 28612 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_316
timestamp 1667941163
transform 1 0 30176 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_328
timestamp 1667941163
transform 1 0 31280 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_355
timestamp 1667941163
transform 1 0 33764 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_367
timestamp 1667941163
transform 1 0 34868 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_376
timestamp 1667941163
transform 1 0 35696 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_384
timestamp 1667941163
transform 1 0 36432 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_389
timestamp 1667941163
transform 1 0 36892 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_400
timestamp 1667941163
transform 1 0 37904 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_412
timestamp 1667941163
transform 1 0 39008 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_431
timestamp 1667941163
transform 1 0 40756 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_442
timestamp 1667941163
transform 1 0 41768 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_23_449
timestamp 1667941163
transform 1 0 42412 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_459
timestamp 1667941163
transform 1 0 43332 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_471
timestamp 1667941163
transform 1 0 44436 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_480
timestamp 1667941163
transform 1 0 45264 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_492
timestamp 1667941163
transform 1 0 46368 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_505
timestamp 1667941163
transform 1 0 47564 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_510
timestamp 1667941163
transform 1 0 48024 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1667941163
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1667941163
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_40
timestamp 1667941163
transform 1 0 4784 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_52
timestamp 1667941163
transform 1 0 5888 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_64
timestamp 1667941163
transform 1 0 6992 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_76
timestamp 1667941163
transform 1 0 8096 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1667941163
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1667941163
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1667941163
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_133
timestamp 1667941163
transform 1 0 13340 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1667941163
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_145
timestamp 1667941163
transform 1 0 14444 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_152
timestamp 1667941163
transform 1 0 15088 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_163
timestamp 1667941163
transform 1 0 16100 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_175
timestamp 1667941163
transform 1 0 17204 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_181
timestamp 1667941163
transform 1 0 17756 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_188
timestamp 1667941163
transform 1 0 18400 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_209
timestamp 1667941163
transform 1 0 20332 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_217
timestamp 1667941163
transform 1 0 21068 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_224
timestamp 1667941163
transform 1 0 21712 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_236
timestamp 1667941163
transform 1 0 22816 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_240
timestamp 1667941163
transform 1 0 23184 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_247
timestamp 1667941163
transform 1 0 23828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1667941163
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_258
timestamp 1667941163
transform 1 0 24840 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_265
timestamp 1667941163
transform 1 0 25484 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_287
timestamp 1667941163
transform 1 0 27508 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_299
timestamp 1667941163
transform 1 0 28612 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1667941163
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_315
timestamp 1667941163
transform 1 0 30084 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_324
timestamp 1667941163
transform 1 0 30912 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_334
timestamp 1667941163
transform 1 0 31832 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_343
timestamp 1667941163
transform 1 0 32660 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_351
timestamp 1667941163
transform 1 0 33396 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_362
timestamp 1667941163
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_373
timestamp 1667941163
transform 1 0 35420 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_389
timestamp 1667941163
transform 1 0 36892 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_400
timestamp 1667941163
transform 1 0 37904 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_407
timestamp 1667941163
transform 1 0 38548 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1667941163
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_421
timestamp 1667941163
transform 1 0 39836 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_427
timestamp 1667941163
transform 1 0 40388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_439
timestamp 1667941163
transform 1 0 41492 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_447
timestamp 1667941163
transform 1 0 42228 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_453
timestamp 1667941163
transform 1 0 42780 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_457
timestamp 1667941163
transform 1 0 43148 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_462
timestamp 1667941163
transform 1 0 43608 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_471
timestamp 1667941163
transform 1 0 44436 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1667941163
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_477
timestamp 1667941163
transform 1 0 44988 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_483
timestamp 1667941163
transform 1 0 45540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_495
timestamp 1667941163
transform 1 0 46644 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_503
timestamp 1667941163
transform 1 0 47380 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_507
timestamp 1667941163
transform 1 0 47748 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_515
timestamp 1667941163
transform 1 0 48484 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1667941163
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1667941163
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1667941163
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1667941163
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1667941163
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1667941163
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1667941163
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1667941163
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1667941163
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1667941163
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1667941163
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_137
timestamp 1667941163
transform 1 0 13708 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_145
timestamp 1667941163
transform 1 0 14444 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_152
timestamp 1667941163
transform 1 0 15088 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1667941163
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_174
timestamp 1667941163
transform 1 0 17112 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_186
timestamp 1667941163
transform 1 0 18216 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_198
timestamp 1667941163
transform 1 0 19320 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_206
timestamp 1667941163
transform 1 0 20056 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_214
timestamp 1667941163
transform 1 0 20792 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1667941163
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_233
timestamp 1667941163
transform 1 0 22540 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_244
timestamp 1667941163
transform 1 0 23552 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_255
timestamp 1667941163
transform 1 0 24564 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_265
timestamp 1667941163
transform 1 0 25484 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_271
timestamp 1667941163
transform 1 0 26036 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1667941163
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_291
timestamp 1667941163
transform 1 0 27876 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_295
timestamp 1667941163
transform 1 0 28244 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_312
timestamp 1667941163
transform 1 0 29808 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_320
timestamp 1667941163
transform 1 0 30544 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_334
timestamp 1667941163
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_355
timestamp 1667941163
transform 1 0 33764 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_375
timestamp 1667941163
transform 1 0 35604 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_384
timestamp 1667941163
transform 1 0 36432 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_399
timestamp 1667941163
transform 1 0 37812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_411
timestamp 1667941163
transform 1 0 38916 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_419
timestamp 1667941163
transform 1 0 39652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_428
timestamp 1667941163
transform 1 0 40480 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_438
timestamp 1667941163
transform 1 0 41400 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_446
timestamp 1667941163
transform 1 0 42136 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1667941163
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_461
timestamp 1667941163
transform 1 0 43516 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_474
timestamp 1667941163
transform 1 0 44712 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_485
timestamp 1667941163
transform 1 0 45724 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_496
timestamp 1667941163
transform 1 0 46736 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_505
timestamp 1667941163
transform 1 0 47564 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_513
timestamp 1667941163
transform 1 0 48300 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_14
timestamp 1667941163
transform 1 0 2392 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1667941163
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1667941163
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1667941163
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1667941163
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1667941163
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1667941163
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1667941163
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1667941163
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1667941163
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1667941163
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1667941163
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1667941163
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_147
timestamp 1667941163
transform 1 0 14628 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_151
timestamp 1667941163
transform 1 0 14996 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_157
timestamp 1667941163
transform 1 0 15548 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_163
timestamp 1667941163
transform 1 0 16100 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_172
timestamp 1667941163
transform 1 0 16928 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_184
timestamp 1667941163
transform 1 0 18032 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1667941163
transform 1 0 20884 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_226
timestamp 1667941163
transform 1 0 21896 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_238
timestamp 1667941163
transform 1 0 23000 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_244
timestamp 1667941163
transform 1 0 23552 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_259
timestamp 1667941163
transform 1 0 24932 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_267
timestamp 1667941163
transform 1 0 25668 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_279
timestamp 1667941163
transform 1 0 26772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_291
timestamp 1667941163
transform 1 0 27876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_303
timestamp 1667941163
transform 1 0 28980 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1667941163
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_319
timestamp 1667941163
transform 1 0 30452 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_331
timestamp 1667941163
transform 1 0 31556 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_343
timestamp 1667941163
transform 1 0 32660 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_355
timestamp 1667941163
transform 1 0 33764 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1667941163
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_383
timestamp 1667941163
transform 1 0 36340 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_398
timestamp 1667941163
transform 1 0 37720 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_418
timestamp 1667941163
transform 1 0 39560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_421
timestamp 1667941163
transform 1 0 39836 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_431
timestamp 1667941163
transform 1 0 40756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_451
timestamp 1667941163
transform 1 0 42596 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_461
timestamp 1667941163
transform 1 0 43516 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_473
timestamp 1667941163
transform 1 0 44620 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_477
timestamp 1667941163
transform 1 0 44988 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_482
timestamp 1667941163
transform 1 0 45448 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_488
timestamp 1667941163
transform 1 0 46000 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_505
timestamp 1667941163
transform 1 0 47564 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_513
timestamp 1667941163
transform 1 0 48300 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_9
timestamp 1667941163
transform 1 0 1932 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_31
timestamp 1667941163
transform 1 0 3956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_43
timestamp 1667941163
transform 1 0 5060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1667941163
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1667941163
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1667941163
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1667941163
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1667941163
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1667941163
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_133
timestamp 1667941163
transform 1 0 13340 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_145
timestamp 1667941163
transform 1 0 14444 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_153
timestamp 1667941163
transform 1 0 15180 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1667941163
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_180
timestamp 1667941163
transform 1 0 17664 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_190
timestamp 1667941163
transform 1 0 18584 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_202
timestamp 1667941163
transform 1 0 19688 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1667941163
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_237
timestamp 1667941163
transform 1 0 22908 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_243
timestamp 1667941163
transform 1 0 23460 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_255
timestamp 1667941163
transform 1 0 24564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_267
timestamp 1667941163
transform 1 0 25668 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1667941163
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_293
timestamp 1667941163
transform 1 0 28060 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_299
timestamp 1667941163
transform 1 0 28612 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_316
timestamp 1667941163
transform 1 0 30176 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_328
timestamp 1667941163
transform 1 0 31280 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_346
timestamp 1667941163
transform 1 0 32936 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_358
timestamp 1667941163
transform 1 0 34040 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_366
timestamp 1667941163
transform 1 0 34776 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_370
timestamp 1667941163
transform 1 0 35144 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_382
timestamp 1667941163
transform 1 0 36248 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_390
timestamp 1667941163
transform 1 0 36984 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1667941163
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_429
timestamp 1667941163
transform 1 0 40572 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_438
timestamp 1667941163
transform 1 0 41400 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_446
timestamp 1667941163
transform 1 0 42136 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_449
timestamp 1667941163
transform 1 0 42412 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_457
timestamp 1667941163
transform 1 0 43148 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1667941163
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1667941163
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1667941163
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1667941163
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_505
timestamp 1667941163
transform 1 0 47564 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_510
timestamp 1667941163
transform 1 0 48024 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_11
timestamp 1667941163
transform 1 0 2116 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1667941163
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1667941163
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1667941163
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1667941163
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1667941163
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1667941163
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1667941163
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1667941163
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_109
timestamp 1667941163
transform 1 0 11132 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_117
timestamp 1667941163
transform 1 0 11868 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp 1667941163
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_151
timestamp 1667941163
transform 1 0 14996 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_158
timestamp 1667941163
transform 1 0 15640 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_170
timestamp 1667941163
transform 1 0 16744 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_190
timestamp 1667941163
transform 1 0 18584 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_205
timestamp 1667941163
transform 1 0 19964 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_225
timestamp 1667941163
transform 1 0 21804 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_233
timestamp 1667941163
transform 1 0 22540 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_242
timestamp 1667941163
transform 1 0 23368 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_249
timestamp 1667941163
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1667941163
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1667941163
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_289
timestamp 1667941163
transform 1 0 27692 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_297
timestamp 1667941163
transform 1 0 28428 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_306
timestamp 1667941163
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_319
timestamp 1667941163
transform 1 0 30452 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_323
timestamp 1667941163
transform 1 0 30820 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_330
timestamp 1667941163
transform 1 0 31464 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_350
timestamp 1667941163
transform 1 0 33304 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_362
timestamp 1667941163
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_372
timestamp 1667941163
transform 1 0 35328 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_380
timestamp 1667941163
transform 1 0 36064 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_387
timestamp 1667941163
transform 1 0 36708 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_399
timestamp 1667941163
transform 1 0 37812 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_411
timestamp 1667941163
transform 1 0 38916 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1667941163
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_421
timestamp 1667941163
transform 1 0 39836 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_429
timestamp 1667941163
transform 1 0 40572 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_440
timestamp 1667941163
transform 1 0 41584 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_452
timestamp 1667941163
transform 1 0 42688 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1667941163
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1667941163
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_477
timestamp 1667941163
transform 1 0 44988 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_483
timestamp 1667941163
transform 1 0 45540 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_491
timestamp 1667941163
transform 1 0 46276 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_514
timestamp 1667941163
transform 1 0 48392 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_9
timestamp 1667941163
transform 1 0 1932 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_31
timestamp 1667941163
transform 1 0 3956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_43
timestamp 1667941163
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1667941163
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1667941163
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1667941163
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1667941163
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1667941163
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1667941163
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_119
timestamp 1667941163
transform 1 0 12052 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_126
timestamp 1667941163
transform 1 0 12696 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_138
timestamp 1667941163
transform 1 0 13800 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_150
timestamp 1667941163
transform 1 0 14904 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_162
timestamp 1667941163
transform 1 0 16008 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1667941163
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1667941163
transform 1 0 17756 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_190
timestamp 1667941163
transform 1 0 18584 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_202
timestamp 1667941163
transform 1 0 19688 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_213
timestamp 1667941163
transform 1 0 20700 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_221
timestamp 1667941163
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_237
timestamp 1667941163
transform 1 0 22908 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_243
timestamp 1667941163
transform 1 0 23460 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_249
timestamp 1667941163
transform 1 0 24012 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_256
timestamp 1667941163
transform 1 0 24656 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_268
timestamp 1667941163
transform 1 0 25760 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_291
timestamp 1667941163
transform 1 0 27876 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_303
timestamp 1667941163
transform 1 0 28980 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_315
timestamp 1667941163
transform 1 0 30084 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_325
timestamp 1667941163
transform 1 0 31004 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_333
timestamp 1667941163
transform 1 0 31740 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_358
timestamp 1667941163
transform 1 0 34040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_368
timestamp 1667941163
transform 1 0 34960 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_379
timestamp 1667941163
transform 1 0 35972 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_390
timestamp 1667941163
transform 1 0 36984 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_411
timestamp 1667941163
transform 1 0 38916 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_428
timestamp 1667941163
transform 1 0 40480 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_434
timestamp 1667941163
transform 1 0 41032 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_439
timestamp 1667941163
transform 1 0 41492 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1667941163
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1667941163
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_461
timestamp 1667941163
transform 1 0 43516 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_469
timestamp 1667941163
transform 1 0 44252 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_489
timestamp 1667941163
transform 1 0 46092 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_501
timestamp 1667941163
transform 1 0 47196 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_505
timestamp 1667941163
transform 1 0 47564 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_510
timestamp 1667941163
transform 1 0 48024 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_9
timestamp 1667941163
transform 1 0 1932 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_13
timestamp 1667941163
transform 1 0 2300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_25
timestamp 1667941163
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1667941163
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1667941163
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1667941163
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1667941163
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1667941163
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1667941163
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1667941163
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1667941163
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1667941163
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1667941163
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_153
timestamp 1667941163
transform 1 0 15180 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_159
timestamp 1667941163
transform 1 0 15732 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1667941163
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1667941163
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1667941163
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_215
timestamp 1667941163
transform 1 0 20884 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_237
timestamp 1667941163
transform 1 0 22908 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1667941163
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_263
timestamp 1667941163
transform 1 0 25300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_291
timestamp 1667941163
transform 1 0 27876 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1667941163
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1667941163
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_315
timestamp 1667941163
transform 1 0 30084 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_332
timestamp 1667941163
transform 1 0 31648 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_347
timestamp 1667941163
transform 1 0 33028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_359
timestamp 1667941163
transform 1 0 34132 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1667941163
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_375
timestamp 1667941163
transform 1 0 35604 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_386
timestamp 1667941163
transform 1 0 36616 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_394
timestamp 1667941163
transform 1 0 37352 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_408
timestamp 1667941163
transform 1 0 38640 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_414
timestamp 1667941163
transform 1 0 39192 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_418
timestamp 1667941163
transform 1 0 39560 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_421
timestamp 1667941163
transform 1 0 39836 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_432
timestamp 1667941163
transform 1 0 40848 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_441
timestamp 1667941163
transform 1 0 41676 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_448
timestamp 1667941163
transform 1 0 42320 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_460
timestamp 1667941163
transform 1 0 43424 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_464
timestamp 1667941163
transform 1 0 43792 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_473
timestamp 1667941163
transform 1 0 44620 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_477
timestamp 1667941163
transform 1 0 44988 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_487
timestamp 1667941163
transform 1 0 45908 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_514
timestamp 1667941163
transform 1 0 48392 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1667941163
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1667941163
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1667941163
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1667941163
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1667941163
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1667941163
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1667941163
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1667941163
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1667941163
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_125
timestamp 1667941163
transform 1 0 12604 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_135
timestamp 1667941163
transform 1 0 13524 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_156
timestamp 1667941163
transform 1 0 15456 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_165
timestamp 1667941163
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_179
timestamp 1667941163
transform 1 0 17572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_191
timestamp 1667941163
transform 1 0 18676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_203
timestamp 1667941163
transform 1 0 19780 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1667941163
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_233
timestamp 1667941163
transform 1 0 22540 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_241
timestamp 1667941163
transform 1 0 23276 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_258
timestamp 1667941163
transform 1 0 24840 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1667941163
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_289
timestamp 1667941163
transform 1 0 27692 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_31_313
timestamp 1667941163
transform 1 0 29900 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_325
timestamp 1667941163
transform 1 0 31004 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_333
timestamp 1667941163
transform 1 0 31740 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_347
timestamp 1667941163
transform 1 0 33028 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_358
timestamp 1667941163
transform 1 0 34040 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_368
timestamp 1667941163
transform 1 0 34960 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_380
timestamp 1667941163
transform 1 0 36064 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_397
timestamp 1667941163
transform 1 0 37628 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_414
timestamp 1667941163
transform 1 0 39192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_426
timestamp 1667941163
transform 1 0 40296 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_436
timestamp 1667941163
transform 1 0 41216 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_445
timestamp 1667941163
transform 1 0 42044 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_449
timestamp 1667941163
transform 1 0 42412 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_457
timestamp 1667941163
transform 1 0 43148 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_463
timestamp 1667941163
transform 1 0 43700 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_471
timestamp 1667941163
transform 1 0 44436 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_478
timestamp 1667941163
transform 1 0 45080 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_490
timestamp 1667941163
transform 1 0 46184 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_498
timestamp 1667941163
transform 1 0 46920 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_502
timestamp 1667941163
transform 1 0 47288 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_505
timestamp 1667941163
transform 1 0 47564 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_510
timestamp 1667941163
transform 1 0 48024 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_11
timestamp 1667941163
transform 1 0 2116 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_16
timestamp 1667941163
transform 1 0 2576 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1667941163
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1667941163
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1667941163
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1667941163
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1667941163
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1667941163
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_109
timestamp 1667941163
transform 1 0 11132 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1667941163
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1667941163
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_159
timestamp 1667941163
transform 1 0 15732 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_176
timestamp 1667941163
transform 1 0 17296 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_183
timestamp 1667941163
transform 1 0 17940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1667941163
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_201
timestamp 1667941163
transform 1 0 19596 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_210
timestamp 1667941163
transform 1 0 20424 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_222
timestamp 1667941163
transform 1 0 21528 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1667941163
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1667941163
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1667941163
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_265
timestamp 1667941163
transform 1 0 25484 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_275
timestamp 1667941163
transform 1 0 26404 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_287
timestamp 1667941163
transform 1 0 27508 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_299
timestamp 1667941163
transform 1 0 28612 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1667941163
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_319
timestamp 1667941163
transform 1 0 30452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_331
timestamp 1667941163
transform 1 0 31556 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_348
timestamp 1667941163
transform 1 0 33120 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_352
timestamp 1667941163
transform 1 0 33488 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1667941163
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1667941163
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_371
timestamp 1667941163
transform 1 0 35236 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_375
timestamp 1667941163
transform 1 0 35604 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_387
timestamp 1667941163
transform 1 0 36708 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_399
timestamp 1667941163
transform 1 0 37812 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_411
timestamp 1667941163
transform 1 0 38916 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_418
timestamp 1667941163
transform 1 0 39560 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_421
timestamp 1667941163
transform 1 0 39836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_431
timestamp 1667941163
transform 1 0 40756 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_442
timestamp 1667941163
transform 1 0 41768 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_454
timestamp 1667941163
transform 1 0 42872 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_466
timestamp 1667941163
transform 1 0 43976 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_474
timestamp 1667941163
transform 1 0 44712 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1667941163
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_489
timestamp 1667941163
transform 1 0 46092 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_514
timestamp 1667941163
transform 1 0 48392 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_9
timestamp 1667941163
transform 1 0 1932 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_31
timestamp 1667941163
transform 1 0 3956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_43
timestamp 1667941163
transform 1 0 5060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1667941163
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1667941163
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1667941163
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1667941163
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1667941163
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1667941163
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_121
timestamp 1667941163
transform 1 0 12236 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_128
timestamp 1667941163
transform 1 0 12880 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_140
timestamp 1667941163
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_144
timestamp 1667941163
transform 1 0 14352 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_155
timestamp 1667941163
transform 1 0 15364 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1667941163
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_178
timestamp 1667941163
transform 1 0 17480 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_186
timestamp 1667941163
transform 1 0 18216 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_194
timestamp 1667941163
transform 1 0 18952 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_213
timestamp 1667941163
transform 1 0 20700 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_221
timestamp 1667941163
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_231
timestamp 1667941163
transform 1 0 22356 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_243
timestamp 1667941163
transform 1 0 23460 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_255
timestamp 1667941163
transform 1 0 24564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_267
timestamp 1667941163
transform 1 0 25668 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1667941163
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1667941163
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_305
timestamp 1667941163
transform 1 0 29164 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_313
timestamp 1667941163
transform 1 0 29900 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_325
timestamp 1667941163
transform 1 0 31004 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_333
timestamp 1667941163
transform 1 0 31740 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_353
timestamp 1667941163
transform 1 0 33580 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_358
timestamp 1667941163
transform 1 0 34040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_367
timestamp 1667941163
transform 1 0 34868 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_382
timestamp 1667941163
transform 1 0 36248 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_390
timestamp 1667941163
transform 1 0 36984 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_405
timestamp 1667941163
transform 1 0 38364 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_429
timestamp 1667941163
transform 1 0 40572 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_446
timestamp 1667941163
transform 1 0 42136 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1667941163
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_461
timestamp 1667941163
transform 1 0 43516 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_471
timestamp 1667941163
transform 1 0 44436 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_483
timestamp 1667941163
transform 1 0 45540 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_489
timestamp 1667941163
transform 1 0 46092 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_493
timestamp 1667941163
transform 1 0 46460 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_500
timestamp 1667941163
transform 1 0 47104 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_505
timestamp 1667941163
transform 1 0 47564 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_513
timestamp 1667941163
transform 1 0 48300 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_14
timestamp 1667941163
transform 1 0 2392 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1667941163
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1667941163
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1667941163
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1667941163
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1667941163
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1667941163
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1667941163
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1667941163
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1667941163
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1667941163
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1667941163
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_151
timestamp 1667941163
transform 1 0 14996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_166
timestamp 1667941163
transform 1 0 16376 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1667941163
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1667941163
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1667941163
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_207
timestamp 1667941163
transform 1 0 20148 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_219
timestamp 1667941163
transform 1 0 21252 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_231
timestamp 1667941163
transform 1 0 22356 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1667941163
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1667941163
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_261
timestamp 1667941163
transform 1 0 25116 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_268
timestamp 1667941163
transform 1 0 25760 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_278
timestamp 1667941163
transform 1 0 26680 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_287
timestamp 1667941163
transform 1 0 27508 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_295
timestamp 1667941163
transform 1 0 28244 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_303
timestamp 1667941163
transform 1 0 28980 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1667941163
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_313
timestamp 1667941163
transform 1 0 29900 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_322
timestamp 1667941163
transform 1 0 30728 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_334
timestamp 1667941163
transform 1 0 31832 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_346
timestamp 1667941163
transform 1 0 32936 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_358
timestamp 1667941163
transform 1 0 34040 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_373
timestamp 1667941163
transform 1 0 35420 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_390
timestamp 1667941163
transform 1 0 36984 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_402
timestamp 1667941163
transform 1 0 38088 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_414
timestamp 1667941163
transform 1 0 39192 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1667941163
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1667941163
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1667941163
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_457
timestamp 1667941163
transform 1 0 43148 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_474
timestamp 1667941163
transform 1 0 44712 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1667941163
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_489
timestamp 1667941163
transform 1 0 46092 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_514
timestamp 1667941163
transform 1 0 48392 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_14
timestamp 1667941163
transform 1 0 2392 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_26
timestamp 1667941163
transform 1 0 3496 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_38
timestamp 1667941163
transform 1 0 4600 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_50
timestamp 1667941163
transform 1 0 5704 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1667941163
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1667941163
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1667941163
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1667941163
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1667941163
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_125
timestamp 1667941163
transform 1 0 12604 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_131
timestamp 1667941163
transform 1 0 13156 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_148
timestamp 1667941163
transform 1 0 14720 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_160
timestamp 1667941163
transform 1 0 15824 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1667941163
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_178
timestamp 1667941163
transform 1 0 17480 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_188
timestamp 1667941163
transform 1 0 18400 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_200
timestamp 1667941163
transform 1 0 19504 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_212
timestamp 1667941163
transform 1 0 20608 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_229
timestamp 1667941163
transform 1 0 22172 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_246
timestamp 1667941163
transform 1 0 23736 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_256
timestamp 1667941163
transform 1 0 24656 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_260
timestamp 1667941163
transform 1 0 25024 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_267
timestamp 1667941163
transform 1 0 25668 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_273
timestamp 1667941163
transform 1 0 26220 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1667941163
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_289
timestamp 1667941163
transform 1 0 27692 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_297
timestamp 1667941163
transform 1 0 28428 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_303
timestamp 1667941163
transform 1 0 28980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_325
timestamp 1667941163
transform 1 0 31004 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_334
timestamp 1667941163
transform 1 0 31832 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_341
timestamp 1667941163
transform 1 0 32476 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_351
timestamp 1667941163
transform 1 0 33396 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_358
timestamp 1667941163
transform 1 0 34040 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_377
timestamp 1667941163
transform 1 0 35788 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_386
timestamp 1667941163
transform 1 0 36616 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_401
timestamp 1667941163
transform 1 0 37996 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_413
timestamp 1667941163
transform 1 0 39100 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_425
timestamp 1667941163
transform 1 0 40204 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_437
timestamp 1667941163
transform 1 0 41308 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_445
timestamp 1667941163
transform 1 0 42044 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_449
timestamp 1667941163
transform 1 0 42412 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_456
timestamp 1667941163
transform 1 0 43056 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_464
timestamp 1667941163
transform 1 0 43792 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_474
timestamp 1667941163
transform 1 0 44712 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_482
timestamp 1667941163
transform 1 0 45448 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_490
timestamp 1667941163
transform 1 0 46184 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_495
timestamp 1667941163
transform 1 0 46644 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_502
timestamp 1667941163
transform 1 0 47288 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_505
timestamp 1667941163
transform 1 0 47564 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_510
timestamp 1667941163
transform 1 0 48024 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1667941163
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1667941163
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1667941163
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1667941163
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1667941163
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1667941163
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_109
timestamp 1667941163
transform 1 0 11132 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_118
timestamp 1667941163
transform 1 0 11960 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_130
timestamp 1667941163
transform 1 0 13064 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1667941163
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_149
timestamp 1667941163
transform 1 0 14812 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_161
timestamp 1667941163
transform 1 0 15916 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_179
timestamp 1667941163
transform 1 0 17572 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_190
timestamp 1667941163
transform 1 0 18584 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_207
timestamp 1667941163
transform 1 0 20148 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_215
timestamp 1667941163
transform 1 0 20884 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_229
timestamp 1667941163
transform 1 0 22172 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_236
timestamp 1667941163
transform 1 0 22816 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_249
timestamp 1667941163
transform 1 0 24012 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_263
timestamp 1667941163
transform 1 0 25300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_282
timestamp 1667941163
transform 1 0 27048 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_286
timestamp 1667941163
transform 1 0 27416 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_294
timestamp 1667941163
transform 1 0 28152 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_306
timestamp 1667941163
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_317
timestamp 1667941163
transform 1 0 30268 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_323
timestamp 1667941163
transform 1 0 30820 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_340
timestamp 1667941163
transform 1 0 32384 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_360
timestamp 1667941163
transform 1 0 34224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_36_374
timestamp 1667941163
transform 1 0 35512 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_380
timestamp 1667941163
transform 1 0 36064 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_389
timestamp 1667941163
transform 1 0 36892 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_400
timestamp 1667941163
transform 1 0 37904 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_407
timestamp 1667941163
transform 1 0 38548 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_411
timestamp 1667941163
transform 1 0 38916 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_418
timestamp 1667941163
transform 1 0 39560 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_421
timestamp 1667941163
transform 1 0 39836 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_425
timestamp 1667941163
transform 1 0 40204 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_432
timestamp 1667941163
transform 1 0 40848 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_436
timestamp 1667941163
transform 1 0 41216 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_453
timestamp 1667941163
transform 1 0 42780 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_463
timestamp 1667941163
transform 1 0 43700 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_471
timestamp 1667941163
transform 1 0 44436 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1667941163
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1667941163
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_489
timestamp 1667941163
transform 1 0 46092 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_514
timestamp 1667941163
transform 1 0 48392 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_11
timestamp 1667941163
transform 1 0 2116 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_17
timestamp 1667941163
transform 1 0 2668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_29
timestamp 1667941163
transform 1 0 3772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_41
timestamp 1667941163
transform 1 0 4876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_53
timestamp 1667941163
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1667941163
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1667941163
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_105
timestamp 1667941163
transform 1 0 10764 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1667941163
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_131
timestamp 1667941163
transform 1 0 13156 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_143
timestamp 1667941163
transform 1 0 14260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1667941163
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_174
timestamp 1667941163
transform 1 0 17112 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_186
timestamp 1667941163
transform 1 0 18216 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_210
timestamp 1667941163
transform 1 0 20424 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1667941163
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_243
timestamp 1667941163
transform 1 0 23460 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_249
timestamp 1667941163
transform 1 0 24012 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_266
timestamp 1667941163
transform 1 0 25576 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_274
timestamp 1667941163
transform 1 0 26312 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1667941163
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_288
timestamp 1667941163
transform 1 0 27600 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_294
timestamp 1667941163
transform 1 0 28152 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_300
timestamp 1667941163
transform 1 0 28704 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_309
timestamp 1667941163
transform 1 0 29532 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_315
timestamp 1667941163
transform 1 0 30084 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_322
timestamp 1667941163
transform 1 0 30728 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_332
timestamp 1667941163
transform 1 0 31648 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_358
timestamp 1667941163
transform 1 0 34040 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_370
timestamp 1667941163
transform 1 0 35144 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1667941163
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1667941163
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_398
timestamp 1667941163
transform 1 0 37720 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_410
timestamp 1667941163
transform 1 0 38824 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_427
timestamp 1667941163
transform 1 0 40388 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_439
timestamp 1667941163
transform 1 0 41492 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_446
timestamp 1667941163
transform 1 0 42136 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_449
timestamp 1667941163
transform 1 0 42412 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_459
timestamp 1667941163
transform 1 0 43332 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_468
timestamp 1667941163
transform 1 0 44160 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_480
timestamp 1667941163
transform 1 0 45264 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_492
timestamp 1667941163
transform 1 0 46368 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_505
timestamp 1667941163
transform 1 0 47564 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_510
timestamp 1667941163
transform 1 0 48024 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1667941163
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1667941163
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1667941163
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1667941163
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1667941163
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1667941163
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_109
timestamp 1667941163
transform 1 0 11132 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_124
timestamp 1667941163
transform 1 0 12512 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1667941163
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_149
timestamp 1667941163
transform 1 0 14812 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_161
timestamp 1667941163
transform 1 0 15916 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_173
timestamp 1667941163
transform 1 0 17020 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_185
timestamp 1667941163
transform 1 0 18124 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_193
timestamp 1667941163
transform 1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_205
timestamp 1667941163
transform 1 0 19964 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_217
timestamp 1667941163
transform 1 0 21068 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_238
timestamp 1667941163
transform 1 0 23000 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1667941163
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_261
timestamp 1667941163
transform 1 0 25116 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_269
timestamp 1667941163
transform 1 0 25852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_277
timestamp 1667941163
transform 1 0 26588 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_285
timestamp 1667941163
transform 1 0 27324 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_293
timestamp 1667941163
transform 1 0 28060 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_302
timestamp 1667941163
transform 1 0 28888 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_325
timestamp 1667941163
transform 1 0 31004 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_335
timestamp 1667941163
transform 1 0 31924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_353
timestamp 1667941163
transform 1 0 33580 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_361
timestamp 1667941163
transform 1 0 34316 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_373
timestamp 1667941163
transform 1 0 35420 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_381
timestamp 1667941163
transform 1 0 36156 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_388
timestamp 1667941163
transform 1 0 36800 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_399
timestamp 1667941163
transform 1 0 37812 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_411
timestamp 1667941163
transform 1 0 38916 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1667941163
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1667941163
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1667941163
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_445
timestamp 1667941163
transform 1 0 42044 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_455
timestamp 1667941163
transform 1 0 42964 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_467
timestamp 1667941163
transform 1 0 44068 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1667941163
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1667941163
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1667941163
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1667941163
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_513
timestamp 1667941163
transform 1 0 48300 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1667941163
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1667941163
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1667941163
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1667941163
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1667941163
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_62
timestamp 1667941163
transform 1 0 6808 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_74
timestamp 1667941163
transform 1 0 7912 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_82
timestamp 1667941163
transform 1 0 8648 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_87
timestamp 1667941163
transform 1 0 9108 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_102
timestamp 1667941163
transform 1 0 10488 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1667941163
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1667941163
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_137
timestamp 1667941163
transform 1 0 13708 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_156
timestamp 1667941163
transform 1 0 15456 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1667941163
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_193
timestamp 1667941163
transform 1 0 18860 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_213
timestamp 1667941163
transform 1 0 20700 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_221
timestamp 1667941163
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_236
timestamp 1667941163
transform 1 0 22816 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_245
timestamp 1667941163
transform 1 0 23644 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_252
timestamp 1667941163
transform 1 0 24288 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_264
timestamp 1667941163
transform 1 0 25392 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1667941163
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_290
timestamp 1667941163
transform 1 0 27784 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_314
timestamp 1667941163
transform 1 0 29992 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_322
timestamp 1667941163
transform 1 0 30728 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1667941163
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_345
timestamp 1667941163
transform 1 0 32844 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_356
timestamp 1667941163
transform 1 0 33856 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_376
timestamp 1667941163
transform 1 0 35696 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_389
timestamp 1667941163
transform 1 0 36892 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_405
timestamp 1667941163
transform 1 0 38364 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_409
timestamp 1667941163
transform 1 0 38732 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_418
timestamp 1667941163
transform 1 0 39560 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_432
timestamp 1667941163
transform 1 0 40848 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_444
timestamp 1667941163
transform 1 0 41952 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1667941163
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_461
timestamp 1667941163
transform 1 0 43516 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_472
timestamp 1667941163
transform 1 0 44528 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_484
timestamp 1667941163
transform 1 0 45632 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_496
timestamp 1667941163
transform 1 0 46736 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_502
timestamp 1667941163
transform 1 0 47288 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_505
timestamp 1667941163
transform 1 0 47564 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_510
timestamp 1667941163
transform 1 0 48024 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1667941163
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_53
timestamp 1667941163
transform 1 0 5980 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_78
timestamp 1667941163
transform 1 0 8280 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_103
timestamp 1667941163
transform 1 0 10580 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_110
timestamp 1667941163
transform 1 0 11224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_117
timestamp 1667941163
transform 1 0 11868 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_130
timestamp 1667941163
transform 1 0 13064 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1667941163
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_152
timestamp 1667941163
transform 1 0 15088 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_165
timestamp 1667941163
transform 1 0 16284 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_172
timestamp 1667941163
transform 1 0 16928 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_185
timestamp 1667941163
transform 1 0 18124 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_193
timestamp 1667941163
transform 1 0 18860 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1667941163
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_221
timestamp 1667941163
transform 1 0 21436 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_246
timestamp 1667941163
transform 1 0 23736 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_265
timestamp 1667941163
transform 1 0 25484 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_271
timestamp 1667941163
transform 1 0 26036 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_284
timestamp 1667941163
transform 1 0 27232 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_304
timestamp 1667941163
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_321
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_327
timestamp 1667941163
transform 1 0 31188 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_337
timestamp 1667941163
transform 1 0 32108 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_361
timestamp 1667941163
transform 1 0 34316 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_396
timestamp 1667941163
transform 1 0 37536 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_418
timestamp 1667941163
transform 1 0 39560 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1667941163
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_433
timestamp 1667941163
transform 1 0 40940 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_453
timestamp 1667941163
transform 1 0 42780 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_462
timestamp 1667941163
transform 1 0 43608 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_471
timestamp 1667941163
transform 1 0 44436 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1667941163
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1667941163
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_489
timestamp 1667941163
transform 1 0 46092 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_514
timestamp 1667941163
transform 1 0 48392 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_11
timestamp 1667941163
transform 1 0 2116 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_17
timestamp 1667941163
transform 1 0 2668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_29
timestamp 1667941163
transform 1 0 3772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_41
timestamp 1667941163
transform 1 0 4876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_53
timestamp 1667941163
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_65
timestamp 1667941163
transform 1 0 7084 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_72
timestamp 1667941163
transform 1 0 7728 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_92
timestamp 1667941163
transform 1 0 9568 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1667941163
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1667941163
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_131
timestamp 1667941163
transform 1 0 13156 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_140
timestamp 1667941163
transform 1 0 13984 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_160
timestamp 1667941163
transform 1 0 15824 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_176
timestamp 1667941163
transform 1 0 17296 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_183
timestamp 1667941163
transform 1 0 17940 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_190
timestamp 1667941163
transform 1 0 18584 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_198
timestamp 1667941163
transform 1 0 19320 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_206
timestamp 1667941163
transform 1 0 20056 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_218
timestamp 1667941163
transform 1 0 21160 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_230
timestamp 1667941163
transform 1 0 22264 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_238
timestamp 1667941163
transform 1 0 23000 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_248
timestamp 1667941163
transform 1 0 23920 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_260
timestamp 1667941163
transform 1 0 25024 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1667941163
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_287
timestamp 1667941163
transform 1 0 27508 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_295
timestamp 1667941163
transform 1 0 28244 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_318
timestamp 1667941163
transform 1 0 30360 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_330
timestamp 1667941163
transform 1 0 31464 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_348
timestamp 1667941163
transform 1 0 33120 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_352
timestamp 1667941163
transform 1 0 33488 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1667941163
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1667941163
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_415
timestamp 1667941163
transform 1 0 39284 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_427
timestamp 1667941163
transform 1 0 40388 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_439
timestamp 1667941163
transform 1 0 41492 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_446
timestamp 1667941163
transform 1 0 42136 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_449
timestamp 1667941163
transform 1 0 42412 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_41_462
timestamp 1667941163
transform 1 0 43608 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_468
timestamp 1667941163
transform 1 0 44160 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_485
timestamp 1667941163
transform 1 0 45724 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_491
timestamp 1667941163
transform 1 0 46276 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_495
timestamp 1667941163
transform 1 0 46644 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_502
timestamp 1667941163
transform 1 0 47288 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_505
timestamp 1667941163
transform 1 0 47564 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_509
timestamp 1667941163
transform 1 0 47932 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_514
timestamp 1667941163
transform 1 0 48392 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_26
timestamp 1667941163
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_53
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_60
timestamp 1667941163
transform 1 0 6624 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_64
timestamp 1667941163
transform 1 0 6992 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_68
timestamp 1667941163
transform 1 0 7360 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_76
timestamp 1667941163
transform 1 0 8096 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1667941163
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_96
timestamp 1667941163
transform 1 0 9936 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_108
timestamp 1667941163
transform 1 0 11040 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_117
timestamp 1667941163
transform 1 0 11868 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_130
timestamp 1667941163
transform 1 0 13064 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1667941163
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_152
timestamp 1667941163
transform 1 0 15088 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_160
timestamp 1667941163
transform 1 0 15824 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_168
timestamp 1667941163
transform 1 0 16560 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_179
timestamp 1667941163
transform 1 0 17572 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1667941163
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_209
timestamp 1667941163
transform 1 0 20332 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_217
timestamp 1667941163
transform 1 0 21068 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_224
timestamp 1667941163
transform 1 0 21712 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_236
timestamp 1667941163
transform 1 0 22816 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_240
timestamp 1667941163
transform 1 0 23184 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1667941163
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_264
timestamp 1667941163
transform 1 0 25392 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_284
timestamp 1667941163
transform 1 0 27232 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_300
timestamp 1667941163
transform 1 0 28704 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_323
timestamp 1667941163
transform 1 0 30820 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_333
timestamp 1667941163
transform 1 0 31740 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_337
timestamp 1667941163
transform 1 0 32108 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_344
timestamp 1667941163
transform 1 0 32752 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_360
timestamp 1667941163
transform 1 0 34224 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1667941163
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1667941163
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1667941163
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1667941163
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_421
timestamp 1667941163
transform 1 0 39836 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_435
timestamp 1667941163
transform 1 0 41124 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_443
timestamp 1667941163
transform 1 0 41860 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_449
timestamp 1667941163
transform 1 0 42412 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_455
timestamp 1667941163
transform 1 0 42964 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_461
timestamp 1667941163
transform 1 0 43516 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_470
timestamp 1667941163
transform 1 0 44344 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_42_477
timestamp 1667941163
transform 1 0 44988 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_484
timestamp 1667941163
transform 1 0 45632 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_492
timestamp 1667941163
transform 1 0 46368 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_514
timestamp 1667941163
transform 1 0 48392 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_14
timestamp 1667941163
transform 1 0 2392 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_26
timestamp 1667941163
transform 1 0 3496 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_38
timestamp 1667941163
transform 1 0 4600 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_50
timestamp 1667941163
transform 1 0 5704 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_75
timestamp 1667941163
transform 1 0 8004 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_87
timestamp 1667941163
transform 1 0 9108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_99
timestamp 1667941163
transform 1 0 10212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1667941163
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_131
timestamp 1667941163
transform 1 0 13156 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_143
timestamp 1667941163
transform 1 0 14260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_155
timestamp 1667941163
transform 1 0 15364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1667941163
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_184
timestamp 1667941163
transform 1 0 18032 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_192
timestamp 1667941163
transform 1 0 18768 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_202
timestamp 1667941163
transform 1 0 19688 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1667941163
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_230
timestamp 1667941163
transform 1 0 22264 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_236
timestamp 1667941163
transform 1 0 22816 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_253
timestamp 1667941163
transform 1 0 24380 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_261
timestamp 1667941163
transform 1 0 25116 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_269
timestamp 1667941163
transform 1 0 25852 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_276
timestamp 1667941163
transform 1 0 26496 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_305
timestamp 1667941163
transform 1 0 29164 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_325
timestamp 1667941163
transform 1 0 31004 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_333
timestamp 1667941163
transform 1 0 31740 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_348
timestamp 1667941163
transform 1 0 33120 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_43_367
timestamp 1667941163
transform 1 0 34868 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_382
timestamp 1667941163
transform 1 0 36248 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_390
timestamp 1667941163
transform 1 0 36984 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_399
timestamp 1667941163
transform 1 0 37812 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_406
timestamp 1667941163
transform 1 0 38456 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_417
timestamp 1667941163
transform 1 0 39468 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_427
timestamp 1667941163
transform 1 0 40388 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_439
timestamp 1667941163
transform 1 0 41492 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1667941163
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1667941163
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_461
timestamp 1667941163
transform 1 0 43516 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_473
timestamp 1667941163
transform 1 0 44620 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_502
timestamp 1667941163
transform 1 0 47288 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_505
timestamp 1667941163
transform 1 0 47564 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_510
timestamp 1667941163
transform 1 0 48024 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1667941163
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1667941163
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1667941163
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1667941163
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1667941163
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1667941163
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_89
timestamp 1667941163
transform 1 0 9292 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1667941163
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_109
timestamp 1667941163
transform 1 0 11132 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_117
timestamp 1667941163
transform 1 0 11868 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_122
timestamp 1667941163
transform 1 0 12328 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_134
timestamp 1667941163
transform 1 0 13432 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_145
timestamp 1667941163
transform 1 0 14444 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_154
timestamp 1667941163
transform 1 0 15272 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_166
timestamp 1667941163
transform 1 0 16376 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_180
timestamp 1667941163
transform 1 0 17664 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_187
timestamp 1667941163
transform 1 0 18308 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1667941163
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_206
timestamp 1667941163
transform 1 0 20056 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_219
timestamp 1667941163
transform 1 0 21252 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_231
timestamp 1667941163
transform 1 0 22356 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_239
timestamp 1667941163
transform 1 0 23092 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1667941163
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_263
timestamp 1667941163
transform 1 0 25300 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_275
timestamp 1667941163
transform 1 0 26404 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_287
timestamp 1667941163
transform 1 0 27508 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_299
timestamp 1667941163
transform 1 0 28612 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1667941163
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_333
timestamp 1667941163
transform 1 0 31740 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_352
timestamp 1667941163
transform 1 0 33488 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_383
timestamp 1667941163
transform 1 0 36340 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_394
timestamp 1667941163
transform 1 0 37352 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_404
timestamp 1667941163
transform 1 0 38272 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_410
timestamp 1667941163
transform 1 0 38824 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_418
timestamp 1667941163
transform 1 0 39560 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_421
timestamp 1667941163
transform 1 0 39836 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_439
timestamp 1667941163
transform 1 0 41492 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_451
timestamp 1667941163
transform 1 0 42596 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_463
timestamp 1667941163
transform 1 0 43700 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1667941163
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1667941163
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1667941163
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_489
timestamp 1667941163
transform 1 0 46092 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_514
timestamp 1667941163
transform 1 0 48392 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1667941163
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1667941163
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1667941163
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1667941163
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_70
timestamp 1667941163
transform 1 0 7544 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_74
timestamp 1667941163
transform 1 0 7912 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_79
timestamp 1667941163
transform 1 0 8372 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_99
timestamp 1667941163
transform 1 0 10212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1667941163
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1667941163
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_137
timestamp 1667941163
transform 1 0 13708 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_157
timestamp 1667941163
transform 1 0 15548 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_165
timestamp 1667941163
transform 1 0 16284 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_178
timestamp 1667941163
transform 1 0 17480 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_187
timestamp 1667941163
transform 1 0 18308 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_199
timestamp 1667941163
transform 1 0 19412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_211
timestamp 1667941163
transform 1 0 20516 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1667941163
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1667941163
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1667941163
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_261
timestamp 1667941163
transform 1 0 25116 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_271
timestamp 1667941163
transform 1 0 26036 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1667941163
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_291
timestamp 1667941163
transform 1 0 27876 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_303
timestamp 1667941163
transform 1 0 28980 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_315
timestamp 1667941163
transform 1 0 30084 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_327
timestamp 1667941163
transform 1 0 31188 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1667941163
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_355
timestamp 1667941163
transform 1 0 33764 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_367
timestamp 1667941163
transform 1 0 34868 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_373
timestamp 1667941163
transform 1 0 35420 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_386
timestamp 1667941163
transform 1 0 36616 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_398
timestamp 1667941163
transform 1 0 37720 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_410
timestamp 1667941163
transform 1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_420
timestamp 1667941163
transform 1 0 39744 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_429
timestamp 1667941163
transform 1 0 40572 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_446
timestamp 1667941163
transform 1 0 42136 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1667941163
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_461
timestamp 1667941163
transform 1 0 43516 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_481
timestamp 1667941163
transform 1 0 45356 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_493
timestamp 1667941163
transform 1 0 46460 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_498
timestamp 1667941163
transform 1 0 46920 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_505
timestamp 1667941163
transform 1 0 47564 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_510
timestamp 1667941163
transform 1 0 48024 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1667941163
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1667941163
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_47
timestamp 1667941163
transform 1 0 5428 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_67
timestamp 1667941163
transform 1 0 7268 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_78
timestamp 1667941163
transform 1 0 8280 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_104
timestamp 1667941163
transform 1 0 10672 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_116
timestamp 1667941163
transform 1 0 11776 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_129
timestamp 1667941163
transform 1 0 12972 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_137
timestamp 1667941163
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_149
timestamp 1667941163
transform 1 0 14812 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_161
timestamp 1667941163
transform 1 0 15916 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_173
timestamp 1667941163
transform 1 0 17020 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_184
timestamp 1667941163
transform 1 0 18032 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1667941163
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1667941163
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_233
timestamp 1667941163
transform 1 0 22540 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_242
timestamp 1667941163
transform 1 0 23368 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_250
timestamp 1667941163
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_257
timestamp 1667941163
transform 1 0 24748 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_274
timestamp 1667941163
transform 1 0 26312 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_278
timestamp 1667941163
transform 1 0 26680 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_295
timestamp 1667941163
transform 1 0 28244 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1667941163
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_319
timestamp 1667941163
transform 1 0 30452 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_331
timestamp 1667941163
transform 1 0 31556 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_349
timestamp 1667941163
transform 1 0 33212 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_361
timestamp 1667941163
transform 1 0 34316 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_386
timestamp 1667941163
transform 1 0 36616 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_398
timestamp 1667941163
transform 1 0 37720 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_408
timestamp 1667941163
transform 1 0 38640 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_421
timestamp 1667941163
transform 1 0 39836 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_427
timestamp 1667941163
transform 1 0 40388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_458
timestamp 1667941163
transform 1 0 43240 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_464
timestamp 1667941163
transform 1 0 43792 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_472
timestamp 1667941163
transform 1 0 44528 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1667941163
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_489
timestamp 1667941163
transform 1 0 46092 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_514
timestamp 1667941163
transform 1 0 48392 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1667941163
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1667941163
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1667941163
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1667941163
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1667941163
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_66
timestamp 1667941163
transform 1 0 7176 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_78
timestamp 1667941163
transform 1 0 8280 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_84
timestamp 1667941163
transform 1 0 8832 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_88
timestamp 1667941163
transform 1 0 9200 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_100
timestamp 1667941163
transform 1 0 10304 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_109
timestamp 1667941163
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_132
timestamp 1667941163
transform 1 0 13248 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_144
timestamp 1667941163
transform 1 0 14352 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_156
timestamp 1667941163
transform 1 0 15456 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_187
timestamp 1667941163
transform 1 0 18308 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_199
timestamp 1667941163
transform 1 0 19412 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_205
timestamp 1667941163
transform 1 0 19964 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_212
timestamp 1667941163
transform 1 0 20608 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_243
timestamp 1667941163
transform 1 0 23460 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_255
timestamp 1667941163
transform 1 0 24564 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_261
timestamp 1667941163
transform 1 0 25116 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_268
timestamp 1667941163
transform 1 0 25760 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_289
timestamp 1667941163
transform 1 0 27692 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1667941163
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1667941163
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1667941163
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_369
timestamp 1667941163
transform 1 0 35052 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_381
timestamp 1667941163
transform 1 0 36156 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_389
timestamp 1667941163
transform 1 0 36892 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_401
timestamp 1667941163
transform 1 0 37996 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_407
timestamp 1667941163
transform 1 0 38548 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_419
timestamp 1667941163
transform 1 0 39652 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_433
timestamp 1667941163
transform 1 0 40940 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_47_445
timestamp 1667941163
transform 1 0 42044 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_449
timestamp 1667941163
transform 1 0 42412 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_461
timestamp 1667941163
transform 1 0 43516 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_468
timestamp 1667941163
transform 1 0 44160 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_472
timestamp 1667941163
transform 1 0 44528 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_490
timestamp 1667941163
transform 1 0 46184 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_502
timestamp 1667941163
transform 1 0 47288 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_505
timestamp 1667941163
transform 1 0 47564 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_510
timestamp 1667941163
transform 1 0 48024 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1667941163
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_66
timestamp 1667941163
transform 1 0 7176 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_74
timestamp 1667941163
transform 1 0 7912 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_79
timestamp 1667941163
transform 1 0 8372 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1667941163
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_96
timestamp 1667941163
transform 1 0 9936 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_108
timestamp 1667941163
transform 1 0 11040 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_122
timestamp 1667941163
transform 1 0 12328 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_129
timestamp 1667941163
transform 1 0 12972 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_138
timestamp 1667941163
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_152
timestamp 1667941163
transform 1 0 15088 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_164
timestamp 1667941163
transform 1 0 16192 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_170
timestamp 1667941163
transform 1 0 16744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_180
timestamp 1667941163
transform 1 0 17664 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_191
timestamp 1667941163
transform 1 0 18676 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1667941163
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_205
timestamp 1667941163
transform 1 0 19964 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_217
timestamp 1667941163
transform 1 0 21068 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_235
timestamp 1667941163
transform 1 0 22724 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1667941163
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_258
timestamp 1667941163
transform 1 0 24840 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_270
timestamp 1667941163
transform 1 0 25944 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_282
timestamp 1667941163
transform 1 0 27048 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_294
timestamp 1667941163
transform 1 0 28152 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_306
timestamp 1667941163
transform 1 0 29256 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_317
timestamp 1667941163
transform 1 0 30268 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_325
timestamp 1667941163
transform 1 0 31004 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_343
timestamp 1667941163
transform 1 0 32660 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_355
timestamp 1667941163
transform 1 0 33764 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1667941163
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_385
timestamp 1667941163
transform 1 0 36524 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_391
timestamp 1667941163
transform 1 0 37076 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_397
timestamp 1667941163
transform 1 0 37628 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_403
timestamp 1667941163
transform 1 0 38180 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_410
timestamp 1667941163
transform 1 0 38824 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_48_417
timestamp 1667941163
transform 1 0 39468 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_421
timestamp 1667941163
transform 1 0 39836 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_427
timestamp 1667941163
transform 1 0 40388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_439
timestamp 1667941163
transform 1 0 41492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_445
timestamp 1667941163
transform 1 0 42044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_453
timestamp 1667941163
transform 1 0 42780 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_461
timestamp 1667941163
transform 1 0 43516 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_468
timestamp 1667941163
transform 1 0 44160 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1667941163
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_489
timestamp 1667941163
transform 1 0 46092 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_514
timestamp 1667941163
transform 1 0 48392 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1667941163
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1667941163
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_39
timestamp 1667941163
transform 1 0 4692 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_49_50
timestamp 1667941163
transform 1 0 5704 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_64
timestamp 1667941163
transform 1 0 6992 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_92
timestamp 1667941163
transform 1 0 9568 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_104
timestamp 1667941163
transform 1 0 10672 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_125
timestamp 1667941163
transform 1 0 12604 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_49_149
timestamp 1667941163
transform 1 0 14812 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_155
timestamp 1667941163
transform 1 0 15364 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1667941163
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1667941163
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_181
timestamp 1667941163
transform 1 0 17756 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_199
timestamp 1667941163
transform 1 0 19412 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_219
timestamp 1667941163
transform 1 0 21252 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1667941163
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_235
timestamp 1667941163
transform 1 0 22724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_247
timestamp 1667941163
transform 1 0 23828 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_255
timestamp 1667941163
transform 1 0 24564 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_267
timestamp 1667941163
transform 1 0 25668 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1667941163
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_290
timestamp 1667941163
transform 1 0 27784 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_296
timestamp 1667941163
transform 1 0 28336 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_313
timestamp 1667941163
transform 1 0 29900 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_323
timestamp 1667941163
transform 1 0 30820 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1667941163
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_347
timestamp 1667941163
transform 1 0 33028 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_357
timestamp 1667941163
transform 1 0 33948 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_377
timestamp 1667941163
transform 1 0 35788 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_389
timestamp 1667941163
transform 1 0 36892 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_401
timestamp 1667941163
transform 1 0 37996 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_410
timestamp 1667941163
transform 1 0 38824 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_418
timestamp 1667941163
transform 1 0 39560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_425
timestamp 1667941163
transform 1 0 40204 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_432
timestamp 1667941163
transform 1 0 40848 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_444
timestamp 1667941163
transform 1 0 41952 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_449
timestamp 1667941163
transform 1 0 42412 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_457
timestamp 1667941163
transform 1 0 43148 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_464
timestamp 1667941163
transform 1 0 43792 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_476
timestamp 1667941163
transform 1 0 44896 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_488
timestamp 1667941163
transform 1 0 46000 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_495
timestamp 1667941163
transform 1 0 46644 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_502
timestamp 1667941163
transform 1 0 47288 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_505
timestamp 1667941163
transform 1 0 47564 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_510
timestamp 1667941163
transform 1 0 48024 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1667941163
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1667941163
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1667941163
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_53
timestamp 1667941163
transform 1 0 5980 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_82
timestamp 1667941163
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_97
timestamp 1667941163
transform 1 0 10028 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_101
timestamp 1667941163
transform 1 0 10396 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1667941163
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_121
timestamp 1667941163
transform 1 0 12236 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_131
timestamp 1667941163
transform 1 0 13156 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1667941163
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_146
timestamp 1667941163
transform 1 0 14536 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_150
timestamp 1667941163
transform 1 0 14904 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_167
timestamp 1667941163
transform 1 0 16468 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_175
timestamp 1667941163
transform 1 0 17204 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_187
timestamp 1667941163
transform 1 0 18308 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1667941163
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_207
timestamp 1667941163
transform 1 0 20148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_235
timestamp 1667941163
transform 1 0 22724 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_244
timestamp 1667941163
transform 1 0 23552 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_266
timestamp 1667941163
transform 1 0 25576 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_286
timestamp 1667941163
transform 1 0 27416 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_298
timestamp 1667941163
transform 1 0 28520 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_306
timestamp 1667941163
transform 1 0 29256 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_319
timestamp 1667941163
transform 1 0 30452 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_327
timestamp 1667941163
transform 1 0 31188 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_346
timestamp 1667941163
transform 1 0 32936 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_354
timestamp 1667941163
transform 1 0 33672 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_362
timestamp 1667941163
transform 1 0 34408 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_378
timestamp 1667941163
transform 1 0 35880 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_390
timestamp 1667941163
transform 1 0 36984 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_394
timestamp 1667941163
transform 1 0 37352 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_404
timestamp 1667941163
transform 1 0 38272 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_414
timestamp 1667941163
transform 1 0 39192 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_421
timestamp 1667941163
transform 1 0 39836 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_439
timestamp 1667941163
transform 1 0 41492 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_451
timestamp 1667941163
transform 1 0 42596 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_459
timestamp 1667941163
transform 1 0 43332 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_468
timestamp 1667941163
transform 1 0 44160 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1667941163
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_489
timestamp 1667941163
transform 1 0 46092 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_514
timestamp 1667941163
transform 1 0 48392 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1667941163
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1667941163
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1667941163
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1667941163
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1667941163
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_66
timestamp 1667941163
transform 1 0 7176 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_78
timestamp 1667941163
transform 1 0 8280 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_106
timestamp 1667941163
transform 1 0 10856 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_124
timestamp 1667941163
transform 1 0 12512 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_131
timestamp 1667941163
transform 1 0 13156 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_143
timestamp 1667941163
transform 1 0 14260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_158
timestamp 1667941163
transform 1 0 15640 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1667941163
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_177
timestamp 1667941163
transform 1 0 17388 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_191
timestamp 1667941163
transform 1 0 18676 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_203
timestamp 1667941163
transform 1 0 19780 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_215
timestamp 1667941163
transform 1 0 20884 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1667941163
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_233
timestamp 1667941163
transform 1 0 22540 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_237
timestamp 1667941163
transform 1 0 22908 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_254
timestamp 1667941163
transform 1 0 24472 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_269
timestamp 1667941163
transform 1 0 25852 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_277
timestamp 1667941163
transform 1 0 26588 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_288
timestamp 1667941163
transform 1 0 27600 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_300
timestamp 1667941163
transform 1 0 28704 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_306
timestamp 1667941163
transform 1 0 29256 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_314
timestamp 1667941163
transform 1 0 29992 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_326
timestamp 1667941163
transform 1 0 31096 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_334
timestamp 1667941163
transform 1 0 31832 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_345
timestamp 1667941163
transform 1 0 32844 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_357
timestamp 1667941163
transform 1 0 33948 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_367
timestamp 1667941163
transform 1 0 34868 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_379
timestamp 1667941163
transform 1 0 35972 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1667941163
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_411
timestamp 1667941163
transform 1 0 38916 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_419
timestamp 1667941163
transform 1 0 39652 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_427
timestamp 1667941163
transform 1 0 40388 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_434
timestamp 1667941163
transform 1 0 41032 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_446
timestamp 1667941163
transform 1 0 42136 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_449
timestamp 1667941163
transform 1 0 42412 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_457
timestamp 1667941163
transform 1 0 43148 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_464
timestamp 1667941163
transform 1 0 43792 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1667941163
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1667941163
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_497
timestamp 1667941163
transform 1 0 46828 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_502
timestamp 1667941163
transform 1 0 47288 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_505
timestamp 1667941163
transform 1 0 47564 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_510
timestamp 1667941163
transform 1 0 48024 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1667941163
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1667941163
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1667941163
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_53
timestamp 1667941163
transform 1 0 5980 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1667941163
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_77
timestamp 1667941163
transform 1 0 8188 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 1667941163
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_91
timestamp 1667941163
transform 1 0 9476 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_96
timestamp 1667941163
transform 1 0 9936 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_118
timestamp 1667941163
transform 1 0 11960 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1667941163
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_153
timestamp 1667941163
transform 1 0 15180 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_157
timestamp 1667941163
transform 1 0 15548 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_161
timestamp 1667941163
transform 1 0 15916 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_167
timestamp 1667941163
transform 1 0 16468 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_184
timestamp 1667941163
transform 1 0 18032 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1667941163
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1667941163
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1667941163
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1667941163
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1667941163
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_261
timestamp 1667941163
transform 1 0 25116 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_272
timestamp 1667941163
transform 1 0 26128 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_284
timestamp 1667941163
transform 1 0 27232 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_296
timestamp 1667941163
transform 1 0 28336 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_52_305
timestamp 1667941163
transform 1 0 29164 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_320
timestamp 1667941163
transform 1 0 30544 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_332
timestamp 1667941163
transform 1 0 31648 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_344
timestamp 1667941163
transform 1 0 32752 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_356
timestamp 1667941163
transform 1 0 33856 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_385
timestamp 1667941163
transform 1 0 36524 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_398
timestamp 1667941163
transform 1 0 37720 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_410
timestamp 1667941163
transform 1 0 38824 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_418
timestamp 1667941163
transform 1 0 39560 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1667941163
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1667941163
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_445
timestamp 1667941163
transform 1 0 42044 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_452
timestamp 1667941163
transform 1 0 42688 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_465
timestamp 1667941163
transform 1 0 43884 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_474
timestamp 1667941163
transform 1 0 44712 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_477
timestamp 1667941163
transform 1 0 44988 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_495
timestamp 1667941163
transform 1 0 46644 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_507
timestamp 1667941163
transform 1 0 47748 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_515
timestamp 1667941163
transform 1 0 48484 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1667941163
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1667941163
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_54
timestamp 1667941163
transform 1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_80
timestamp 1667941163
transform 1 0 8464 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_90
timestamp 1667941163
transform 1 0 9384 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_98
timestamp 1667941163
transform 1 0 10120 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_103
timestamp 1667941163
transform 1 0 10580 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1667941163
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_121
timestamp 1667941163
transform 1 0 12236 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_126
timestamp 1667941163
transform 1 0 12696 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_139
timestamp 1667941163
transform 1 0 13892 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_151
timestamp 1667941163
transform 1 0 14996 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_155
timestamp 1667941163
transform 1 0 15364 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_162
timestamp 1667941163
transform 1 0 16008 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_178
timestamp 1667941163
transform 1 0 17480 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_185
timestamp 1667941163
transform 1 0 18124 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_197
timestamp 1667941163
transform 1 0 19228 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_208
timestamp 1667941163
transform 1 0 20240 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_220
timestamp 1667941163
transform 1 0 21344 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_249
timestamp 1667941163
transform 1 0 24012 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_255
timestamp 1667941163
transform 1 0 24564 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_263
timestamp 1667941163
transform 1 0 25300 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_270
timestamp 1667941163
transform 1 0 25944 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_278
timestamp 1667941163
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_312
timestamp 1667941163
transform 1 0 29808 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_319
timestamp 1667941163
transform 1 0 30452 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_327
timestamp 1667941163
transform 1 0 31188 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_331
timestamp 1667941163
transform 1 0 31556 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1667941163
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_353
timestamp 1667941163
transform 1 0 33580 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_370
timestamp 1667941163
transform 1 0 35144 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_380
timestamp 1667941163
transform 1 0 36064 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_402
timestamp 1667941163
transform 1 0 38088 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_410
timestamp 1667941163
transform 1 0 38824 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_415
timestamp 1667941163
transform 1 0 39284 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_427
timestamp 1667941163
transform 1 0 40388 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_439
timestamp 1667941163
transform 1 0 41492 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1667941163
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_449
timestamp 1667941163
transform 1 0 42412 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_453
timestamp 1667941163
transform 1 0 42780 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_470
timestamp 1667941163
transform 1 0 44344 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_477
timestamp 1667941163
transform 1 0 44988 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_489
timestamp 1667941163
transform 1 0 46092 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_501
timestamp 1667941163
transform 1 0 47196 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1667941163
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_513
timestamp 1667941163
transform 1 0 48300 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1667941163
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_35
timestamp 1667941163
transform 1 0 4324 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_39
timestamp 1667941163
transform 1 0 4692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_57
timestamp 1667941163
transform 1 0 6348 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_68
timestamp 1667941163
transform 1 0 7360 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_80
timestamp 1667941163
transform 1 0 8464 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_91
timestamp 1667941163
transform 1 0 9476 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_99
timestamp 1667941163
transform 1 0 10212 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1667941163
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1667941163
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1667941163
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1667941163
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_149
timestamp 1667941163
transform 1 0 14812 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_169
timestamp 1667941163
transform 1 0 16652 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_182
timestamp 1667941163
transform 1 0 17848 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_194
timestamp 1667941163
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_215
timestamp 1667941163
transform 1 0 20884 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_223
timestamp 1667941163
transform 1 0 21620 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_234
timestamp 1667941163
transform 1 0 22632 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_242
timestamp 1667941163
transform 1 0 23368 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_250
timestamp 1667941163
transform 1 0 24104 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_261
timestamp 1667941163
transform 1 0 25116 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_271
timestamp 1667941163
transform 1 0 26036 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_283
timestamp 1667941163
transform 1 0 27140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_295
timestamp 1667941163
transform 1 0 28244 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1667941163
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_327
timestamp 1667941163
transform 1 0 31188 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_338
timestamp 1667941163
transform 1 0 32200 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_350
timestamp 1667941163
transform 1 0 33304 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_362
timestamp 1667941163
transform 1 0 34408 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_371
timestamp 1667941163
transform 1 0 35236 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_388
timestamp 1667941163
transform 1 0 36800 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_54_405
timestamp 1667941163
transform 1 0 38364 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_416
timestamp 1667941163
transform 1 0 39376 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_421
timestamp 1667941163
transform 1 0 39836 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_439
timestamp 1667941163
transform 1 0 41492 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_451
timestamp 1667941163
transform 1 0 42596 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_463
timestamp 1667941163
transform 1 0 43700 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1667941163
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_477
timestamp 1667941163
transform 1 0 44988 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_485
timestamp 1667941163
transform 1 0 45724 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_507
timestamp 1667941163
transform 1 0 47748 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_515
timestamp 1667941163
transform 1 0 48484 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_8
timestamp 1667941163
transform 1 0 1840 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_20
timestamp 1667941163
transform 1 0 2944 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_28
timestamp 1667941163
transform 1 0 3680 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_50
timestamp 1667941163
transform 1 0 5704 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_63
timestamp 1667941163
transform 1 0 6900 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_75
timestamp 1667941163
transform 1 0 8004 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_83
timestamp 1667941163
transform 1 0 8740 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_101
timestamp 1667941163
transform 1 0 10396 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_108
timestamp 1667941163
transform 1 0 11040 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_122
timestamp 1667941163
transform 1 0 12328 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_130
timestamp 1667941163
transform 1 0 13064 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_147
timestamp 1667941163
transform 1 0 14628 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_160
timestamp 1667941163
transform 1 0 15824 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_186
timestamp 1667941163
transform 1 0 18216 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_199
timestamp 1667941163
transform 1 0 19412 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_207
timestamp 1667941163
transform 1 0 20148 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_214
timestamp 1667941163
transform 1 0 20792 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_222
timestamp 1667941163
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_243
timestamp 1667941163
transform 1 0 23460 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_264
timestamp 1667941163
transform 1 0 25392 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_278
timestamp 1667941163
transform 1 0 26680 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_300
timestamp 1667941163
transform 1 0 28704 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_312
timestamp 1667941163
transform 1 0 29808 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_324
timestamp 1667941163
transform 1 0 30912 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_332
timestamp 1667941163
transform 1 0 31648 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_362
timestamp 1667941163
transform 1 0 34408 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_377
timestamp 1667941163
transform 1 0 35788 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_386
timestamp 1667941163
transform 1 0 36616 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_417
timestamp 1667941163
transform 1 0 39468 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1667941163
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1667941163
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1667941163
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1667941163
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1667941163
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_473
timestamp 1667941163
transform 1 0 44620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_477
timestamp 1667941163
transform 1 0 44988 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_502
timestamp 1667941163
transform 1 0 47288 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_505
timestamp 1667941163
transform 1 0 47564 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_510
timestamp 1667941163
transform 1 0 48024 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1667941163
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1667941163
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_34
timestamp 1667941163
transform 1 0 4232 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_42
timestamp 1667941163
transform 1 0 4968 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_49
timestamp 1667941163
transform 1 0 5612 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_69
timestamp 1667941163
transform 1 0 7452 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_79
timestamp 1667941163
transform 1 0 8372 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1667941163
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_93
timestamp 1667941163
transform 1 0 9660 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_103
timestamp 1667941163
transform 1 0 10580 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_115
timestamp 1667941163
transform 1 0 11684 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_119
timestamp 1667941163
transform 1 0 12052 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_129
timestamp 1667941163
transform 1 0 12972 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_138
timestamp 1667941163
transform 1 0 13800 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1667941163
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1667941163
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_177
timestamp 1667941163
transform 1 0 17388 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1667941163
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1667941163
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_205
timestamp 1667941163
transform 1 0 19964 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_218
timestamp 1667941163
transform 1 0 21160 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_227
timestamp 1667941163
transform 1 0 21988 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_235
timestamp 1667941163
transform 1 0 22724 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_243
timestamp 1667941163
transform 1 0 23460 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1667941163
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_56_275
timestamp 1667941163
transform 1 0 26404 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_283
timestamp 1667941163
transform 1 0 27140 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_288
timestamp 1667941163
transform 1 0 27600 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_300
timestamp 1667941163
transform 1 0 28704 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_327
timestamp 1667941163
transform 1 0 31188 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_336
timestamp 1667941163
transform 1 0 32016 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_344
timestamp 1667941163
transform 1 0 32752 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_356
timestamp 1667941163
transform 1 0 33856 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_371
timestamp 1667941163
transform 1 0 35236 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_375
timestamp 1667941163
transform 1 0 35604 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_387
timestamp 1667941163
transform 1 0 36708 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_399
timestamp 1667941163
transform 1 0 37812 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_414
timestamp 1667941163
transform 1 0 39192 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_421
timestamp 1667941163
transform 1 0 39836 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_429
timestamp 1667941163
transform 1 0 40572 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_441
timestamp 1667941163
transform 1 0 41676 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_453
timestamp 1667941163
transform 1 0 42780 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_465
timestamp 1667941163
transform 1 0 43884 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_473
timestamp 1667941163
transform 1 0 44620 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_56_477
timestamp 1667941163
transform 1 0 44988 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_56_486
timestamp 1667941163
transform 1 0 45816 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_492
timestamp 1667941163
transform 1 0 46368 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_514
timestamp 1667941163
transform 1 0 48392 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1667941163
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_27
timestamp 1667941163
transform 1 0 3588 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_33
timestamp 1667941163
transform 1 0 4140 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_38
timestamp 1667941163
transform 1 0 4600 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_48
timestamp 1667941163
transform 1 0 5520 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_64
timestamp 1667941163
transform 1 0 6992 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_84
timestamp 1667941163
transform 1 0 8832 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_94
timestamp 1667941163
transform 1 0 9752 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_101
timestamp 1667941163
transform 1 0 10396 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_109
timestamp 1667941163
transform 1 0 11132 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_131
timestamp 1667941163
transform 1 0 13156 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_143
timestamp 1667941163
transform 1 0 14260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_155
timestamp 1667941163
transform 1 0 15364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1667941163
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_173
timestamp 1667941163
transform 1 0 17020 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_177
timestamp 1667941163
transform 1 0 17388 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_186
timestamp 1667941163
transform 1 0 18216 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_190
timestamp 1667941163
transform 1 0 18584 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_194
timestamp 1667941163
transform 1 0 18952 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_198
timestamp 1667941163
transform 1 0 19320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_203
timestamp 1667941163
transform 1 0 19780 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_210
timestamp 1667941163
transform 1 0 20424 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_216
timestamp 1667941163
transform 1 0 20976 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_220
timestamp 1667941163
transform 1 0 21344 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_245
timestamp 1667941163
transform 1 0 23644 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_257
timestamp 1667941163
transform 1 0 24748 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_271
timestamp 1667941163
transform 1 0 26036 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_278
timestamp 1667941163
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_288
timestamp 1667941163
transform 1 0 27600 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_295
timestamp 1667941163
transform 1 0 28244 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_307
timestamp 1667941163
transform 1 0 29348 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_321
timestamp 1667941163
transform 1 0 30636 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_333
timestamp 1667941163
transform 1 0 31740 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_343
timestamp 1667941163
transform 1 0 32660 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_347
timestamp 1667941163
transform 1 0 33028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_359
timestamp 1667941163
transform 1 0 34132 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_367
timestamp 1667941163
transform 1 0 34868 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_375
timestamp 1667941163
transform 1 0 35604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_387
timestamp 1667941163
transform 1 0 36708 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1667941163
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1667941163
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1667941163
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1667941163
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1667941163
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1667941163
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1667941163
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1667941163
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1667941163
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_497
timestamp 1667941163
transform 1 0 46828 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_501
timestamp 1667941163
transform 1 0 47196 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_505
timestamp 1667941163
transform 1 0 47564 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_513
timestamp 1667941163
transform 1 0 48300 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1667941163
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_49
timestamp 1667941163
transform 1 0 5612 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_61
timestamp 1667941163
transform 1 0 6716 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_68
timestamp 1667941163
transform 1 0 7360 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_76
timestamp 1667941163
transform 1 0 8096 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_89
timestamp 1667941163
transform 1 0 9292 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_106
timestamp 1667941163
transform 1 0 10856 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_118
timestamp 1667941163
transform 1 0 11960 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_122
timestamp 1667941163
transform 1 0 12328 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_130
timestamp 1667941163
transform 1 0 13064 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_136
timestamp 1667941163
transform 1 0 13616 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_146
timestamp 1667941163
transform 1 0 14536 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_154
timestamp 1667941163
transform 1 0 15272 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_171
timestamp 1667941163
transform 1 0 16836 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_183
timestamp 1667941163
transform 1 0 17940 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_58_193
timestamp 1667941163
transform 1 0 18860 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_208
timestamp 1667941163
transform 1 0 20240 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_219
timestamp 1667941163
transform 1 0 21252 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_231
timestamp 1667941163
transform 1 0 22356 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_243
timestamp 1667941163
transform 1 0 23460 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_274
timestamp 1667941163
transform 1 0 26312 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_282
timestamp 1667941163
transform 1 0 27048 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1667941163
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1667941163
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1667941163
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_319
timestamp 1667941163
transform 1 0 30452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_331
timestamp 1667941163
transform 1 0 31556 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_339
timestamp 1667941163
transform 1 0 32292 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_356
timestamp 1667941163
transform 1 0 33856 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_369
timestamp 1667941163
transform 1 0 35052 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_378
timestamp 1667941163
transform 1 0 35880 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_386
timestamp 1667941163
transform 1 0 36616 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_394
timestamp 1667941163
transform 1 0 37352 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_405
timestamp 1667941163
transform 1 0 38364 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_415
timestamp 1667941163
transform 1 0 39284 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1667941163
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1667941163
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1667941163
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1667941163
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1667941163
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1667941163
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1667941163
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1667941163
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1667941163
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1667941163
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_513
timestamp 1667941163
transform 1 0 48300 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_9
timestamp 1667941163
transform 1 0 1932 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_21
timestamp 1667941163
transform 1 0 3036 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_33
timestamp 1667941163
transform 1 0 4140 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_39
timestamp 1667941163
transform 1 0 4692 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_46
timestamp 1667941163
transform 1 0 5336 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_53
timestamp 1667941163
transform 1 0 5980 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_81
timestamp 1667941163
transform 1 0 8556 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_87
timestamp 1667941163
transform 1 0 9108 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_95
timestamp 1667941163
transform 1 0 9844 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_107
timestamp 1667941163
transform 1 0 10948 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1667941163
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_144
timestamp 1667941163
transform 1 0 14352 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_154
timestamp 1667941163
transform 1 0 15272 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_166
timestamp 1667941163
transform 1 0 16376 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_179
timestamp 1667941163
transform 1 0 17572 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_187
timestamp 1667941163
transform 1 0 18308 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_192
timestamp 1667941163
transform 1 0 18768 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_204
timestamp 1667941163
transform 1 0 19872 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_212
timestamp 1667941163
transform 1 0 20608 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1667941163
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1667941163
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_234
timestamp 1667941163
transform 1 0 22632 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_242
timestamp 1667941163
transform 1 0 23368 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_253
timestamp 1667941163
transform 1 0 24380 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_260
timestamp 1667941163
transform 1 0 25024 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_272
timestamp 1667941163
transform 1 0 26128 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_288
timestamp 1667941163
transform 1 0 27600 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_300
timestamp 1667941163
transform 1 0 28704 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_306
timestamp 1667941163
transform 1 0 29256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_313
timestamp 1667941163
transform 1 0 29900 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_325
timestamp 1667941163
transform 1 0 31004 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_333
timestamp 1667941163
transform 1 0 31740 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_353
timestamp 1667941163
transform 1 0 33580 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_357
timestamp 1667941163
transform 1 0 33948 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_366
timestamp 1667941163
transform 1 0 34776 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_374
timestamp 1667941163
transform 1 0 35512 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_380
timestamp 1667941163
transform 1 0 36064 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_390
timestamp 1667941163
transform 1 0 36984 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_398
timestamp 1667941163
transform 1 0 37720 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_420
timestamp 1667941163
transform 1 0 39744 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_432
timestamp 1667941163
transform 1 0 40848 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_444
timestamp 1667941163
transform 1 0 41952 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1667941163
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1667941163
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1667941163
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1667941163
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1667941163
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1667941163
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_505
timestamp 1667941163
transform 1 0 47564 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_513
timestamp 1667941163
transform 1 0 48300 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1667941163
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_51
timestamp 1667941163
transform 1 0 5796 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_63
timestamp 1667941163
transform 1 0 6900 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_71
timestamp 1667941163
transform 1 0 7636 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_81
timestamp 1667941163
transform 1 0 8556 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1667941163
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1667941163
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1667941163
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_153
timestamp 1667941163
transform 1 0 15180 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_157
timestamp 1667941163
transform 1 0 15548 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_174
timestamp 1667941163
transform 1 0 17112 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_185
timestamp 1667941163
transform 1 0 18124 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_193
timestamp 1667941163
transform 1 0 18860 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_217
timestamp 1667941163
transform 1 0 21068 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_227
timestamp 1667941163
transform 1 0 21988 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_60_249
timestamp 1667941163
transform 1 0 24012 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_264
timestamp 1667941163
transform 1 0 25392 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_274
timestamp 1667941163
transform 1 0 26312 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_282
timestamp 1667941163
transform 1 0 27048 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_292
timestamp 1667941163
transform 1 0 27968 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_303
timestamp 1667941163
transform 1 0 28980 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1667941163
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_60_328
timestamp 1667941163
transform 1 0 31280 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_334
timestamp 1667941163
transform 1 0 31832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_343
timestamp 1667941163
transform 1 0 32660 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_353
timestamp 1667941163
transform 1 0 33580 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_361
timestamp 1667941163
transform 1 0 34316 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_384
timestamp 1667941163
transform 1 0 36432 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_388
timestamp 1667941163
transform 1 0 36800 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_405
timestamp 1667941163
transform 1 0 38364 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_417
timestamp 1667941163
transform 1 0 39468 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1667941163
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1667941163
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1667941163
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1667941163
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1667941163
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1667941163
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1667941163
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1667941163
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1667941163
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_513
timestamp 1667941163
transform 1 0 48300 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1667941163
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1667941163
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_39
timestamp 1667941163
transform 1 0 4692 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_43
timestamp 1667941163
transform 1 0 5060 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_50
timestamp 1667941163
transform 1 0 5704 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1667941163
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_137
timestamp 1667941163
transform 1 0 13708 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_147
timestamp 1667941163
transform 1 0 14628 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_159
timestamp 1667941163
transform 1 0 15732 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1667941163
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_188
timestamp 1667941163
transform 1 0 18400 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_200
timestamp 1667941163
transform 1 0 19504 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_212
timestamp 1667941163
transform 1 0 20608 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_218
timestamp 1667941163
transform 1 0 21160 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_222
timestamp 1667941163
transform 1 0 21528 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_231
timestamp 1667941163
transform 1 0 22356 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_61_246
timestamp 1667941163
transform 1 0 23736 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_254
timestamp 1667941163
transform 1 0 24472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_261
timestamp 1667941163
transform 1 0 25116 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_269
timestamp 1667941163
transform 1 0 25852 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_276
timestamp 1667941163
transform 1 0 26496 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_287
timestamp 1667941163
transform 1 0 27508 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_299
timestamp 1667941163
transform 1 0 28612 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_311
timestamp 1667941163
transform 1 0 29716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_323
timestamp 1667941163
transform 1 0 30820 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1667941163
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_355
timestamp 1667941163
transform 1 0 33764 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_367
timestamp 1667941163
transform 1 0 34868 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_374
timestamp 1667941163
transform 1 0 35512 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_386
timestamp 1667941163
transform 1 0 36616 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1667941163
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1667941163
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1667941163
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1667941163
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1667941163
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1667941163
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1667941163
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1667941163
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1667941163
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1667941163
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_505
timestamp 1667941163
transform 1 0 47564 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_510
timestamp 1667941163
transform 1 0 48024 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1667941163
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1667941163
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_33
timestamp 1667941163
transform 1 0 4140 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_38
timestamp 1667941163
transform 1 0 4600 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_42
timestamp 1667941163
transform 1 0 4968 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_49
timestamp 1667941163
transform 1 0 5612 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_56
timestamp 1667941163
transform 1 0 6256 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_68
timestamp 1667941163
transform 1 0 7360 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_80
timestamp 1667941163
transform 1 0 8464 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_93
timestamp 1667941163
transform 1 0 9660 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_100
timestamp 1667941163
transform 1 0 10304 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_112
timestamp 1667941163
transform 1 0 11408 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_124
timestamp 1667941163
transform 1 0 12512 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_136
timestamp 1667941163
transform 1 0 13616 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_165
timestamp 1667941163
transform 1 0 16284 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_171
timestamp 1667941163
transform 1 0 16836 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_178
timestamp 1667941163
transform 1 0 17480 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_190
timestamp 1667941163
transform 1 0 18584 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_217
timestamp 1667941163
transform 1 0 21068 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_225
timestamp 1667941163
transform 1 0 21804 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_237
timestamp 1667941163
transform 1 0 22908 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_245
timestamp 1667941163
transform 1 0 23644 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_250
timestamp 1667941163
transform 1 0 24104 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_262
timestamp 1667941163
transform 1 0 25208 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_269
timestamp 1667941163
transform 1 0 25852 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_273
timestamp 1667941163
transform 1 0 26220 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_279
timestamp 1667941163
transform 1 0 26772 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_285
timestamp 1667941163
transform 1 0 27324 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_293
timestamp 1667941163
transform 1 0 28060 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_305
timestamp 1667941163
transform 1 0 29164 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1667941163
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1667941163
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1667941163
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1667941163
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1667941163
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1667941163
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1667941163
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1667941163
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1667941163
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1667941163
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1667941163
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1667941163
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_489
timestamp 1667941163
transform 1 0 46092 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_514
timestamp 1667941163
transform 1 0 48392 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1667941163
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_27
timestamp 1667941163
transform 1 0 3588 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_33
timestamp 1667941163
transform 1 0 4140 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_50
timestamp 1667941163
transform 1 0 5704 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_69
timestamp 1667941163
transform 1 0 7452 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_89
timestamp 1667941163
transform 1 0 9292 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_101
timestamp 1667941163
transform 1 0 10396 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_109
timestamp 1667941163
transform 1 0 11132 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_125
timestamp 1667941163
transform 1 0 12604 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_144
timestamp 1667941163
transform 1 0 14352 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_152
timestamp 1667941163
transform 1 0 15088 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_159
timestamp 1667941163
transform 1 0 15732 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1667941163
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1667941163
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_193
timestamp 1667941163
transform 1 0 18860 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_197
timestamp 1667941163
transform 1 0 19228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_205
timestamp 1667941163
transform 1 0 19964 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_216
timestamp 1667941163
transform 1 0 20976 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_233
timestamp 1667941163
transform 1 0 22540 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_245
timestamp 1667941163
transform 1 0 23644 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_253
timestamp 1667941163
transform 1 0 24380 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_260
timestamp 1667941163
transform 1 0 25024 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_267
timestamp 1667941163
transform 1 0 25668 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1667941163
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1667941163
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1667941163
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1667941163
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1667941163
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1667941163
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1667941163
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1667941163
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1667941163
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1667941163
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1667941163
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1667941163
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1667941163
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1667941163
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1667941163
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1667941163
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1667941163
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1667941163
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1667941163
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1667941163
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1667941163
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_505
timestamp 1667941163
transform 1 0 47564 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_510
timestamp 1667941163
transform 1 0 48024 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_11
timestamp 1667941163
transform 1 0 2116 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1667941163
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1667941163
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_36
timestamp 1667941163
transform 1 0 4416 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_56
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_66
timestamp 1667941163
transform 1 0 7176 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_70
timestamp 1667941163
transform 1 0 7544 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1667941163
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1667941163
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_90
timestamp 1667941163
transform 1 0 9384 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_102
timestamp 1667941163
transform 1 0 10488 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_114
timestamp 1667941163
transform 1 0 11592 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_129
timestamp 1667941163
transform 1 0 12972 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_138
timestamp 1667941163
transform 1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_151
timestamp 1667941163
transform 1 0 14996 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_162
timestamp 1667941163
transform 1 0 16008 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_174
timestamp 1667941163
transform 1 0 17112 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_192
timestamp 1667941163
transform 1 0 18768 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_208
timestamp 1667941163
transform 1 0 20240 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_228
timestamp 1667941163
transform 1 0 22080 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_240
timestamp 1667941163
transform 1 0 23184 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_265
timestamp 1667941163
transform 1 0 25484 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_287
timestamp 1667941163
transform 1 0 27508 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_299
timestamp 1667941163
transform 1 0 28612 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1667941163
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1667941163
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1667941163
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1667941163
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1667941163
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1667941163
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1667941163
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1667941163
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1667941163
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1667941163
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1667941163
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1667941163
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1667941163
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1667941163
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1667941163
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1667941163
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1667941163
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1667941163
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_489
timestamp 1667941163
transform 1 0 46092 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_514
timestamp 1667941163
transform 1 0 48392 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1667941163
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1667941163
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_27
timestamp 1667941163
transform 1 0 3588 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_35
timestamp 1667941163
transform 1 0 4324 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_42
timestamp 1667941163
transform 1 0 4968 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_50
timestamp 1667941163
transform 1 0 5704 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_54
timestamp 1667941163
transform 1 0 6072 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_57
timestamp 1667941163
transform 1 0 6348 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_75
timestamp 1667941163
transform 1 0 8004 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_83
timestamp 1667941163
transform 1 0 8740 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_95
timestamp 1667941163
transform 1 0 9844 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_107
timestamp 1667941163
transform 1 0 10948 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1667941163
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1667941163
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_125
timestamp 1667941163
transform 1 0 12604 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_131
timestamp 1667941163
transform 1 0 13156 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_135
timestamp 1667941163
transform 1 0 13524 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_145
timestamp 1667941163
transform 1 0 14444 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_154
timestamp 1667941163
transform 1 0 15272 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_166
timestamp 1667941163
transform 1 0 16376 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_169
timestamp 1667941163
transform 1 0 16652 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_177
timestamp 1667941163
transform 1 0 17388 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_181
timestamp 1667941163
transform 1 0 17756 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_192
timestamp 1667941163
transform 1 0 18768 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_198
timestamp 1667941163
transform 1 0 19320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_206
timestamp 1667941163
transform 1 0 20056 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_216
timestamp 1667941163
transform 1 0 20976 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1667941163
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_237
timestamp 1667941163
transform 1 0 22908 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_255
timestamp 1667941163
transform 1 0 24564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_267
timestamp 1667941163
transform 1 0 25668 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1667941163
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1667941163
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1667941163
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1667941163
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1667941163
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1667941163
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1667941163
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_337
timestamp 1667941163
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_349
timestamp 1667941163
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1667941163
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_373
timestamp 1667941163
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1667941163
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1667941163
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1667941163
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1667941163
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1667941163
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1667941163
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1667941163
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1667941163
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1667941163
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1667941163
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1667941163
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1667941163
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1667941163
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1667941163
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_505
timestamp 1667941163
transform 1 0 47564 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_510
timestamp 1667941163
transform 1 0 48024 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1667941163
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1667941163
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1667941163
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1667941163
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1667941163
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_53
timestamp 1667941163
transform 1 0 5980 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_57
timestamp 1667941163
transform 1 0 6348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_62
timestamp 1667941163
transform 1 0 6808 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_74
timestamp 1667941163
transform 1 0 7912 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_82
timestamp 1667941163
transform 1 0 8648 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1667941163
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1667941163
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_109
timestamp 1667941163
transform 1 0 11132 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_117
timestamp 1667941163
transform 1 0 11868 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_136
timestamp 1667941163
transform 1 0 13616 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_141
timestamp 1667941163
transform 1 0 14076 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_153
timestamp 1667941163
transform 1 0 15180 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_173
timestamp 1667941163
transform 1 0 17020 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_177
timestamp 1667941163
transform 1 0 17388 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_194
timestamp 1667941163
transform 1 0 18952 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1667941163
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1667941163
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_221
timestamp 1667941163
transform 1 0 21436 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_229
timestamp 1667941163
transform 1 0 22172 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_235
timestamp 1667941163
transform 1 0 22724 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1667941163
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1667941163
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_253
timestamp 1667941163
transform 1 0 24380 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_271
timestamp 1667941163
transform 1 0 26036 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_283
timestamp 1667941163
transform 1 0 27140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_295
timestamp 1667941163
transform 1 0 28244 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1667941163
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1667941163
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1667941163
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_333
timestamp 1667941163
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_345
timestamp 1667941163
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1667941163
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1667941163
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1667941163
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1667941163
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1667941163
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1667941163
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1667941163
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1667941163
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1667941163
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1667941163
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1667941163
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1667941163
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1667941163
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1667941163
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1667941163
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1667941163
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_501
timestamp 1667941163
transform 1 0 47196 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_507
timestamp 1667941163
transform 1 0 47748 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_515
timestamp 1667941163
transform 1 0 48484 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_3
timestamp 1667941163
transform 1 0 1380 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_11
timestamp 1667941163
transform 1 0 2116 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_23
timestamp 1667941163
transform 1 0 3220 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_35
timestamp 1667941163
transform 1 0 4324 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_47
timestamp 1667941163
transform 1 0 5428 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1667941163
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1667941163
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1667941163
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1667941163
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1667941163
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1667941163
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1667941163
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1667941163
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1667941163
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_137
timestamp 1667941163
transform 1 0 13708 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_145
timestamp 1667941163
transform 1 0 14444 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_67_153
timestamp 1667941163
transform 1 0 15180 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_67_166
timestamp 1667941163
transform 1 0 16376 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1667941163
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_181
timestamp 1667941163
transform 1 0 17756 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_190
timestamp 1667941163
transform 1 0 18584 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_202
timestamp 1667941163
transform 1 0 19688 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_208
timestamp 1667941163
transform 1 0 20240 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_216
timestamp 1667941163
transform 1 0 20976 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_225
timestamp 1667941163
transform 1 0 21804 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_233
timestamp 1667941163
transform 1 0 22540 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_67_249
timestamp 1667941163
transform 1 0 24012 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_260
timestamp 1667941163
transform 1 0 25024 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_272
timestamp 1667941163
transform 1 0 26128 0 -1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1667941163
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1667941163
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_305
timestamp 1667941163
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_317
timestamp 1667941163
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1667941163
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1667941163
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1667941163
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1667941163
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1667941163
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1667941163
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1667941163
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1667941163
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1667941163
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1667941163
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1667941163
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1667941163
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1667941163
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1667941163
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1667941163
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1667941163
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1667941163
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1667941163
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1667941163
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1667941163
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_505
timestamp 1667941163
transform 1 0 47564 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_67_510
timestamp 1667941163
transform 1 0 48024 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1667941163
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1667941163
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1667941163
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1667941163
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1667941163
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1667941163
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1667941163
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1667941163
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1667941163
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1667941163
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1667941163
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1667941163
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_121
timestamp 1667941163
transform 1 0 12236 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_129
timestamp 1667941163
transform 1 0 12972 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1667941163
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1667941163
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1667941163
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1667941163
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1667941163
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1667941163
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1667941163
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1667941163
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1667941163
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1667941163
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_238
timestamp 1667941163
transform 1 0 23000 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_242
timestamp 1667941163
transform 1 0 23368 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_250
timestamp 1667941163
transform 1 0 24104 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_253
timestamp 1667941163
transform 1 0 24380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_260
timestamp 1667941163
transform 1 0 25024 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_267
timestamp 1667941163
transform 1 0 25668 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_279
timestamp 1667941163
transform 1 0 26772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_291
timestamp 1667941163
transform 1 0 27876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_303
timestamp 1667941163
transform 1 0 28980 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1667941163
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1667941163
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1667941163
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1667941163
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1667941163
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1667941163
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1667941163
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1667941163
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1667941163
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1667941163
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1667941163
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1667941163
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1667941163
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1667941163
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1667941163
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1667941163
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1667941163
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1667941163
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1667941163
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1667941163
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_489
timestamp 1667941163
transform 1 0 46092 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_514
timestamp 1667941163
transform 1 0 48392 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1667941163
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1667941163
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1667941163
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1667941163
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1667941163
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1667941163
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1667941163
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1667941163
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1667941163
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1667941163
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1667941163
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1667941163
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1667941163
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_125
timestamp 1667941163
transform 1 0 12604 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_150
timestamp 1667941163
transform 1 0 14904 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_158
timestamp 1667941163
transform 1 0 15640 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_164
timestamp 1667941163
transform 1 0 16192 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_169
timestamp 1667941163
transform 1 0 16652 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_177
timestamp 1667941163
transform 1 0 17388 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_200
timestamp 1667941163
transform 1 0 19504 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_212
timestamp 1667941163
transform 1 0 20608 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_225
timestamp 1667941163
transform 1 0 21804 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_232
timestamp 1667941163
transform 1 0 22448 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_240
timestamp 1667941163
transform 1 0 23184 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_250
timestamp 1667941163
transform 1 0 24104 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_258
timestamp 1667941163
transform 1 0 24840 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_270
timestamp 1667941163
transform 1 0 25944 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_278
timestamp 1667941163
transform 1 0 26680 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1667941163
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1667941163
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1667941163
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1667941163
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1667941163
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1667941163
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1667941163
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1667941163
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1667941163
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1667941163
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1667941163
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1667941163
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1667941163
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1667941163
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1667941163
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1667941163
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1667941163
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1667941163
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1667941163
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1667941163
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1667941163
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1667941163
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_497
timestamp 1667941163
transform 1 0 46828 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_502
timestamp 1667941163
transform 1 0 47288 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_505
timestamp 1667941163
transform 1 0 47564 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_510
timestamp 1667941163
transform 1 0 48024 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1667941163
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1667941163
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1667941163
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1667941163
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1667941163
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1667941163
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1667941163
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1667941163
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1667941163
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1667941163
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1667941163
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1667941163
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1667941163
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1667941163
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1667941163
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1667941163
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_153
timestamp 1667941163
transform 1 0 15180 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_159
timestamp 1667941163
transform 1 0 15732 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_181
timestamp 1667941163
transform 1 0 17756 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_188
timestamp 1667941163
transform 1 0 18400 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1667941163
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1667941163
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1667941163
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1667941163
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_248
timestamp 1667941163
transform 1 0 23920 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1667941163
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1667941163
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_277
timestamp 1667941163
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_289
timestamp 1667941163
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1667941163
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1667941163
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1667941163
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_321
timestamp 1667941163
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_333
timestamp 1667941163
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_345
timestamp 1667941163
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1667941163
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1667941163
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1667941163
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1667941163
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1667941163
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1667941163
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1667941163
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1667941163
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1667941163
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1667941163
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1667941163
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1667941163
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1667941163
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1667941163
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1667941163
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_489
timestamp 1667941163
transform 1 0 46092 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_514
timestamp 1667941163
transform 1 0 48392 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1667941163
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1667941163
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1667941163
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1667941163
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1667941163
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1667941163
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_57
timestamp 1667941163
transform 1 0 6348 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_62
timestamp 1667941163
transform 1 0 6808 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_74
timestamp 1667941163
transform 1 0 7912 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_86
timestamp 1667941163
transform 1 0 9016 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_98
timestamp 1667941163
transform 1 0 10120 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_110
timestamp 1667941163
transform 1 0 11224 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1667941163
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1667941163
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1667941163
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1667941163
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1667941163
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1667941163
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1667941163
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1667941163
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1667941163
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1667941163
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1667941163
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1667941163
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1667941163
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1667941163
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1667941163
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1667941163
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1667941163
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1667941163
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1667941163
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1667941163
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1667941163
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1667941163
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1667941163
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1667941163
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1667941163
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1667941163
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1667941163
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1667941163
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1667941163
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1667941163
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1667941163
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1667941163
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1667941163
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1667941163
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1667941163
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1667941163
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1667941163
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1667941163
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1667941163
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1667941163
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_497
timestamp 1667941163
transform 1 0 46828 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_502
timestamp 1667941163
transform 1 0 47288 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_505
timestamp 1667941163
transform 1 0 47564 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_510
timestamp 1667941163
transform 1 0 48024 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1667941163
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1667941163
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1667941163
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1667941163
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_41
timestamp 1667941163
transform 1 0 4876 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_68
timestamp 1667941163
transform 1 0 7360 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_80
timestamp 1667941163
transform 1 0 8464 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1667941163
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1667941163
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1667941163
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1667941163
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1667941163
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1667941163
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1667941163
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1667941163
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1667941163
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1667941163
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1667941163
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1667941163
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1667941163
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1667941163
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1667941163
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1667941163
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1667941163
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1667941163
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1667941163
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1667941163
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_277
timestamp 1667941163
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_289
timestamp 1667941163
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1667941163
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1667941163
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1667941163
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1667941163
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1667941163
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1667941163
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1667941163
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1667941163
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1667941163
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1667941163
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1667941163
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1667941163
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1667941163
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1667941163
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1667941163
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1667941163
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1667941163
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1667941163
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1667941163
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1667941163
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1667941163
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_489
timestamp 1667941163
transform 1 0 46092 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_514
timestamp 1667941163
transform 1 0 48392 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1667941163
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1667941163
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1667941163
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_39
timestamp 1667941163
transform 1 0 4692 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_73_50
timestamp 1667941163
transform 1 0 5704 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1667941163
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1667941163
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1667941163
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1667941163
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1667941163
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1667941163
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1667941163
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1667941163
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1667941163
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1667941163
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1667941163
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1667941163
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1667941163
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1667941163
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1667941163
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1667941163
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1667941163
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1667941163
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1667941163
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1667941163
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1667941163
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 1667941163
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1667941163
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1667941163
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_281
timestamp 1667941163
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_293
timestamp 1667941163
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_305
timestamp 1667941163
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_317
timestamp 1667941163
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1667941163
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1667941163
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1667941163
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1667941163
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1667941163
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1667941163
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1667941163
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1667941163
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1667941163
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1667941163
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1667941163
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1667941163
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1667941163
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1667941163
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1667941163
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1667941163
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1667941163
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1667941163
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1667941163
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1667941163
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_505
timestamp 1667941163
transform 1 0 47564 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_73_510
timestamp 1667941163
transform 1 0 48024 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_74_3
timestamp 1667941163
transform 1 0 1380 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_11
timestamp 1667941163
transform 1 0 2116 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_16
timestamp 1667941163
transform 1 0 2576 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_23
timestamp 1667941163
transform 1 0 3220 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1667941163
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1667941163
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_41
timestamp 1667941163
transform 1 0 4876 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_52
timestamp 1667941163
transform 1 0 5888 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_64
timestamp 1667941163
transform 1 0 6992 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_76
timestamp 1667941163
transform 1 0 8096 0 1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1667941163
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1667941163
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1667941163
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1667941163
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1667941163
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1667941163
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1667941163
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1667941163
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1667941163
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1667941163
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1667941163
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1667941163
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1667941163
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1667941163
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1667941163
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1667941163
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1667941163
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1667941163
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1667941163
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1667941163
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_277
timestamp 1667941163
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_289
timestamp 1667941163
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1667941163
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1667941163
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1667941163
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1667941163
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1667941163
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_345
timestamp 1667941163
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1667941163
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1667941163
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1667941163
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1667941163
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_389
timestamp 1667941163
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_401
timestamp 1667941163
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1667941163
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1667941163
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1667941163
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1667941163
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1667941163
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1667941163
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1667941163
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1667941163
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1667941163
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_489
timestamp 1667941163
transform 1 0 46092 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_514
timestamp 1667941163
transform 1 0 48392 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_75_3
timestamp 1667941163
transform 1 0 1380 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_9
timestamp 1667941163
transform 1 0 1932 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_31
timestamp 1667941163
transform 1 0 3956 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_47
timestamp 1667941163
transform 1 0 5428 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_54
timestamp 1667941163
transform 1 0 6072 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1667941163
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1667941163
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1667941163
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1667941163
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1667941163
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1667941163
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1667941163
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1667941163
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1667941163
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1667941163
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1667941163
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1667941163
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1667941163
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1667941163
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1667941163
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1667941163
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1667941163
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1667941163
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1667941163
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1667941163
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1667941163
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1667941163
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1667941163
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1667941163
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1667941163
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1667941163
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1667941163
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1667941163
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1667941163
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1667941163
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1667941163
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1667941163
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1667941163
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_373
timestamp 1667941163
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1667941163
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1667941163
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1667941163
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1667941163
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1667941163
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1667941163
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1667941163
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1667941163
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1667941163
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1667941163
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1667941163
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1667941163
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_497
timestamp 1667941163
transform 1 0 46828 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_502
timestamp 1667941163
transform 1 0 47288 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_505
timestamp 1667941163
transform 1 0 47564 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_75_510
timestamp 1667941163
transform 1 0 48024 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_76_3
timestamp 1667941163
transform 1 0 1380 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_10
timestamp 1667941163
transform 1 0 2024 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_26
timestamp 1667941163
transform 1 0 3496 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_29
timestamp 1667941163
transform 1 0 3772 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_43
timestamp 1667941163
transform 1 0 5060 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_68
timestamp 1667941163
transform 1 0 7360 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_80
timestamp 1667941163
transform 1 0 8464 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1667941163
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1667941163
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1667941163
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1667941163
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1667941163
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1667941163
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1667941163
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1667941163
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1667941163
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1667941163
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1667941163
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1667941163
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1667941163
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1667941163
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1667941163
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1667941163
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1667941163
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1667941163
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1667941163
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1667941163
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1667941163
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_289
timestamp 1667941163
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1667941163
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1667941163
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1667941163
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1667941163
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1667941163
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1667941163
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1667941163
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1667941163
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1667941163
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1667941163
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1667941163
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1667941163
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1667941163
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1667941163
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1667941163
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1667941163
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1667941163
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1667941163
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1667941163
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1667941163
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1667941163
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1667941163
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1667941163
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_513
timestamp 1667941163
transform 1 0 48300 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_77_3
timestamp 1667941163
transform 1 0 1380 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_9
timestamp 1667941163
transform 1 0 1932 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_31
timestamp 1667941163
transform 1 0 3956 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_38
timestamp 1667941163
transform 1 0 4600 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_54
timestamp 1667941163
transform 1 0 6072 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_57
timestamp 1667941163
transform 1 0 6348 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_62
timestamp 1667941163
transform 1 0 6808 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_74
timestamp 1667941163
transform 1 0 7912 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_86
timestamp 1667941163
transform 1 0 9016 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_98
timestamp 1667941163
transform 1 0 10120 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_110
timestamp 1667941163
transform 1 0 11224 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1667941163
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1667941163
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1667941163
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1667941163
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1667941163
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1667941163
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1667941163
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1667941163
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1667941163
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1667941163
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1667941163
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1667941163
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1667941163
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1667941163
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1667941163
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1667941163
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1667941163
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1667941163
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1667941163
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1667941163
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1667941163
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1667941163
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1667941163
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1667941163
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1667941163
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1667941163
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1667941163
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1667941163
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1667941163
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1667941163
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1667941163
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1667941163
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1667941163
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1667941163
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1667941163
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1667941163
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1667941163
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1667941163
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1667941163
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1667941163
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_497
timestamp 1667941163
transform 1 0 46828 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_502
timestamp 1667941163
transform 1 0 47288 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_505
timestamp 1667941163
transform 1 0 47564 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_77_510
timestamp 1667941163
transform 1 0 48024 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_78_3
timestamp 1667941163
transform 1 0 1380 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_10
timestamp 1667941163
transform 1 0 2024 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_26
timestamp 1667941163
transform 1 0 3496 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_29
timestamp 1667941163
transform 1 0 3772 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_51
timestamp 1667941163
transform 1 0 5796 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_67
timestamp 1667941163
transform 1 0 7268 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_79
timestamp 1667941163
transform 1 0 8372 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1667941163
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1667941163
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1667941163
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1667941163
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1667941163
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1667941163
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1667941163
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1667941163
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1667941163
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1667941163
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1667941163
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1667941163
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1667941163
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1667941163
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1667941163
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1667941163
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1667941163
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1667941163
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1667941163
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1667941163
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1667941163
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1667941163
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1667941163
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1667941163
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1667941163
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1667941163
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1667941163
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1667941163
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1667941163
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1667941163
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1667941163
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1667941163
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1667941163
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 1667941163
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_401
timestamp 1667941163
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1667941163
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1667941163
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_421
timestamp 1667941163
transform 1 0 39836 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_425
timestamp 1667941163
transform 1 0 40204 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_429
timestamp 1667941163
transform 1 0 40572 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_441
timestamp 1667941163
transform 1 0 41676 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_453
timestamp 1667941163
transform 1 0 42780 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_465
timestamp 1667941163
transform 1 0 43884 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_473
timestamp 1667941163
transform 1 0 44620 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1667941163
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_489
timestamp 1667941163
transform 1 0 46092 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_514
timestamp 1667941163
transform 1 0 48392 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_3
timestamp 1667941163
transform 1 0 1380 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_79_32
timestamp 1667941163
transform 1 0 4048 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_52
timestamp 1667941163
transform 1 0 5888 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_57
timestamp 1667941163
transform 1 0 6348 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_71
timestamp 1667941163
transform 1 0 7636 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_83
timestamp 1667941163
transform 1 0 8740 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_95
timestamp 1667941163
transform 1 0 9844 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_101
timestamp 1667941163
transform 1 0 10396 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1667941163
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1667941163
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1667941163
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1667941163
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_137
timestamp 1667941163
transform 1 0 13708 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_148
timestamp 1667941163
transform 1 0 14720 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_155
timestamp 1667941163
transform 1 0 15364 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1667941163
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1667941163
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1667941163
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1667941163
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1667941163
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1667941163
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1667941163
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1667941163
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1667941163
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_249
timestamp 1667941163
transform 1 0 24012 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_253
timestamp 1667941163
transform 1 0 24380 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_257
timestamp 1667941163
transform 1 0 24748 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_264
timestamp 1667941163
transform 1 0 25392 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_276
timestamp 1667941163
transform 1 0 26496 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1667941163
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1667941163
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_305
timestamp 1667941163
transform 1 0 29164 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_311
timestamp 1667941163
transform 1 0 29716 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_315
timestamp 1667941163
transform 1 0 30084 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_327
timestamp 1667941163
transform 1 0 31188 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1667941163
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1667941163
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1667941163
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1667941163
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_373
timestamp 1667941163
transform 1 0 35420 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_377
timestamp 1667941163
transform 1 0 35788 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_384
timestamp 1667941163
transform 1 0 36432 0 -1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1667941163
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_405
timestamp 1667941163
transform 1 0 38364 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_79_432
timestamp 1667941163
transform 1 0 40848 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_438
timestamp 1667941163
transform 1 0 41400 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_442
timestamp 1667941163
transform 1 0 41768 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1667941163
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1667941163
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1667941163
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_485
timestamp 1667941163
transform 1 0 45724 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_490
timestamp 1667941163
transform 1 0 46184 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_498
timestamp 1667941163
transform 1 0 46920 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_502
timestamp 1667941163
transform 1 0 47288 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_505
timestamp 1667941163
transform 1 0 47564 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_79_510
timestamp 1667941163
transform 1 0 48024 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_80_3
timestamp 1667941163
transform 1 0 1380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_26
timestamp 1667941163
transform 1 0 3496 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_29
timestamp 1667941163
transform 1 0 3772 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_51
timestamp 1667941163
transform 1 0 5796 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_58
timestamp 1667941163
transform 1 0 6440 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1667941163
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1667941163
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1667941163
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1667941163
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_97
timestamp 1667941163
transform 1 0 10028 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_101
timestamp 1667941163
transform 1 0 10396 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_123
timestamp 1667941163
transform 1 0 12420 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_130
timestamp 1667941163
transform 1 0 13064 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_134
timestamp 1667941163
transform 1 0 13432 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_138
timestamp 1667941163
transform 1 0 13800 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_80_141
timestamp 1667941163
transform 1 0 14076 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_147
timestamp 1667941163
transform 1 0 14628 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_172
timestamp 1667941163
transform 1 0 16928 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_184
timestamp 1667941163
transform 1 0 18032 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1667941163
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1667941163
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1667941163
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_236
timestamp 1667941163
transform 1 0 22816 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_244
timestamp 1667941163
transform 1 0 23552 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_80_250
timestamp 1667941163
transform 1 0 24104 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_253
timestamp 1667941163
transform 1 0 24380 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_276
timestamp 1667941163
transform 1 0 26496 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_288
timestamp 1667941163
transform 1 0 27600 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_300
timestamp 1667941163
transform 1 0 28704 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_80_306
timestamp 1667941163
transform 1 0 29256 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_309
timestamp 1667941163
transform 1 0 29532 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_332
timestamp 1667941163
transform 1 0 31648 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_344
timestamp 1667941163
transform 1 0 32752 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_351
timestamp 1667941163
transform 1 0 33396 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1667941163
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_365
timestamp 1667941163
transform 1 0 34684 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_371
timestamp 1667941163
transform 1 0 35236 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_393
timestamp 1667941163
transform 1 0 37260 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_401
timestamp 1667941163
transform 1 0 37996 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_407
timestamp 1667941163
transform 1 0 38548 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_414
timestamp 1667941163
transform 1 0 39192 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_80_421
timestamp 1667941163
transform 1 0 39836 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1667941163
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1667941163
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1667941163
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1667941163
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_477
timestamp 1667941163
transform 1 0 44988 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_482
timestamp 1667941163
transform 1 0 45448 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_489
timestamp 1667941163
transform 1 0 46092 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_514
timestamp 1667941163
transform 1 0 48392 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_3
timestamp 1667941163
transform 1 0 1380 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_7
timestamp 1667941163
transform 1 0 1748 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_29
timestamp 1667941163
transform 1 0 3772 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_54
timestamp 1667941163
transform 1 0 6072 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_57
timestamp 1667941163
transform 1 0 6348 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_62
timestamp 1667941163
transform 1 0 6808 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1667941163
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1667941163
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_93
timestamp 1667941163
transform 1 0 9660 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_101
timestamp 1667941163
transform 1 0 10396 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1667941163
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1667941163
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_113
timestamp 1667941163
transform 1 0 11500 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_140
timestamp 1667941163
transform 1 0 13984 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_165
timestamp 1667941163
transform 1 0 16284 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_81_169
timestamp 1667941163
transform 1 0 16652 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_174
timestamp 1667941163
transform 1 0 17112 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_186
timestamp 1667941163
transform 1 0 18216 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_198
timestamp 1667941163
transform 1 0 19320 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_210
timestamp 1667941163
transform 1 0 20424 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_222
timestamp 1667941163
transform 1 0 21528 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_81_225
timestamp 1667941163
transform 1 0 21804 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_231
timestamp 1667941163
transform 1 0 22356 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_253
timestamp 1667941163
transform 1 0 24380 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_278
timestamp 1667941163
transform 1 0 26680 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1667941163
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_293
timestamp 1667941163
transform 1 0 28060 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_297
timestamp 1667941163
transform 1 0 28428 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_301
timestamp 1667941163
transform 1 0 28796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_326
timestamp 1667941163
transform 1 0 31096 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_334
timestamp 1667941163
transform 1 0 31832 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_337
timestamp 1667941163
transform 1 0 32108 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_345
timestamp 1667941163
transform 1 0 32844 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_368
timestamp 1667941163
transform 1 0 34960 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_372
timestamp 1667941163
transform 1 0 35328 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_376
timestamp 1667941163
transform 1 0 35696 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_383
timestamp 1667941163
transform 1 0 36340 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1667941163
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_393
timestamp 1667941163
transform 1 0 37260 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_416
timestamp 1667941163
transform 1 0 39376 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1667941163
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1667941163
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_449
timestamp 1667941163
transform 1 0 42412 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_472
timestamp 1667941163
transform 1 0 44528 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_480
timestamp 1667941163
transform 1 0 45264 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_502
timestamp 1667941163
transform 1 0 47288 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_505
timestamp 1667941163
transform 1 0 47564 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_81_510
timestamp 1667941163
transform 1 0 48024 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_82_3
timestamp 1667941163
transform 1 0 1380 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_9
timestamp 1667941163
transform 1 0 1932 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_19
timestamp 1667941163
transform 1 0 2852 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_26
timestamp 1667941163
transform 1 0 3496 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_29
timestamp 1667941163
transform 1 0 3772 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_37
timestamp 1667941163
transform 1 0 4508 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_44
timestamp 1667941163
transform 1 0 5152 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_51
timestamp 1667941163
transform 1 0 5796 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_55
timestamp 1667941163
transform 1 0 6164 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_57
timestamp 1667941163
transform 1 0 6348 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_62
timestamp 1667941163
transform 1 0 6808 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_74
timestamp 1667941163
transform 1 0 7912 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_82
timestamp 1667941163
transform 1 0 8648 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_85
timestamp 1667941163
transform 1 0 8924 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_90
timestamp 1667941163
transform 1 0 9384 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_102
timestamp 1667941163
transform 1 0 10488 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_110
timestamp 1667941163
transform 1 0 11224 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_113
timestamp 1667941163
transform 1 0 11500 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_121
timestamp 1667941163
transform 1 0 12236 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_126
timestamp 1667941163
transform 1 0 12696 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_134
timestamp 1667941163
transform 1 0 13432 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_138
timestamp 1667941163
transform 1 0 13800 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_141
timestamp 1667941163
transform 1 0 14076 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_164
timestamp 1667941163
transform 1 0 16192 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_169
timestamp 1667941163
transform 1 0 16652 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_177
timestamp 1667941163
transform 1 0 17388 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_182
timestamp 1667941163
transform 1 0 17848 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_194
timestamp 1667941163
transform 1 0 18952 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_197
timestamp 1667941163
transform 1 0 19228 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_203
timestamp 1667941163
transform 1 0 19780 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_215
timestamp 1667941163
transform 1 0 20884 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_223
timestamp 1667941163
transform 1 0 21620 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_225
timestamp 1667941163
transform 1 0 21804 0 1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_82_236
timestamp 1667941163
transform 1 0 22816 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_248
timestamp 1667941163
transform 1 0 23920 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_253
timestamp 1667941163
transform 1 0 24380 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_259
timestamp 1667941163
transform 1 0 24932 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_266
timestamp 1667941163
transform 1 0 25576 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_278
timestamp 1667941163
transform 1 0 26680 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_281
timestamp 1667941163
transform 1 0 26956 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_293
timestamp 1667941163
transform 1 0 28060 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_305
timestamp 1667941163
transform 1 0 29164 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_82_309
timestamp 1667941163
transform 1 0 29532 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_315
timestamp 1667941163
transform 1 0 30084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_327
timestamp 1667941163
transform 1 0 31188 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_335
timestamp 1667941163
transform 1 0 31924 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_337
timestamp 1667941163
transform 1 0 32108 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_343
timestamp 1667941163
transform 1 0 32660 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_347
timestamp 1667941163
transform 1 0 33028 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_351
timestamp 1667941163
transform 1 0 33396 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1667941163
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1667941163
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1667941163
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_389
timestamp 1667941163
transform 1 0 36892 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_393
timestamp 1667941163
transform 1 0 37260 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_401
timestamp 1667941163
transform 1 0 37996 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_405
timestamp 1667941163
transform 1 0 38364 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_82_414
timestamp 1667941163
transform 1 0 39192 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_82_421
timestamp 1667941163
transform 1 0 39836 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_427
timestamp 1667941163
transform 1 0 40388 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_435
timestamp 1667941163
transform 1 0 41124 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_440
timestamp 1667941163
transform 1 0 41584 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_449
timestamp 1667941163
transform 1 0 42412 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_455
timestamp 1667941163
transform 1 0 42964 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_467
timestamp 1667941163
transform 1 0 44068 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1667941163
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_477
timestamp 1667941163
transform 1 0 44988 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_502
timestamp 1667941163
transform 1 0 47288 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_82_505
timestamp 1667941163
transform 1 0 47564 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_82_514
timestamp 1667941163
transform 1 0 48392 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1667941163
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1667941163
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1667941163
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1667941163
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1667941163
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1667941163
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1667941163
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1667941163
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1667941163
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1667941163
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1667941163
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1667941163
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1667941163
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1667941163
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1667941163
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1667941163
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1667941163
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1667941163
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1667941163
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1667941163
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1667941163
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1667941163
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1667941163
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1667941163
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1667941163
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1667941163
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1667941163
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1667941163
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1667941163
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1667941163
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1667941163
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1667941163
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1667941163
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1667941163
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1667941163
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1667941163
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1667941163
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1667941163
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1667941163
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1667941163
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1667941163
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1667941163
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1667941163
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1667941163
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1667941163
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1667941163
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1667941163
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1667941163
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1667941163
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1667941163
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1667941163
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1667941163
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1667941163
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1667941163
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1667941163
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1667941163
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1667941163
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1667941163
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1667941163
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1667941163
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1667941163
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1667941163
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1667941163
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1667941163
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1667941163
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1667941163
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1667941163
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1667941163
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1667941163
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1667941163
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1667941163
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1667941163
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1667941163
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1667941163
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1667941163
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1667941163
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1667941163
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1667941163
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1667941163
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1667941163
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1667941163
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1667941163
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1667941163
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1667941163
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1667941163
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1667941163
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1667941163
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1667941163
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1667941163
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1667941163
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1667941163
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1667941163
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1667941163
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1667941163
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1667941163
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1667941163
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1667941163
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1667941163
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1667941163
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1667941163
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1667941163
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1667941163
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1667941163
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1667941163
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1667941163
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1667941163
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1667941163
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1667941163
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1667941163
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1667941163
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1667941163
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1667941163
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1667941163
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1667941163
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1667941163
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1667941163
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1667941163
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1667941163
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1667941163
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1667941163
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1667941163
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1667941163
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1667941163
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1667941163
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1667941163
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1667941163
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1667941163
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1667941163
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1667941163
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1667941163
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1667941163
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1667941163
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1667941163
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1667941163
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1667941163
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1667941163
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1667941163
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1667941163
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1667941163
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1667941163
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1667941163
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1667941163
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1667941163
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1667941163
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1667941163
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1667941163
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1667941163
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1667941163
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1667941163
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1667941163
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1667941163
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1667941163
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1667941163
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1667941163
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1667941163
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1667941163
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1667941163
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1667941163
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1667941163
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1667941163
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1667941163
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1667941163
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1667941163
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1667941163
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1667941163
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1667941163
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1667941163
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1667941163
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1667941163
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1667941163
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1667941163
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1667941163
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1667941163
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1667941163
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1667941163
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1667941163
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1667941163
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1667941163
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1667941163
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1667941163
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1667941163
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1667941163
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1667941163
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1667941163
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1667941163
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1667941163
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1667941163
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1667941163
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1667941163
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1667941163
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1667941163
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1667941163
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1667941163
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1667941163
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1667941163
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1667941163
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1667941163
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1667941163
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1667941163
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1667941163
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1667941163
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1667941163
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1667941163
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1667941163
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1667941163
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1667941163
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1667941163
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1667941163
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1667941163
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1667941163
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1667941163
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1667941163
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1667941163
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1667941163
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1667941163
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1667941163
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1667941163
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1667941163
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1667941163
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1667941163
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1667941163
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1667941163
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1667941163
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1667941163
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1667941163
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1667941163
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1667941163
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1667941163
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1667941163
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1667941163
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1667941163
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1667941163
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1667941163
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1667941163
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1667941163
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1667941163
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1667941163
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1667941163
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1667941163
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1667941163
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1667941163
transform 1 0 42320 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1667941163
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1667941163
transform 1 0 47472 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0956_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 5612 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _0957_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 9108 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0958_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0959_
timestamp 1667941163
transform 1 0 7636 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0960_
timestamp 1667941163
transform 1 0 9108 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0961_
timestamp 1667941163
transform -1 0 7176 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0962_
timestamp 1667941163
transform -1 0 6072 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0963_
timestamp 1667941163
transform -1 0 5612 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0964_
timestamp 1667941163
transform -1 0 4416 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0965_
timestamp 1667941163
transform 1 0 5152 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0966_
timestamp 1667941163
transform 1 0 5980 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0967_
timestamp 1667941163
transform 1 0 4968 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0968_
timestamp 1667941163
transform 1 0 5704 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0969_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 10396 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0970_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 5336 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0971_
timestamp 1667941163
transform 1 0 9200 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0972_
timestamp 1667941163
transform -1 0 9108 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0973_
timestamp 1667941163
transform -1 0 8372 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0974_
timestamp 1667941163
transform -1 0 6992 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0975_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 7452 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0976_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6808 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  _0977_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 2852 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  _0978_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 3496 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  _0979_
timestamp 1667941163
transform 1 0 6532 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0980_
timestamp 1667941163
transform -1 0 47288 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0981_
timestamp 1667941163
transform 1 0 6532 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0982_
timestamp 1667941163
transform 1 0 47748 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0983_
timestamp 1667941163
transform -1 0 46092 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0984_
timestamp 1667941163
transform -1 0 47104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp 1667941163
transform 1 0 6532 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0986_
timestamp 1667941163
transform -1 0 40572 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0987_
timestamp 1667941163
transform -1 0 6072 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0988_
timestamp 1667941163
transform -1 0 32568 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0989_
timestamp 1667941163
transform 1 0 47748 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0990_
timestamp 1667941163
transform 1 0 4324 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1667941163
transform 1 0 27140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0992_
timestamp 1667941163
transform 1 0 36156 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0993_
timestamp 1667941163
transform -1 0 4232 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0994_
timestamp 1667941163
transform 1 0 38272 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0995_
timestamp 1667941163
transform -1 0 17664 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0996_
timestamp 1667941163
transform 1 0 43056 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0997_
timestamp 1667941163
transform -1 0 2576 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0998_
timestamp 1667941163
transform -1 0 2576 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0999_
timestamp 1667941163
transform -1 0 4600 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1000_
timestamp 1667941163
transform 1 0 42964 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1001_
timestamp 1667941163
transform 1 0 6164 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1002_
timestamp 1667941163
transform -1 0 47288 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1003_
timestamp 1667941163
transform 1 0 47748 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1004_
timestamp 1667941163
transform 1 0 15088 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1005_
timestamp 1667941163
transform 1 0 47748 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1006_
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1007_
timestamp 1667941163
transform 1 0 41492 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1008_
timestamp 1667941163
transform -1 0 25576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1009_
timestamp 1667941163
transform -1 0 47288 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1010_
timestamp 1667941163
transform -1 0 4692 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1011_
timestamp 1667941163
transform 1 0 47748 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1012_
timestamp 1667941163
transform 1 0 2392 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1013_
timestamp 1667941163
transform -1 0 13064 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1014_
timestamp 1667941163
transform 1 0 4048 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1015_
timestamp 1667941163
transform 1 0 10488 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1016_
timestamp 1667941163
transform -1 0 3036 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1017_
timestamp 1667941163
transform -1 0 47288 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1018_
timestamp 1667941163
transform 1 0 47748 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1019_
timestamp 1667941163
transform 1 0 47748 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1020_
timestamp 1667941163
transform 1 0 2944 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1021_
timestamp 1667941163
transform 1 0 13524 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1022_
timestamp 1667941163
transform -1 0 47748 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1023_
timestamp 1667941163
transform 1 0 4784 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1024_
timestamp 1667941163
transform 1 0 13156 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1025_
timestamp 1667941163
transform -1 0 35788 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1026_
timestamp 1667941163
transform 1 0 14352 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1027_
timestamp 1667941163
transform 1 0 46368 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1028_
timestamp 1667941163
transform -1 0 6440 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1667941163
transform -1 0 4876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1030_
timestamp 1667941163
transform 1 0 23828 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1031_
timestamp 1667941163
transform -1 0 25392 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1032_
timestamp 1667941163
transform 1 0 46368 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1033_
timestamp 1667941163
transform 1 0 47748 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _1034_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3956 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _1035_
timestamp 1667941163
transform 1 0 28980 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1036_
timestamp 1667941163
transform -1 0 43148 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1037_
timestamp 1667941163
transform 1 0 46920 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1038_
timestamp 1667941163
transform -1 0 3496 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1039_
timestamp 1667941163
transform -1 0 41584 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1040_
timestamp 1667941163
transform -1 0 2668 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1041_
timestamp 1667941163
transform -1 0 45724 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1042_
timestamp 1667941163
transform 1 0 10488 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1043_
timestamp 1667941163
transform -1 0 2668 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1044_
timestamp 1667941163
transform 1 0 7544 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1045_
timestamp 1667941163
transform -1 0 5060 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1046_
timestamp 1667941163
transform -1 0 2484 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1047_
timestamp 1667941163
transform -1 0 3220 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1048_
timestamp 1667941163
transform -1 0 2484 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1049_
timestamp 1667941163
transform 1 0 19412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1050_
timestamp 1667941163
transform -1 0 3036 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1051_
timestamp 1667941163
transform 1 0 47748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1052_
timestamp 1667941163
transform -1 0 4232 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1053_
timestamp 1667941163
transform 1 0 46184 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1054_
timestamp 1667941163
transform 1 0 6716 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1055_
timestamp 1667941163
transform 1 0 44712 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1056_
timestamp 1667941163
transform 1 0 5060 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1057_
timestamp 1667941163
transform -1 0 45816 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1058_
timestamp 1667941163
transform -1 0 46920 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1059_
timestamp 1667941163
transform -1 0 22264 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1060_
timestamp 1667941163
transform 1 0 15916 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1061_
timestamp 1667941163
transform 1 0 13064 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1062_
timestamp 1667941163
transform -1 0 18400 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1063_
timestamp 1667941163
transform -1 0 5704 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1064_
timestamp 1667941163
transform 1 0 47748 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1065_
timestamp 1667941163
transform 1 0 47748 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1066_
timestamp 1667941163
transform -1 0 6072 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _1067_
timestamp 1667941163
transform -1 0 5796 0 1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _1068_
timestamp 1667941163
transform 1 0 46368 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1069_
timestamp 1667941163
transform -1 0 3036 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1070_
timestamp 1667941163
transform 1 0 47748 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1071_
timestamp 1667941163
transform 1 0 29808 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1072_
timestamp 1667941163
transform -1 0 12604 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1073_
timestamp 1667941163
transform -1 0 47288 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1074_
timestamp 1667941163
transform -1 0 4692 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1075_
timestamp 1667941163
transform 1 0 47748 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1076_
timestamp 1667941163
transform -1 0 7084 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1077_
timestamp 1667941163
transform 1 0 45172 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1078_
timestamp 1667941163
transform 1 0 4968 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1079_
timestamp 1667941163
transform 1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1080_
timestamp 1667941163
transform 1 0 46368 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1081_
timestamp 1667941163
transform 1 0 47748 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1082_
timestamp 1667941163
transform 1 0 33120 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1083_
timestamp 1667941163
transform -1 0 47288 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1084_
timestamp 1667941163
transform 1 0 6624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1085_
timestamp 1667941163
transform 1 0 18584 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1086_
timestamp 1667941163
transform -1 0 5244 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1087_
timestamp 1667941163
transform 1 0 47748 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1088_
timestamp 1667941163
transform 1 0 47748 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1089_
timestamp 1667941163
transform -1 0 2576 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1090_
timestamp 1667941163
transform 1 0 22540 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1091_
timestamp 1667941163
transform -1 0 2576 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1092_
timestamp 1667941163
transform -1 0 5520 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1093_
timestamp 1667941163
transform 1 0 2760 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1094_
timestamp 1667941163
transform 1 0 38088 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1095_
timestamp 1667941163
transform -1 0 26220 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1096_
timestamp 1667941163
transform 1 0 38916 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1097_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 7636 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1098_
timestamp 1667941163
transform -1 0 11132 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1099_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 9384 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1100_
timestamp 1667941163
transform 1 0 10028 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1101_
timestamp 1667941163
transform 1 0 10488 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1102_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1103_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 13156 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1104_
timestamp 1667941163
transform 1 0 12880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1105_
timestamp 1667941163
transform 1 0 13064 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1106_
timestamp 1667941163
transform 1 0 12420 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1107_
timestamp 1667941163
transform 1 0 11684 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1108_
timestamp 1667941163
transform 1 0 10304 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1109_
timestamp 1667941163
transform -1 0 11132 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1110_
timestamp 1667941163
transform 1 0 10764 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1111_
timestamp 1667941163
transform 1 0 9752 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1112_
timestamp 1667941163
transform 1 0 8372 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1113_
timestamp 1667941163
transform 1 0 9108 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1114_
timestamp 1667941163
transform 1 0 8924 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1115_
timestamp 1667941163
transform -1 0 10764 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1116_
timestamp 1667941163
transform 1 0 10948 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1117_
timestamp 1667941163
transform 1 0 9660 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1118_
timestamp 1667941163
transform 1 0 8832 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1119_
timestamp 1667941163
transform 1 0 9108 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1120_
timestamp 1667941163
transform 1 0 7084 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1121_
timestamp 1667941163
transform 1 0 6716 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1122_
timestamp 1667941163
transform -1 0 6072 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1123_
timestamp 1667941163
transform -1 0 8556 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1124_
timestamp 1667941163
transform 1 0 6532 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1125_
timestamp 1667941163
transform -1 0 7360 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1126_
timestamp 1667941163
transform -1 0 7176 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1127_
timestamp 1667941163
transform -1 0 30452 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1128_
timestamp 1667941163
transform 1 0 29348 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _1129_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 32292 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1130_
timestamp 1667941163
transform -1 0 32936 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1131_
timestamp 1667941163
transform 1 0 29716 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1132_
timestamp 1667941163
transform 1 0 28888 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1133_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 30728 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1134_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 31556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _1135_
timestamp 1667941163
transform 1 0 41308 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1136_
timestamp 1667941163
transform -1 0 31648 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1137_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 31188 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1138_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 36892 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1139_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 31556 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1140_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 31556 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1141_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 33028 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1142_
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1143_
timestamp 1667941163
transform 1 0 33672 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1144_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 31556 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_2  _1145_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 32292 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1146_
timestamp 1667941163
transform 1 0 35604 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1147_
timestamp 1667941163
transform 1 0 37444 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1148_
timestamp 1667941163
transform -1 0 36432 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1149_
timestamp 1667941163
transform -1 0 36616 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1150_
timestamp 1667941163
transform -1 0 35604 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1151_
timestamp 1667941163
transform -1 0 36064 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1152_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 35788 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1153_
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1154_
timestamp 1667941163
transform 1 0 33672 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1155_
timestamp 1667941163
transform 1 0 35236 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1156_
timestamp 1667941163
transform 1 0 36248 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1157_
timestamp 1667941163
transform -1 0 35604 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1158_
timestamp 1667941163
transform 1 0 33580 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1159_
timestamp 1667941163
transform 1 0 33028 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1160_
timestamp 1667941163
transform 1 0 32752 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1161_
timestamp 1667941163
transform 1 0 39008 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1162_
timestamp 1667941163
transform -1 0 39376 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1163_
timestamp 1667941163
transform -1 0 39192 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1164_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 35420 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _1165_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 35880 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1166_
timestamp 1667941163
transform -1 0 38088 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1167_
timestamp 1667941163
transform 1 0 36064 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1168_
timestamp 1667941163
transform 1 0 37536 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1169_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 38916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1170_
timestamp 1667941163
transform 1 0 40756 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1171_
timestamp 1667941163
transform -1 0 40848 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1172_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 40204 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1173_
timestamp 1667941163
transform 1 0 37168 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1174_
timestamp 1667941163
transform 1 0 38180 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1175_
timestamp 1667941163
transform -1 0 39652 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1176_
timestamp 1667941163
transform 1 0 38640 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1177_
timestamp 1667941163
transform -1 0 38272 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1178_
timestamp 1667941163
transform 1 0 39100 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1179_
timestamp 1667941163
transform -1 0 40388 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1180_
timestamp 1667941163
transform 1 0 40112 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1181_
timestamp 1667941163
transform -1 0 40388 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1182_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 38824 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1183_
timestamp 1667941163
transform 1 0 39836 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1184_
timestamp 1667941163
transform -1 0 37720 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1185_
timestamp 1667941163
transform 1 0 36340 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1186_
timestamp 1667941163
transform -1 0 38272 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1187_
timestamp 1667941163
transform -1 0 39560 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1188_
timestamp 1667941163
transform -1 0 37352 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1189_
timestamp 1667941163
transform 1 0 35788 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1190_
timestamp 1667941163
transform 1 0 35420 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1191_
timestamp 1667941163
transform 1 0 35144 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1192_
timestamp 1667941163
transform -1 0 40848 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _1193_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37904 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1194_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37996 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _1195_
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1196_
timestamp 1667941163
transform 1 0 40020 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1197_
timestamp 1667941163
transform 1 0 39192 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1198_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 38088 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1199_
timestamp 1667941163
transform -1 0 38548 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1200_
timestamp 1667941163
transform -1 0 36524 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1201_
timestamp 1667941163
transform -1 0 36800 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1202_
timestamp 1667941163
transform -1 0 37720 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1203_
timestamp 1667941163
transform 1 0 37260 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1204_
timestamp 1667941163
transform -1 0 37812 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1205_
timestamp 1667941163
transform -1 0 36892 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1206_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 36892 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1207_
timestamp 1667941163
transform 1 0 33580 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1208_
timestamp 1667941163
transform -1 0 34040 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1209_
timestamp 1667941163
transform 1 0 35236 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1210_
timestamp 1667941163
transform -1 0 35788 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1211_
timestamp 1667941163
transform 1 0 31372 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1212_
timestamp 1667941163
transform 1 0 32568 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _1213_
timestamp 1667941163
transform -1 0 35420 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1214_
timestamp 1667941163
transform 1 0 33396 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1215_
timestamp 1667941163
transform 1 0 33672 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1216_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 34868 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1217_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 33948 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1218_
timestamp 1667941163
transform -1 0 33028 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1219_
timestamp 1667941163
transform -1 0 42044 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1220_
timestamp 1667941163
transform -1 0 34040 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1221_
timestamp 1667941163
transform 1 0 34868 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1222_
timestamp 1667941163
transform -1 0 35144 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1223_
timestamp 1667941163
transform -1 0 34960 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1224_
timestamp 1667941163
transform 1 0 34960 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1225_
timestamp 1667941163
transform 1 0 36340 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1226_
timestamp 1667941163
transform -1 0 36708 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1227_
timestamp 1667941163
transform 1 0 36340 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1228_
timestamp 1667941163
transform 1 0 35328 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1229_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 36524 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1230_
timestamp 1667941163
transform 1 0 37444 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1231_
timestamp 1667941163
transform -1 0 36616 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1232_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 35604 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _1233_
timestamp 1667941163
transform 1 0 34408 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1234_
timestamp 1667941163
transform 1 0 35328 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1235_
timestamp 1667941163
transform 1 0 36064 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1236_
timestamp 1667941163
transform 1 0 35512 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1237_
timestamp 1667941163
transform 1 0 35972 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1238_
timestamp 1667941163
transform 1 0 36616 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1239_
timestamp 1667941163
transform 1 0 37260 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1240_
timestamp 1667941163
transform 1 0 38272 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1241_
timestamp 1667941163
transform -1 0 34408 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1242_
timestamp 1667941163
transform -1 0 36892 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1243_
timestamp 1667941163
transform -1 0 34040 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1244_
timestamp 1667941163
transform 1 0 33028 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1245_
timestamp 1667941163
transform 1 0 34960 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1246_
timestamp 1667941163
transform -1 0 35696 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1247_
timestamp 1667941163
transform 1 0 32200 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1248_
timestamp 1667941163
transform -1 0 33396 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1249_
timestamp 1667941163
transform 1 0 35880 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1250_
timestamp 1667941163
transform 1 0 36156 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1251_
timestamp 1667941163
transform -1 0 35788 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1252_
timestamp 1667941163
transform -1 0 37260 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1253_
timestamp 1667941163
transform 1 0 36340 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1254_
timestamp 1667941163
transform 1 0 36340 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1255_
timestamp 1667941163
transform 1 0 37444 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1256_
timestamp 1667941163
transform 1 0 37352 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1257_
timestamp 1667941163
transform -1 0 35144 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1258_
timestamp 1667941163
transform 1 0 34500 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1259_
timestamp 1667941163
transform -1 0 35144 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1260_
timestamp 1667941163
transform 1 0 35328 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1261_
timestamp 1667941163
transform 1 0 35880 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1262_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 35512 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1263_
timestamp 1667941163
transform 1 0 33396 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1264_
timestamp 1667941163
transform 1 0 33304 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1265_
timestamp 1667941163
transform 1 0 24564 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1266_
timestamp 1667941163
transform -1 0 24656 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1267_
timestamp 1667941163
transform -1 0 25484 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1268_
timestamp 1667941163
transform -1 0 23828 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1269_
timestamp 1667941163
transform -1 0 24104 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1270_
timestamp 1667941163
transform 1 0 23736 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1271_
timestamp 1667941163
transform -1 0 23552 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1272_
timestamp 1667941163
transform -1 0 13800 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1273_
timestamp 1667941163
transform -1 0 14996 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1274_
timestamp 1667941163
transform -1 0 14444 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1275_
timestamp 1667941163
transform -1 0 15088 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1276_
timestamp 1667941163
transform -1 0 23552 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1277_
timestamp 1667941163
transform 1 0 21436 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1278_
timestamp 1667941163
transform 1 0 23184 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1279_
timestamp 1667941163
transform -1 0 27784 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1280_
timestamp 1667941163
transform -1 0 27600 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1281_
timestamp 1667941163
transform 1 0 24932 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1282_
timestamp 1667941163
transform 1 0 22540 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_2  _1283_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 23092 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1284_
timestamp 1667941163
transform 1 0 16836 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1285_
timestamp 1667941163
transform 1 0 17756 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1286_
timestamp 1667941163
transform 1 0 21988 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1287_
timestamp 1667941163
transform 1 0 16836 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1288_
timestamp 1667941163
transform 1 0 16652 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1289_
timestamp 1667941163
transform 1 0 17664 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _1290_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 18124 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1291_
timestamp 1667941163
transform -1 0 15364 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1292_
timestamp 1667941163
transform 1 0 16100 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1293_
timestamp 1667941163
transform 1 0 15916 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1294_
timestamp 1667941163
transform -1 0 18584 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1295_
timestamp 1667941163
transform 1 0 15456 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1296_
timestamp 1667941163
transform 1 0 16836 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1297_
timestamp 1667941163
transform -1 0 17112 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1298_
timestamp 1667941163
transform 1 0 16836 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1299_
timestamp 1667941163
transform 1 0 14536 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1300_
timestamp 1667941163
transform 1 0 14720 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1301_
timestamp 1667941163
transform 1 0 15364 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1302_
timestamp 1667941163
transform 1 0 15640 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1303_
timestamp 1667941163
transform -1 0 17664 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1304_
timestamp 1667941163
transform 1 0 19412 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1305_
timestamp 1667941163
transform 1 0 19780 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1306_
timestamp 1667941163
transform -1 0 20148 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _1307_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 21068 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1308_
timestamp 1667941163
transform 1 0 23000 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1309_
timestamp 1667941163
transform -1 0 22908 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1310_
timestamp 1667941163
transform 1 0 23644 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1311_
timestamp 1667941163
transform 1 0 21252 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1312_
timestamp 1667941163
transform 1 0 21068 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1313_
timestamp 1667941163
transform 1 0 21988 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1314_
timestamp 1667941163
transform 1 0 23828 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1315_
timestamp 1667941163
transform -1 0 18952 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1316_
timestamp 1667941163
transform 1 0 18032 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1317_
timestamp 1667941163
transform 1 0 18952 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1318_
timestamp 1667941163
transform -1 0 20240 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1319_
timestamp 1667941163
transform 1 0 21436 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1320_
timestamp 1667941163
transform 1 0 21988 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _1321_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 21988 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1322_
timestamp 1667941163
transform -1 0 21988 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1323_
timestamp 1667941163
transform -1 0 20332 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1324_
timestamp 1667941163
transform 1 0 20700 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1325_
timestamp 1667941163
transform -1 0 21344 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1326_
timestamp 1667941163
transform -1 0 21988 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1327_
timestamp 1667941163
transform -1 0 25392 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1328_
timestamp 1667941163
transform 1 0 25300 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1329_
timestamp 1667941163
transform 1 0 25668 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1330_
timestamp 1667941163
transform 1 0 24564 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1331_
timestamp 1667941163
transform 1 0 22356 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _1332_
timestamp 1667941163
transform -1 0 25116 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1333_
timestamp 1667941163
transform 1 0 23552 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _1334_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 21896 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1335_
timestamp 1667941163
transform 1 0 16928 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1336_
timestamp 1667941163
transform 1 0 18768 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1337_
timestamp 1667941163
transform -1 0 21528 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1338_
timestamp 1667941163
transform -1 0 20792 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1339_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 20240 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1340_
timestamp 1667941163
transform 1 0 20148 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1341_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 20700 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1342_
timestamp 1667941163
transform -1 0 19780 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1343_
timestamp 1667941163
transform 1 0 17112 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1344_
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1345_
timestamp 1667941163
transform -1 0 18216 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1346_
timestamp 1667941163
transform 1 0 18308 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1347_
timestamp 1667941163
transform -1 0 18768 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1348_
timestamp 1667941163
transform 1 0 25484 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1349_
timestamp 1667941163
transform 1 0 17204 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1350_
timestamp 1667941163
transform -1 0 18400 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1351_
timestamp 1667941163
transform -1 0 16376 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1352_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 23736 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1353_
timestamp 1667941163
transform 1 0 17480 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1354_
timestamp 1667941163
transform 1 0 16836 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1355_
timestamp 1667941163
transform 1 0 27140 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1356_
timestamp 1667941163
transform 1 0 27968 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1357_
timestamp 1667941163
transform 1 0 27324 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1358_
timestamp 1667941163
transform -1 0 18952 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1359_
timestamp 1667941163
transform -1 0 21252 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_1  _1360_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 20240 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _1361_
timestamp 1667941163
transform -1 0 22632 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1362_
timestamp 1667941163
transform -1 0 26312 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1363_
timestamp 1667941163
transform -1 0 26680 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1364_
timestamp 1667941163
transform 1 0 25300 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1365_
timestamp 1667941163
transform -1 0 28980 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1366_
timestamp 1667941163
transform -1 0 27692 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1367_
timestamp 1667941163
transform -1 0 27968 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1368_
timestamp 1667941163
transform 1 0 27416 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1369_
timestamp 1667941163
transform -1 0 24104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1370_
timestamp 1667941163
transform 1 0 24748 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1371_
timestamp 1667941163
transform 1 0 25576 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1372_
timestamp 1667941163
transform -1 0 27600 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1373_
timestamp 1667941163
transform -1 0 27508 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1374_
timestamp 1667941163
transform 1 0 26312 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1375_
timestamp 1667941163
transform 1 0 25944 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1376_
timestamp 1667941163
transform -1 0 25668 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1377_
timestamp 1667941163
transform 1 0 27876 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1378_
timestamp 1667941163
transform 1 0 23092 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1379_
timestamp 1667941163
transform 1 0 24748 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1380_
timestamp 1667941163
transform -1 0 25024 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1381_
timestamp 1667941163
transform 1 0 24564 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1382_
timestamp 1667941163
transform 1 0 23644 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1383_
timestamp 1667941163
transform 1 0 21252 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1384_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 26312 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1385_
timestamp 1667941163
transform -1 0 22356 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _1386_
timestamp 1667941163
transform 1 0 24564 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__a31oi_1  _1387_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 20608 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1388_
timestamp 1667941163
transform -1 0 21804 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1389_
timestamp 1667941163
transform -1 0 20056 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1390_
timestamp 1667941163
transform 1 0 19320 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1391_
timestamp 1667941163
transform 1 0 20332 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1392_
timestamp 1667941163
transform -1 0 18584 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1393_
timestamp 1667941163
transform 1 0 19504 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1394_
timestamp 1667941163
transform 1 0 17480 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1395_
timestamp 1667941163
transform 1 0 18216 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1396_
timestamp 1667941163
transform 1 0 18124 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1397_
timestamp 1667941163
transform 1 0 20424 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1398_
timestamp 1667941163
transform -1 0 22540 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1399_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 20332 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1400_
timestamp 1667941163
transform -1 0 25024 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1401_
timestamp 1667941163
transform -1 0 25668 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1402_
timestamp 1667941163
transform 1 0 23644 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1403_
timestamp 1667941163
transform -1 0 22540 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _1404_
timestamp 1667941163
transform 1 0 21988 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1405_
timestamp 1667941163
transform 1 0 24380 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1406_
timestamp 1667941163
transform -1 0 24104 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1407_
timestamp 1667941163
transform 1 0 23276 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1408_
timestamp 1667941163
transform 1 0 23460 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1409_
timestamp 1667941163
transform 1 0 23276 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1410_
timestamp 1667941163
transform -1 0 22724 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1411_
timestamp 1667941163
transform -1 0 24840 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_4  _1412_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 23000 0 1 39168
box -38 -48 1602 592
use sky130_fd_sc_hd__a31oi_1  _1413_
timestamp 1667941163
transform 1 0 15272 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1414_
timestamp 1667941163
transform 1 0 14444 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1415_
timestamp 1667941163
transform -1 0 13800 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1416_
timestamp 1667941163
transform -1 0 12972 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1417_
timestamp 1667941163
transform -1 0 15272 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1418_
timestamp 1667941163
transform 1 0 13616 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1419_
timestamp 1667941163
transform 1 0 12880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1420_
timestamp 1667941163
transform 1 0 14720 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1421_
timestamp 1667941163
transform -1 0 15180 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1422_
timestamp 1667941163
transform 1 0 15732 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1423_
timestamp 1667941163
transform 1 0 15640 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1424_
timestamp 1667941163
transform -1 0 13616 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1425_
timestamp 1667941163
transform -1 0 14536 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1426_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 16008 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _1427_
timestamp 1667941163
transform 1 0 14720 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _1428_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 13892 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1429_
timestamp 1667941163
transform 1 0 24564 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1430_
timestamp 1667941163
transform -1 0 24564 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_8  _1431_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 26680 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _1432_
timestamp 1667941163
transform 1 0 23276 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1433_
timestamp 1667941163
transform 1 0 23276 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1434_
timestamp 1667941163
transform -1 0 25668 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a311oi_1  _1435_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24656 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1436_
timestamp 1667941163
transform 1 0 25392 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1437_
timestamp 1667941163
transform -1 0 24288 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1438_
timestamp 1667941163
transform -1 0 23920 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1439_
timestamp 1667941163
transform 1 0 23184 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1440_
timestamp 1667941163
transform -1 0 23000 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1441_
timestamp 1667941163
transform 1 0 22540 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1442_
timestamp 1667941163
transform 1 0 19136 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1443_
timestamp 1667941163
transform 1 0 20424 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1444_
timestamp 1667941163
transform 1 0 20700 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1445_
timestamp 1667941163
transform 1 0 20424 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1446_
timestamp 1667941163
transform -1 0 20056 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1447_
timestamp 1667941163
transform 1 0 18400 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1448_
timestamp 1667941163
transform 1 0 18032 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1449_
timestamp 1667941163
transform -1 0 18308 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1450_
timestamp 1667941163
transform -1 0 18676 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1451_
timestamp 1667941163
transform 1 0 17388 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1452_
timestamp 1667941163
transform -1 0 17664 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1453_
timestamp 1667941163
transform 1 0 16928 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1454_
timestamp 1667941163
transform 1 0 17296 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1455_
timestamp 1667941163
transform 1 0 15456 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1456_
timestamp 1667941163
transform 1 0 14812 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1457_
timestamp 1667941163
transform 1 0 15916 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_1  _1458_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17848 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1459_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 17388 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1460_
timestamp 1667941163
transform -1 0 18584 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1461_
timestamp 1667941163
transform 1 0 16836 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1462_
timestamp 1667941163
transform 1 0 15824 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1463_
timestamp 1667941163
transform -1 0 17940 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1464_
timestamp 1667941163
transform 1 0 17848 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1465_
timestamp 1667941163
transform 1 0 16836 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1466_
timestamp 1667941163
transform 1 0 15732 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1467_
timestamp 1667941163
transform 1 0 14628 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1468_
timestamp 1667941163
transform -1 0 14352 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1469_
timestamp 1667941163
transform 1 0 16192 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1470_
timestamp 1667941163
transform 1 0 15916 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1471_
timestamp 1667941163
transform 1 0 16100 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1472_
timestamp 1667941163
transform 1 0 16468 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1473_
timestamp 1667941163
transform 1 0 17940 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1474_
timestamp 1667941163
transform -1 0 18584 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1475_
timestamp 1667941163
transform -1 0 17112 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1476_
timestamp 1667941163
transform 1 0 15456 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1477_
timestamp 1667941163
transform 1 0 16100 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1478_
timestamp 1667941163
transform 1 0 14352 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1479_
timestamp 1667941163
transform 1 0 13524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1480_
timestamp 1667941163
transform -1 0 16376 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1481_
timestamp 1667941163
transform 1 0 22724 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1482_
timestamp 1667941163
transform 1 0 23552 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1483_
timestamp 1667941163
transform 1 0 24564 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1484_
timestamp 1667941163
transform 1 0 23092 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1485_
timestamp 1667941163
transform 1 0 23920 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1486_
timestamp 1667941163
transform -1 0 25668 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1487_
timestamp 1667941163
transform -1 0 25484 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1488_
timestamp 1667941163
transform 1 0 20516 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1489_
timestamp 1667941163
transform 1 0 21436 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1490_
timestamp 1667941163
transform -1 0 21896 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1491_
timestamp 1667941163
transform 1 0 20240 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1492_
timestamp 1667941163
transform -1 0 20240 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1493_
timestamp 1667941163
transform 1 0 19688 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1494_
timestamp 1667941163
transform 1 0 20056 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1495_
timestamp 1667941163
transform 1 0 16836 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1496_
timestamp 1667941163
transform 1 0 16836 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1497_
timestamp 1667941163
transform -1 0 21528 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1498_
timestamp 1667941163
transform 1 0 22356 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1499_
timestamp 1667941163
transform 1 0 23000 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1500_
timestamp 1667941163
transform 1 0 19872 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1501_
timestamp 1667941163
transform 1 0 19504 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1502_
timestamp 1667941163
transform -1 0 23460 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1503_
timestamp 1667941163
transform 1 0 23276 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1504_
timestamp 1667941163
transform 1 0 24932 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1505_
timestamp 1667941163
transform 1 0 24564 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1506_
timestamp 1667941163
transform -1 0 24932 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1507_
timestamp 1667941163
transform 1 0 27232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1508_
timestamp 1667941163
transform 1 0 27600 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1509_
timestamp 1667941163
transform 1 0 28244 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1510_
timestamp 1667941163
transform 1 0 28612 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1511_
timestamp 1667941163
transform 1 0 29532 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1512_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 28428 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1513_
timestamp 1667941163
transform 1 0 30360 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1514_
timestamp 1667941163
transform -1 0 28704 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1515_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 30452 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1516_
timestamp 1667941163
transform 1 0 30268 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1517_
timestamp 1667941163
transform 1 0 29716 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1518_
timestamp 1667941163
transform 1 0 29716 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1519_
timestamp 1667941163
transform 1 0 34132 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1520_
timestamp 1667941163
transform 1 0 33856 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1521_
timestamp 1667941163
transform 1 0 32292 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1522_
timestamp 1667941163
transform 1 0 32292 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1523_
timestamp 1667941163
transform 1 0 36156 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1524_
timestamp 1667941163
transform -1 0 33948 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1525_
timestamp 1667941163
transform 1 0 35236 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1526_
timestamp 1667941163
transform -1 0 35052 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1527_
timestamp 1667941163
transform 1 0 27140 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1528_
timestamp 1667941163
transform 1 0 27692 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1529_
timestamp 1667941163
transform -1 0 30820 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1530_
timestamp 1667941163
transform 1 0 31188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1531_
timestamp 1667941163
transform 1 0 33488 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1532_
timestamp 1667941163
transform 1 0 32200 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1533_
timestamp 1667941163
transform 1 0 33120 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1534_
timestamp 1667941163
transform 1 0 33028 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1535_
timestamp 1667941163
transform 1 0 29992 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1536_
timestamp 1667941163
transform 1 0 29716 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1537_
timestamp 1667941163
transform 1 0 29716 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1538_
timestamp 1667941163
transform 1 0 28704 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1539_
timestamp 1667941163
transform 1 0 29716 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1540_
timestamp 1667941163
transform -1 0 29256 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1541_
timestamp 1667941163
transform 1 0 30176 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1542_
timestamp 1667941163
transform 1 0 28704 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1543_
timestamp 1667941163
transform -1 0 30452 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1544_
timestamp 1667941163
transform -1 0 31372 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1545_
timestamp 1667941163
transform 1 0 28428 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1546_
timestamp 1667941163
transform 1 0 28152 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1547_
timestamp 1667941163
transform 1 0 30176 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1548_
timestamp 1667941163
transform -1 0 30452 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  _1549_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6072 0 1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_2  _1550_
timestamp 1667941163
transform 1 0 9568 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1551_
timestamp 1667941163
transform 1 0 9016 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1552_
timestamp 1667941163
transform -1 0 9476 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1553_
timestamp 1667941163
transform -1 0 8372 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1554_
timestamp 1667941163
transform 1 0 8004 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1555_
timestamp 1667941163
transform 1 0 8280 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1556_
timestamp 1667941163
transform 1 0 7360 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1557_
timestamp 1667941163
transform 1 0 6256 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1558_
timestamp 1667941163
transform -1 0 5428 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1559_
timestamp 1667941163
transform -1 0 6900 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1560_
timestamp 1667941163
transform -1 0 8096 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1561_
timestamp 1667941163
transform -1 0 9844 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1562_
timestamp 1667941163
transform -1 0 4600 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1563_
timestamp 1667941163
transform -1 0 4692 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1564_
timestamp 1667941163
transform -1 0 4600 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1565_
timestamp 1667941163
transform 1 0 4600 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1566_
timestamp 1667941163
transform -1 0 6808 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1567_
timestamp 1667941163
transform -1 0 8740 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1568_
timestamp 1667941163
transform 1 0 8096 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1569_
timestamp 1667941163
transform 1 0 36064 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1570_
timestamp 1667941163
transform 1 0 37444 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1571_
timestamp 1667941163
transform -1 0 37812 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _1572_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 35972 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1573_
timestamp 1667941163
transform 1 0 37444 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1574_
timestamp 1667941163
transform -1 0 35972 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1575_
timestamp 1667941163
transform 1 0 42320 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1576_
timestamp 1667941163
transform 1 0 40296 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1577_
timestamp 1667941163
transform 1 0 42688 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1578_
timestamp 1667941163
transform 1 0 44804 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1579_
timestamp 1667941163
transform 1 0 43240 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1580_
timestamp 1667941163
transform 1 0 43700 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1581_
timestamp 1667941163
transform 1 0 44068 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1582_
timestamp 1667941163
transform 1 0 45080 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1583_
timestamp 1667941163
transform -1 0 45540 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1584_
timestamp 1667941163
transform 1 0 45080 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1585_
timestamp 1667941163
transform 1 0 46092 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1586_
timestamp 1667941163
transform -1 0 44620 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1587_
timestamp 1667941163
transform 1 0 45172 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1588_
timestamp 1667941163
transform -1 0 45080 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1589_
timestamp 1667941163
transform -1 0 44620 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1590_
timestamp 1667941163
transform -1 0 43792 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1591_
timestamp 1667941163
transform 1 0 43700 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1592_
timestamp 1667941163
transform -1 0 45540 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1593_
timestamp 1667941163
transform 1 0 45172 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1594_
timestamp 1667941163
transform -1 0 44712 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1595_
timestamp 1667941163
transform 1 0 44068 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1596_
timestamp 1667941163
transform 1 0 44068 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1597_
timestamp 1667941163
transform 1 0 43700 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o41a_1  _1598_
timestamp 1667941163
transform 1 0 43424 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1599_
timestamp 1667941163
transform -1 0 43700 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1600_
timestamp 1667941163
transform -1 0 44436 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1601_
timestamp 1667941163
transform -1 0 43516 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1602_
timestamp 1667941163
transform 1 0 39836 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1603_
timestamp 1667941163
transform 1 0 40848 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _1604_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 42596 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _1605_
timestamp 1667941163
transform 1 0 40020 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1606_
timestamp 1667941163
transform -1 0 41768 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1607_
timestamp 1667941163
transform -1 0 40388 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1608_
timestamp 1667941163
transform 1 0 40112 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1609_
timestamp 1667941163
transform -1 0 41124 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1610_
timestamp 1667941163
transform 1 0 40388 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1611_
timestamp 1667941163
transform 1 0 42044 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1612_
timestamp 1667941163
transform -1 0 42044 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1613_
timestamp 1667941163
transform -1 0 41400 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1614_
timestamp 1667941163
transform 1 0 40020 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1615_
timestamp 1667941163
transform 1 0 40020 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1616_
timestamp 1667941163
transform -1 0 39560 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1617_
timestamp 1667941163
transform 1 0 39560 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _1618_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 42136 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _1619_
timestamp 1667941163
transform -1 0 39560 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1620_
timestamp 1667941163
transform 1 0 41124 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1621_
timestamp 1667941163
transform 1 0 40020 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1622_
timestamp 1667941163
transform -1 0 41216 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1623_
timestamp 1667941163
transform 1 0 41216 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _1624_
timestamp 1667941163
transform 1 0 41124 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _1625_
timestamp 1667941163
transform 1 0 40940 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1626_
timestamp 1667941163
transform -1 0 42596 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1627_
timestamp 1667941163
transform 1 0 41676 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1628_
timestamp 1667941163
transform 1 0 43700 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1629_
timestamp 1667941163
transform 1 0 43148 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1630_
timestamp 1667941163
transform -1 0 44436 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1631_
timestamp 1667941163
transform -1 0 43056 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1632_
timestamp 1667941163
transform 1 0 42596 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1633_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 42320 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1634_
timestamp 1667941163
transform 1 0 43148 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1635_
timestamp 1667941163
transform 1 0 42044 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _1636_
timestamp 1667941163
transform -1 0 42136 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _1637_
timestamp 1667941163
transform -1 0 43516 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1638_
timestamp 1667941163
transform -1 0 43608 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1639_
timestamp 1667941163
transform 1 0 43976 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1640_
timestamp 1667941163
transform -1 0 44528 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1641_
timestamp 1667941163
transform -1 0 45632 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1642_
timestamp 1667941163
transform 1 0 43792 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1643_
timestamp 1667941163
transform -1 0 44252 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1644_
timestamp 1667941163
transform -1 0 44344 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_1  _1645_
timestamp 1667941163
transform -1 0 43332 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1646_
timestamp 1667941163
transform -1 0 43792 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1647_
timestamp 1667941163
transform 1 0 43700 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1648_
timestamp 1667941163
transform -1 0 44988 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1649_
timestamp 1667941163
transform -1 0 44620 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1650_
timestamp 1667941163
transform 1 0 43056 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1651_
timestamp 1667941163
transform -1 0 42688 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1652_
timestamp 1667941163
transform -1 0 44712 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1653_
timestamp 1667941163
transform -1 0 44160 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _1654_
timestamp 1667941163
transform -1 0 43792 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1655_
timestamp 1667941163
transform 1 0 43884 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1656_
timestamp 1667941163
transform 1 0 43884 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _1657_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 42780 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1658_
timestamp 1667941163
transform 1 0 42136 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1659_
timestamp 1667941163
transform -1 0 26588 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1660_
timestamp 1667941163
transform -1 0 19964 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1661_
timestamp 1667941163
transform 1 0 16836 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1662_
timestamp 1667941163
transform -1 0 15916 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1663_
timestamp 1667941163
transform 1 0 15364 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1664_
timestamp 1667941163
transform -1 0 25668 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1665_
timestamp 1667941163
transform 1 0 17020 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1666_
timestamp 1667941163
transform 1 0 15456 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1667_
timestamp 1667941163
transform 1 0 15640 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1668_
timestamp 1667941163
transform 1 0 17480 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1669_
timestamp 1667941163
transform 1 0 16928 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1670_
timestamp 1667941163
transform 1 0 17848 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1671_
timestamp 1667941163
transform 1 0 14996 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1672_
timestamp 1667941163
transform -1 0 14812 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1673_
timestamp 1667941163
transform 1 0 13524 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1674_
timestamp 1667941163
transform 1 0 12144 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1675_
timestamp 1667941163
transform 1 0 11776 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1676_
timestamp 1667941163
transform -1 0 12328 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1677_
timestamp 1667941163
transform 1 0 14260 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1678_
timestamp 1667941163
transform -1 0 13800 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1679_
timestamp 1667941163
transform -1 0 14536 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1680_
timestamp 1667941163
transform -1 0 13064 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1681_
timestamp 1667941163
transform 1 0 13524 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1682_
timestamp 1667941163
transform -1 0 11868 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1683_
timestamp 1667941163
transform 1 0 11684 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1684_
timestamp 1667941163
transform -1 0 11960 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1685_
timestamp 1667941163
transform -1 0 11224 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1686_
timestamp 1667941163
transform 1 0 12236 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1687_
timestamp 1667941163
transform -1 0 11868 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1688_
timestamp 1667941163
transform 1 0 12052 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1689_
timestamp 1667941163
transform 1 0 12144 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1690_
timestamp 1667941163
transform 1 0 11776 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1691_
timestamp 1667941163
transform -1 0 12972 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1692_
timestamp 1667941163
transform 1 0 26404 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1693_
timestamp 1667941163
transform -1 0 27232 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _1694_
timestamp 1667941163
transform -1 0 27048 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1695_
timestamp 1667941163
transform 1 0 26312 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1696_
timestamp 1667941163
transform 1 0 25208 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1697_
timestamp 1667941163
transform 1 0 27140 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1698_
timestamp 1667941163
transform -1 0 26496 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1699_
timestamp 1667941163
transform -1 0 29072 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1700_
timestamp 1667941163
transform 1 0 30728 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1701_
timestamp 1667941163
transform -1 0 29532 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1702_
timestamp 1667941163
transform 1 0 28888 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1703_
timestamp 1667941163
transform -1 0 30728 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1704_
timestamp 1667941163
transform 1 0 27508 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1705_
timestamp 1667941163
transform 1 0 28612 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1706_
timestamp 1667941163
transform 1 0 31372 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1707_
timestamp 1667941163
transform 1 0 31464 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1708_
timestamp 1667941163
transform 1 0 30268 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1709_
timestamp 1667941163
transform 1 0 29348 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1710_
timestamp 1667941163
transform -1 0 30636 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1711_
timestamp 1667941163
transform 1 0 29900 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1712_
timestamp 1667941163
transform 1 0 37628 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1713_
timestamp 1667941163
transform -1 0 36984 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1714_
timestamp 1667941163
transform -1 0 32660 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1715_
timestamp 1667941163
transform 1 0 33028 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1716_
timestamp 1667941163
transform -1 0 39468 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1717_
timestamp 1667941163
transform 1 0 38732 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1718_
timestamp 1667941163
transform -1 0 40572 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1719_
timestamp 1667941163
transform 1 0 40020 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1720_
timestamp 1667941163
transform 1 0 38824 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1721_
timestamp 1667941163
transform -1 0 39284 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1722_
timestamp 1667941163
transform -1 0 33120 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1723_
timestamp 1667941163
transform 1 0 32660 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1724_
timestamp 1667941163
transform -1 0 34316 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1725_
timestamp 1667941163
transform 1 0 34868 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1726_
timestamp 1667941163
transform -1 0 31004 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1727_
timestamp 1667941163
transform 1 0 31096 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1728_
timestamp 1667941163
transform 1 0 28520 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1729_
timestamp 1667941163
transform -1 0 31004 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1730_
timestamp 1667941163
transform 1 0 30452 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1731_
timestamp 1667941163
transform -1 0 30452 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1732_
timestamp 1667941163
transform 1 0 30912 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1733_
timestamp 1667941163
transform -1 0 31280 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1734_
timestamp 1667941163
transform 1 0 31280 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1735_
timestamp 1667941163
transform -1 0 30636 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1736_
timestamp 1667941163
transform 1 0 33120 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1737_
timestamp 1667941163
transform -1 0 29256 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1738_
timestamp 1667941163
transform 1 0 29532 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1739_
timestamp 1667941163
transform -1 0 31372 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1740_
timestamp 1667941163
transform 1 0 32292 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1741_
timestamp 1667941163
transform 1 0 39008 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1742_
timestamp 1667941163
transform -1 0 27784 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1743_
timestamp 1667941163
transform -1 0 26680 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1744_
timestamp 1667941163
transform 1 0 25852 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _1745_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 27692 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1746_
timestamp 1667941163
transform 1 0 26128 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1747_
timestamp 1667941163
transform 1 0 25300 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1748_
timestamp 1667941163
transform 1 0 25208 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1749_
timestamp 1667941163
transform -1 0 27876 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1750_
timestamp 1667941163
transform 1 0 27140 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1751_
timestamp 1667941163
transform 1 0 24564 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1752_
timestamp 1667941163
transform 1 0 24564 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1753_
timestamp 1667941163
transform 1 0 24564 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1754_
timestamp 1667941163
transform 1 0 23368 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1755_
timestamp 1667941163
transform 1 0 25668 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1756_
timestamp 1667941163
transform 1 0 14536 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1757_
timestamp 1667941163
transform 1 0 14260 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1758_
timestamp 1667941163
transform 1 0 14352 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1759_
timestamp 1667941163
transform 1 0 14260 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1760_
timestamp 1667941163
transform 1 0 14260 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1761_
timestamp 1667941163
transform 1 0 14260 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1762_
timestamp 1667941163
transform 1 0 12788 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1763_
timestamp 1667941163
transform 1 0 12328 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1764_
timestamp 1667941163
transform 1 0 13064 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1765_
timestamp 1667941163
transform 1 0 12144 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1766_
timestamp 1667941163
transform 1 0 14260 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1767_
timestamp 1667941163
transform -1 0 11868 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1768_
timestamp 1667941163
transform -1 0 26404 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1769_
timestamp 1667941163
transform 1 0 27140 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1770_
timestamp 1667941163
transform 1 0 25760 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1771_
timestamp 1667941163
transform 1 0 25944 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1772_
timestamp 1667941163
transform 1 0 18124 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1773_
timestamp 1667941163
transform 1 0 17848 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1774_
timestamp 1667941163
transform 1 0 18032 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1775_
timestamp 1667941163
transform 1 0 17020 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1776_
timestamp 1667941163
transform 1 0 25392 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1777_
timestamp 1667941163
transform 1 0 18216 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1778_
timestamp 1667941163
transform 1 0 17756 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1779_
timestamp 1667941163
transform 1 0 26220 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1780_
timestamp 1667941163
transform -1 0 26956 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1781_
timestamp 1667941163
transform -1 0 26680 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1782_
timestamp 1667941163
transform 1 0 27048 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1783_
timestamp 1667941163
transform 1 0 27876 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1784_
timestamp 1667941163
transform 1 0 21988 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1785_
timestamp 1667941163
transform 1 0 22632 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1786_
timestamp 1667941163
transform 1 0 22172 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1787_
timestamp 1667941163
transform 1 0 21988 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1788_
timestamp 1667941163
transform 1 0 21988 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1789_
timestamp 1667941163
transform -1 0 23644 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1790_
timestamp 1667941163
transform 1 0 24104 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1791_
timestamp 1667941163
transform 1 0 20332 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1792_
timestamp 1667941163
transform 1 0 20056 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1793_
timestamp 1667941163
transform -1 0 20148 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1794_
timestamp 1667941163
transform 1 0 19412 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1795_
timestamp 1667941163
transform 1 0 19596 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1796_
timestamp 1667941163
transform 1 0 19504 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1797_
timestamp 1667941163
transform -1 0 20148 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1798_
timestamp 1667941163
transform 1 0 20792 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1799_
timestamp 1667941163
transform 1 0 19688 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1800_
timestamp 1667941163
transform 1 0 19596 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1801_
timestamp 1667941163
transform -1 0 22540 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1802_
timestamp 1667941163
transform 1 0 21988 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1803_
timestamp 1667941163
transform 1 0 19964 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1804_
timestamp 1667941163
transform -1 0 19780 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1805_
timestamp 1667941163
transform -1 0 27876 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1806_
timestamp 1667941163
transform 1 0 28244 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1807_
timestamp 1667941163
transform 1 0 27140 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1808_
timestamp 1667941163
transform 1 0 26128 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1809_
timestamp 1667941163
transform 1 0 20792 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1810_
timestamp 1667941163
transform -1 0 19964 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1811_
timestamp 1667941163
transform 1 0 20976 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1812_
timestamp 1667941163
transform 1 0 20884 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1813_
timestamp 1667941163
transform 1 0 23276 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1814_
timestamp 1667941163
transform 1 0 23184 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1815_
timestamp 1667941163
transform -1 0 26772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1816_
timestamp 1667941163
transform 1 0 26128 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1817_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 28336 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1818_
timestamp 1667941163
transform -1 0 32660 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1819_
timestamp 1667941163
transform 1 0 35328 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1820_
timestamp 1667941163
transform 1 0 32384 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1821_
timestamp 1667941163
transform 1 0 37996 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1822_
timestamp 1667941163
transform 1 0 40020 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1823_
timestamp 1667941163
transform -1 0 41492 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1824_
timestamp 1667941163
transform 1 0 34868 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1825_
timestamp 1667941163
transform 1 0 36064 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1826_
timestamp 1667941163
transform 1 0 32752 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1827_
timestamp 1667941163
transform 1 0 31648 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1828_
timestamp 1667941163
transform -1 0 38916 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1829_
timestamp 1667941163
transform 1 0 34132 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1830_
timestamp 1667941163
transform 1 0 32292 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1831_
timestamp 1667941163
transform -1 0 39100 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1832_
timestamp 1667941163
transform 1 0 33120 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1833_
timestamp 1667941163
transform 1 0 21988 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1834_
timestamp 1667941163
transform -1 0 20884 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1835_
timestamp 1667941163
transform 1 0 15364 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1836_
timestamp 1667941163
transform 1 0 15640 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1837_
timestamp 1667941163
transform 1 0 24932 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1838_
timestamp 1667941163
transform 1 0 27692 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1839_
timestamp 1667941163
transform -1 0 27508 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1840_
timestamp 1667941163
transform -1 0 24012 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1841_
timestamp 1667941163
transform -1 0 22080 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1842_
timestamp 1667941163
transform 1 0 17480 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1843_
timestamp 1667941163
transform 1 0 24564 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1844_
timestamp 1667941163
transform 1 0 23092 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1845_
timestamp 1667941163
transform 1 0 12880 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1846_
timestamp 1667941163
transform 1 0 12144 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1847_
timestamp 1667941163
transform 1 0 15548 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1848_
timestamp 1667941163
transform -1 0 14352 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1849_
timestamp 1667941163
transform 1 0 23000 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1850_
timestamp 1667941163
transform 1 0 25944 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1851_
timestamp 1667941163
transform 1 0 21988 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1852_
timestamp 1667941163
transform 1 0 20056 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1853_
timestamp 1667941163
transform 1 0 16836 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1854_
timestamp 1667941163
transform 1 0 14352 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1855_
timestamp 1667941163
transform 1 0 16100 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1856_
timestamp 1667941163
transform 1 0 14260 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1857_
timestamp 1667941163
transform -1 0 18584 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1858_
timestamp 1667941163
transform 1 0 13156 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1859_
timestamp 1667941163
transform 1 0 23368 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1860_
timestamp 1667941163
transform 1 0 24012 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1861_
timestamp 1667941163
transform -1 0 20884 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1862_
timestamp 1667941163
transform 1 0 15916 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1863_
timestamp 1667941163
transform 1 0 19136 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1864_
timestamp 1667941163
transform -1 0 26036 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1865_
timestamp 1667941163
transform 1 0 28428 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1866_
timestamp 1667941163
transform 1 0 28796 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1867_
timestamp 1667941163
transform 1 0 33672 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1868_
timestamp 1667941163
transform 1 0 31464 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1869_
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1870_
timestamp 1667941163
transform 1 0 35052 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1871_
timestamp 1667941163
transform -1 0 31004 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1872_
timestamp 1667941163
transform 1 0 32016 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1873_
timestamp 1667941163
transform 1 0 32844 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1874_
timestamp 1667941163
transform 1 0 29532 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1875_
timestamp 1667941163
transform 1 0 28428 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1876_
timestamp 1667941163
transform 1 0 28704 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1877_
timestamp 1667941163
transform 1 0 28336 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1878_
timestamp 1667941163
transform 1 0 28704 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1879_
timestamp 1667941163
transform 1 0 27692 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1880_
timestamp 1667941163
transform 1 0 29992 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1881_
timestamp 1667941163
transform 1 0 12328 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1882_
timestamp 1667941163
transform 1 0 10488 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1883_
timestamp 1667941163
transform 1 0 9384 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1884_
timestamp 1667941163
transform 1 0 8924 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1885_
timestamp 1667941163
transform 1 0 8096 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1886_
timestamp 1667941163
transform 1 0 8740 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1887_
timestamp 1667941163
transform 1 0 9108 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1888_
timestamp 1667941163
transform 1 0 8096 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1889_
timestamp 1667941163
transform 1 0 6532 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1890_
timestamp 1667941163
transform 1 0 5796 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1891_
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1892_
timestamp 1667941163
transform 1 0 7360 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1893_
timestamp 1667941163
transform 1 0 9384 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1894_
timestamp 1667941163
transform 1 0 4140 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1895_
timestamp 1667941163
transform 1 0 4324 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1896_
timestamp 1667941163
transform 1 0 4232 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1897_
timestamp 1667941163
transform 1 0 4784 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1898_
timestamp 1667941163
transform 1 0 6532 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1899_
timestamp 1667941163
transform 1 0 7820 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1900_
timestamp 1667941163
transform -1 0 9660 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1901_
timestamp 1667941163
transform 1 0 43240 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1902_
timestamp 1667941163
transform 1 0 46092 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1903_
timestamp 1667941163
transform 1 0 44620 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1904_
timestamp 1667941163
transform 1 0 43240 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1905_
timestamp 1667941163
transform 1 0 38088 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1906_
timestamp 1667941163
transform 1 0 40204 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1907_
timestamp 1667941163
transform 1 0 37720 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1908_
timestamp 1667941163
transform 1 0 39100 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1909_
timestamp 1667941163
transform -1 0 42780 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1910_
timestamp 1667941163
transform 1 0 41308 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1911_
timestamp 1667941163
transform 1 0 44252 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1912_
timestamp 1667941163
transform 1 0 43884 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1913_
timestamp 1667941163
transform 1 0 45172 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1914_
timestamp 1667941163
transform 1 0 42872 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1915_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 44620 0 -1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1916_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 41492 0 1 27200
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1917_
timestamp 1667941163
transform 1 0 14996 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1918_
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1919_
timestamp 1667941163
transform -1 0 18032 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1920_
timestamp 1667941163
transform 1 0 13156 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1921_
timestamp 1667941163
transform -1 0 13156 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1922_
timestamp 1667941163
transform -1 0 14812 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1923_
timestamp 1667941163
transform 1 0 11684 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1924_
timestamp 1667941163
transform -1 0 13156 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1925_
timestamp 1667941163
transform 1 0 11684 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1926_
timestamp 1667941163
transform -1 0 13248 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1927_
timestamp 1667941163
transform 1 0 25760 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1928_
timestamp 1667941163
transform -1 0 29992 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1929_
timestamp 1667941163
transform 1 0 29808 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1930_
timestamp 1667941163
transform 1 0 29716 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1931_
timestamp 1667941163
transform 1 0 36892 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1932_
timestamp 1667941163
transform 1 0 32292 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1933_
timestamp 1667941163
transform 1 0 38272 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1934_
timestamp 1667941163
transform 1 0 40020 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1935_
timestamp 1667941163
transform -1 0 39560 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1936_
timestamp 1667941163
transform 1 0 32292 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1937_
timestamp 1667941163
transform 1 0 34224 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1938_
timestamp 1667941163
transform 1 0 30912 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1939_
timestamp 1667941163
transform 1 0 30176 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1940_
timestamp 1667941163
transform -1 0 33304 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1941_
timestamp 1667941163
transform 1 0 32292 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1942_
timestamp 1667941163
transform 1 0 31280 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1943_
timestamp 1667941163
transform 1 0 29716 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1944_
timestamp 1667941163
transform 1 0 31648 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1945_
timestamp 1667941163
transform 1 0 38916 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1946_
timestamp 1667941163
transform 1 0 24840 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1947_
timestamp 1667941163
transform 1 0 26772 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1948_
timestamp 1667941163
transform 1 0 24104 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1949_
timestamp 1667941163
transform 1 0 22908 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1950_
timestamp 1667941163
transform 1 0 14076 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1951_
timestamp 1667941163
transform 1 0 13984 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1952_
timestamp 1667941163
transform 1 0 13248 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1953_
timestamp 1667941163
transform 1 0 11868 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1954_
timestamp 1667941163
transform 1 0 12236 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1955_
timestamp 1667941163
transform 1 0 11868 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1956_
timestamp 1667941163
transform -1 0 26680 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1957_
timestamp 1667941163
transform -1 0 26956 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1958_
timestamp 1667941163
transform 1 0 17480 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1959_
timestamp 1667941163
transform 1 0 16192 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1960_
timestamp 1667941163
transform 1 0 17296 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1961_
timestamp 1667941163
transform -1 0 28612 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1962_
timestamp 1667941163
transform 1 0 27140 0 -1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1963_
timestamp 1667941163
transform 1 0 21988 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1964_
timestamp 1667941163
transform 1 0 21252 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1965_
timestamp 1667941163
transform -1 0 23736 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1966_
timestamp 1667941163
transform 1 0 19780 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1967_
timestamp 1667941163
transform -1 0 19412 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1968_
timestamp 1667941163
transform 1 0 19228 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1969_
timestamp 1667941163
transform -1 0 20424 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1970_
timestamp 1667941163
transform 1 0 19228 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1971_
timestamp 1667941163
transform -1 0 22908 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1972_
timestamp 1667941163
transform 1 0 19412 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1973_
timestamp 1667941163
transform -1 0 27876 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1974_
timestamp 1667941163
transform 1 0 26036 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1975_
timestamp 1667941163
transform 1 0 20332 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1976_
timestamp 1667941163
transform 1 0 20056 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1977_
timestamp 1667941163
transform 1 0 22632 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1978_
timestamp 1667941163
transform -1 0 26680 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _2076__26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 8464 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2076_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 7452 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2077__27
timestamp 1667941163
transform 1 0 1748 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2077_
timestamp 1667941163
transform 1 0 2024 0 -1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2078__28
timestamp 1667941163
transform -1 0 20332 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2078_
timestamp 1667941163
transform 1 0 19596 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2079_
timestamp 1667941163
transform 1 0 2024 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2079__29
timestamp 1667941163
transform -1 0 2392 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2080__30
timestamp 1667941163
transform 1 0 45816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2080_
timestamp 1667941163
transform -1 0 46828 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2081__31
timestamp 1667941163
transform 1 0 2852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2081_
timestamp 1667941163
transform -1 0 3772 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2082__32
timestamp 1667941163
transform -1 0 47104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2082_
timestamp 1667941163
transform 1 0 46460 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2083_
timestamp 1667941163
transform 1 0 6716 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2084_
timestamp 1667941163
transform 1 0 45816 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2085_
timestamp 1667941163
transform 1 0 45356 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2086_
timestamp 1667941163
transform 1 0 46460 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2087_
timestamp 1667941163
transform 1 0 21804 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2088_
timestamp 1667941163
transform 1 0 15824 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2089_
timestamp 1667941163
transform -1 0 14904 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2090_
timestamp 1667941163
transform 1 0 17572 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2091_
timestamp 1667941163
transform -1 0 7176 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2092__33
timestamp 1667941163
transform -1 0 47288 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2092_
timestamp 1667941163
transform 1 0 46460 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2093__34
timestamp 1667941163
transform 1 0 47748 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2093_
timestamp 1667941163
transform -1 0 48392 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2094__35
timestamp 1667941163
transform 1 0 6532 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2094_
timestamp 1667941163
transform -1 0 7360 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2095_
timestamp 1667941163
transform -1 0 47288 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2095__36
timestamp 1667941163
transform 1 0 47012 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2096__37
timestamp 1667941163
transform 1 0 2116 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2096_
timestamp 1667941163
transform -1 0 3496 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2097__38
timestamp 1667941163
transform -1 0 47288 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2097_
timestamp 1667941163
transform 1 0 46460 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2098__39
timestamp 1667941163
transform -1 0 30084 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2098_
timestamp 1667941163
transform 1 0 29716 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2099_
timestamp 1667941163
transform 1 0 11868 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2099__40
timestamp 1667941163
transform -1 0 12696 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2100__41
timestamp 1667941163
transform -1 0 48024 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2100_
timestamp 1667941163
transform 1 0 46460 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2101__42
timestamp 1667941163
transform -1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2101_
timestamp 1667941163
transform -1 0 3496 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2102__43
timestamp 1667941163
transform 1 0 47748 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2102_
timestamp 1667941163
transform -1 0 48392 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2103__44
timestamp 1667941163
transform -1 0 6808 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2103_
timestamp 1667941163
transform -1 0 4048 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2104__45
timestamp 1667941163
transform 1 0 44344 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2104_
timestamp 1667941163
transform 1 0 45172 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2105__46
timestamp 1667941163
transform 1 0 5244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2105_
timestamp 1667941163
transform 1 0 5888 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2106__47
timestamp 1667941163
transform -1 0 47288 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2106_
timestamp 1667941163
transform 1 0 46460 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2107_
timestamp 1667941163
transform -1 0 47288 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2107__48
timestamp 1667941163
transform 1 0 47012 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2108__49
timestamp 1667941163
transform -1 0 39192 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2108_
timestamp 1667941163
transform 1 0 38916 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2109__50
timestamp 1667941163
transform -1 0 33396 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2109_
timestamp 1667941163
transform 1 0 33028 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2110__51
timestamp 1667941163
transform -1 0 6900 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2110_
timestamp 1667941163
transform 1 0 6624 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2111__52
timestamp 1667941163
transform 1 0 1748 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2111_
timestamp 1667941163
transform 1 0 2024 0 -1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2112__53
timestamp 1667941163
transform -1 0 47288 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2112_
timestamp 1667941163
transform 1 0 46460 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2113__54
timestamp 1667941163
transform -1 0 22816 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2113_
timestamp 1667941163
transform 1 0 22448 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2114_
timestamp 1667941163
transform 1 0 46460 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2114__55
timestamp 1667941163
transform 1 0 45172 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2115__56
timestamp 1667941163
transform -1 0 2392 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2115_
timestamp 1667941163
transform 1 0 2024 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2116__57
timestamp 1667941163
transform 1 0 18676 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2116_
timestamp 1667941163
transform 1 0 19412 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2117__58
timestamp 1667941163
transform 1 0 4508 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2117_
timestamp 1667941163
transform -1 0 6072 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2118__59
timestamp 1667941163
transform 1 0 47748 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2118_
timestamp 1667941163
transform -1 0 48392 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2119__60
timestamp 1667941163
transform 1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2119_
timestamp 1667941163
transform -1 0 3496 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2120_
timestamp 1667941163
transform -1 0 3496 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2120__61
timestamp 1667941163
transform 1 0 2116 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2121__62
timestamp 1667941163
transform -1 0 39284 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2121_
timestamp 1667941163
transform 1 0 39008 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2122__63
timestamp 1667941163
transform -1 0 48024 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2122_
timestamp 1667941163
transform 1 0 46460 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2123__64
timestamp 1667941163
transform 1 0 5428 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2123_
timestamp 1667941163
transform -1 0 7360 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2124__65
timestamp 1667941163
transform 1 0 47748 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2124_
timestamp 1667941163
transform -1 0 48392 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2125_
timestamp 1667941163
transform 1 0 45356 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2125__66
timestamp 1667941163
transform -1 0 46184 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2126__67
timestamp 1667941163
transform -1 0 46460 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2126_
timestamp 1667941163
transform 1 0 46092 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2127_
timestamp 1667941163
transform -1 0 8280 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2128__68
timestamp 1667941163
transform -1 0 40388 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2128_
timestamp 1667941163
transform 1 0 40112 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2129_
timestamp 1667941163
transform 1 0 6532 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2130_
timestamp 1667941163
transform 1 0 31832 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2130__69
timestamp 1667941163
transform 1 0 31188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2131__70
timestamp 1667941163
transform 1 0 47748 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2131_
timestamp 1667941163
transform -1 0 48392 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2132__71
timestamp 1667941163
transform -1 0 28336 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2132_
timestamp 1667941163
transform 1 0 27140 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2133_
timestamp 1667941163
transform 1 0 37444 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2133__72
timestamp 1667941163
transform 1 0 36064 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2134_
timestamp 1667941163
transform -1 0 3496 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2134__73
timestamp 1667941163
transform 1 0 2944 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2135__74
timestamp 1667941163
transform 1 0 38088 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2135_
timestamp 1667941163
transform 1 0 39744 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2136__75
timestamp 1667941163
transform 1 0 16744 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2136_
timestamp 1667941163
transform 1 0 16836 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2137__76
timestamp 1667941163
transform 1 0 43700 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2137_
timestamp 1667941163
transform 1 0 44896 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2138__77
timestamp 1667941163
transform -1 0 3680 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2138_
timestamp 1667941163
transform -1 0 3496 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2139__78
timestamp 1667941163
transform 1 0 2116 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2139_
timestamp 1667941163
transform -1 0 3496 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2140__79
timestamp 1667941163
transform -1 0 6808 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2140_
timestamp 1667941163
transform -1 0 3496 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2141__80
timestamp 1667941163
transform -1 0 43516 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2141_
timestamp 1667941163
transform 1 0 42780 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2142__81
timestamp 1667941163
transform -1 0 48024 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2142_
timestamp 1667941163
transform 1 0 46460 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2143__82
timestamp 1667941163
transform 1 0 47472 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2143_
timestamp 1667941163
transform -1 0 48392 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2144__83
timestamp 1667941163
transform -1 0 17112 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2144_
timestamp 1667941163
transform -1 0 16928 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2145__84
timestamp 1667941163
transform 1 0 47748 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2145_
timestamp 1667941163
transform -1 0 48392 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2146_
timestamp 1667941163
transform 1 0 25760 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2146__85
timestamp 1667941163
transform 1 0 25116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2147__86
timestamp 1667941163
transform -1 0 39008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2147_
timestamp 1667941163
transform 1 0 38732 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2148__87
timestamp 1667941163
transform 1 0 41308 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2148_
timestamp 1667941163
transform 1 0 42596 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2149__88
timestamp 1667941163
transform -1 0 25576 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2149_
timestamp 1667941163
transform 1 0 24748 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2150_
timestamp 1667941163
transform -1 0 47288 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2150__89
timestamp 1667941163
transform -1 0 48024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2151__90
timestamp 1667941163
transform -1 0 4232 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2151_
timestamp 1667941163
transform 1 0 3772 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2152__91
timestamp 1667941163
transform 1 0 47748 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2152_
timestamp 1667941163
transform -1 0 48392 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2153__92
timestamp 1667941163
transform -1 0 12696 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2153_
timestamp 1667941163
transform 1 0 12052 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2154__93
timestamp 1667941163
transform 1 0 3956 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2154_
timestamp 1667941163
transform 1 0 4048 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2155_
timestamp 1667941163
transform 1 0 10488 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2155__94
timestamp 1667941163
transform -1 0 10764 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2156_
timestamp 1667941163
transform 1 0 2024 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2156__95
timestamp 1667941163
transform -1 0 2392 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2157__96
timestamp 1667941163
transform 1 0 46368 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2157_
timestamp 1667941163
transform 1 0 46460 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2158__97
timestamp 1667941163
transform 1 0 47472 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2158_
timestamp 1667941163
transform -1 0 48392 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2159__98
timestamp 1667941163
transform 1 0 47748 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2159_
timestamp 1667941163
transform -1 0 48392 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2160_
timestamp 1667941163
transform -1 0 4048 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2160__99
timestamp 1667941163
transform 1 0 2300 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2161__100
timestamp 1667941163
transform 1 0 13524 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2161_
timestamp 1667941163
transform 1 0 14260 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2162__101
timestamp 1667941163
transform -1 0 48392 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2162_
timestamp 1667941163
transform -1 0 44528 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2163__102
timestamp 1667941163
transform -1 0 13432 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2163_
timestamp 1667941163
transform 1 0 13156 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2164__103
timestamp 1667941163
transform -1 0 35696 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2164_
timestamp 1667941163
transform 1 0 35328 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2165_
timestamp 1667941163
transform 1 0 14352 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2165__104
timestamp 1667941163
transform -1 0 14720 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2166__105
timestamp 1667941163
transform -1 0 47288 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2166_
timestamp 1667941163
transform 1 0 46460 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2167__106
timestamp 1667941163
transform 1 0 4876 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2167_
timestamp 1667941163
transform -1 0 6072 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2168__107
timestamp 1667941163
transform -1 0 5244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2168_
timestamp 1667941163
transform 1 0 4140 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2169_
timestamp 1667941163
transform 1 0 24564 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2169__108
timestamp 1667941163
transform 1 0 24472 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2170__109
timestamp 1667941163
transform -1 0 25576 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2170_
timestamp 1667941163
transform 1 0 24748 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2171__110
timestamp 1667941163
transform -1 0 48024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2171_
timestamp 1667941163
transform -1 0 47288 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2172__111
timestamp 1667941163
transform 1 0 47748 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2172_
timestamp 1667941163
transform -1 0 48392 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2173__112
timestamp 1667941163
transform 1 0 28520 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2173_
timestamp 1667941163
transform 1 0 29164 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2174_
timestamp 1667941163
transform 1 0 42596 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2174__113
timestamp 1667941163
transform 1 0 41676 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2175_
timestamp 1667941163
transform 1 0 46460 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2175__114
timestamp 1667941163
transform -1 0 48024 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2176__115
timestamp 1667941163
transform -1 0 5796 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2176_
timestamp 1667941163
transform -1 0 3772 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2177_
timestamp 1667941163
transform 1 0 40572 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2177__116
timestamp 1667941163
transform -1 0 41308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2178__117
timestamp 1667941163
transform 1 0 2116 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2178_
timestamp 1667941163
transform -1 0 3496 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2179__118
timestamp 1667941163
transform -1 0 44988 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2179_
timestamp 1667941163
transform -1 0 44712 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2180__119
timestamp 1667941163
transform -1 0 10764 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2180_
timestamp 1667941163
transform 1 0 10488 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2181_
timestamp 1667941163
transform -1 0 3496 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2181__120
timestamp 1667941163
transform 1 0 2116 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2182_
timestamp 1667941163
transform 1 0 2024 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2182__121
timestamp 1667941163
transform -1 0 2300 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2183__122
timestamp 1667941163
transform -1 0 2300 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2183_
timestamp 1667941163
transform 1 0 2024 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i
timestamp 1667941163
transform -1 0 30360 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_wb_clk_i
timestamp 1667941163
transform 1 0 16284 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_wb_clk_i
timestamp 1667941163
transform -1 0 16376 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_wb_clk_i
timestamp 1667941163
transform -1 0 21528 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_wb_clk_i
timestamp 1667941163
transform 1 0 21160 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_wb_clk_i
timestamp 1667941163
transform 1 0 17664 0 -1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_wb_clk_i
timestamp 1667941163
transform -1 0 18492 0 1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_wb_clk_i
timestamp 1667941163
transform -1 0 25852 0 -1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_wb_clk_i
timestamp 1667941163
transform -1 0 24748 0 -1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_wb_clk_i
timestamp 1667941163
transform -1 0 31832 0 -1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_wb_clk_i
timestamp 1667941163
transform 1 0 32016 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_wb_clk_i
timestamp 1667941163
transform 1 0 36708 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_wb_clk_i
timestamp 1667941163
transform 1 0 37628 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_wb_clk_i
timestamp 1667941163
transform 1 0 33856 0 -1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_wb_clk_i
timestamp 1667941163
transform 1 0 34868 0 1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_wb_clk_i
timestamp 1667941163
transform 1 0 40112 0 1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_wb_clk_i
timestamp 1667941163
transform 1 0 39928 0 -1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1667941163
transform 1 0 7176 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1667941163
transform 1 0 9108 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input3
timestamp 1667941163
transform -1 0 48392 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1667941163
transform 1 0 32292 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1667941163
transform 1 0 24564 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input6
timestamp 1667941163
transform 1 0 43884 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input7
timestamp 1667941163
transform 1 0 17480 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input8
timestamp 1667941163
transform 1 0 20056 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input9
timestamp 1667941163
transform 1 0 1564 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input10
timestamp 1667941163
transform -1 0 48392 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input11
timestamp 1667941163
transform -1 0 48392 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input12
timestamp 1667941163
transform 1 0 1564 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input13
timestamp 1667941163
transform 1 0 14260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input14
timestamp 1667941163
transform 1 0 1564 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1667941163
transform -1 0 48392 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1667941163
transform 1 0 1564 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input18
timestamp 1667941163
transform 1 0 3956 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input19
timestamp 1667941163
transform 1 0 11684 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input20
timestamp 1667941163
transform 1 0 1564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1667941163
transform -1 0 39100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1667941163
transform -1 0 1840 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input23
timestamp 1667941163
transform 1 0 42596 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1667941163
transform -1 0 48392 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input25
timestamp 1667941163
transform 1 0 19412 0 1 46784
box -38 -48 406 592
<< labels >>
flabel metal3 s 200 46188 800 46428 0 FreeSans 960 0 0 0 active
port 0 nsew signal input
flabel metal2 s 15446 200 15558 800 0 FreeSans 448 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 27682 49200 27794 49800 0 FreeSans 448 90 0 0 io_in[10]
port 2 nsew signal input
flabel metal2 s -10 49200 102 49800 0 FreeSans 448 90 0 0 io_in[11]
port 3 nsew signal input
flabel metal3 s 49200 42108 49800 42348 0 FreeSans 960 0 0 0 io_in[12]
port 4 nsew signal input
flabel metal2 s 23818 200 23930 800 0 FreeSans 448 90 0 0 io_in[13]
port 5 nsew signal input
flabel metal2 s 18666 49200 18778 49800 0 FreeSans 448 90 0 0 io_in[14]
port 6 nsew signal input
flabel metal3 s 49200 44148 49800 44388 0 FreeSans 960 0 0 0 io_in[15]
port 7 nsew signal input
flabel metal3 s 49200 4028 49800 4268 0 FreeSans 960 0 0 0 io_in[16]
port 8 nsew signal input
flabel metal2 s 10294 49200 10406 49800 0 FreeSans 448 90 0 0 io_in[17]
port 9 nsew signal input
flabel metal2 s 12226 49200 12338 49800 0 FreeSans 448 90 0 0 io_in[18]
port 10 nsew signal input
flabel metal2 s 43138 200 43250 800 0 FreeSans 448 90 0 0 io_in[19]
port 11 nsew signal input
flabel metal3 s 200 16268 800 16508 0 FreeSans 960 0 0 0 io_in[1]
port 12 nsew signal input
flabel metal3 s 200 29188 800 29428 0 FreeSans 960 0 0 0 io_in[20]
port 13 nsew signal input
flabel metal3 s 200 18988 800 19228 0 FreeSans 960 0 0 0 io_in[21]
port 14 nsew signal input
flabel metal3 s 49200 15588 49800 15828 0 FreeSans 960 0 0 0 io_in[22]
port 15 nsew signal input
flabel metal2 s 9006 49200 9118 49800 0 FreeSans 448 90 0 0 io_in[23]
port 16 nsew signal input
flabel metal2 s 6430 49200 6542 49800 0 FreeSans 448 90 0 0 io_in[24]
port 17 nsew signal input
flabel metal2 s 37342 200 37454 800 0 FreeSans 448 90 0 0 io_in[25]
port 18 nsew signal input
flabel metal2 s 36698 200 36810 800 0 FreeSans 448 90 0 0 io_in[26]
port 19 nsew signal input
flabel metal3 s 49200 10828 49800 11068 0 FreeSans 960 0 0 0 io_in[27]
port 20 nsew signal input
flabel metal2 s 32834 200 32946 800 0 FreeSans 448 90 0 0 io_in[28]
port 21 nsew signal input
flabel metal2 s 49578 49200 49690 49800 0 FreeSans 448 90 0 0 io_in[29]
port 22 nsew signal input
flabel metal2 s 16090 200 16202 800 0 FreeSans 448 90 0 0 io_in[2]
port 23 nsew signal input
flabel metal3 s 49200 19668 49800 19908 0 FreeSans 960 0 0 0 io_in[30]
port 24 nsew signal input
flabel metal3 s 200 44148 800 44388 0 FreeSans 960 0 0 0 io_in[31]
port 25 nsew signal input
flabel metal2 s 30902 200 31014 800 0 FreeSans 448 90 0 0 io_in[32]
port 26 nsew signal input
flabel metal3 s 200 25788 800 26028 0 FreeSans 960 0 0 0 io_in[33]
port 27 nsew signal input
flabel metal2 s 37986 49200 38098 49800 0 FreeSans 448 90 0 0 io_in[34]
port 28 nsew signal input
flabel metal2 s 43138 49200 43250 49800 0 FreeSans 448 90 0 0 io_in[35]
port 29 nsew signal input
flabel metal3 s 49200 31228 49800 31468 0 FreeSans 960 0 0 0 io_in[36]
port 30 nsew signal input
flabel metal2 s 44426 49200 44538 49800 0 FreeSans 448 90 0 0 io_in[37]
port 31 nsew signal input
flabel metal2 s 28970 49200 29082 49800 0 FreeSans 448 90 0 0 io_in[3]
port 32 nsew signal input
flabel metal3 s 49200 30548 49800 30788 0 FreeSans 960 0 0 0 io_in[4]
port 33 nsew signal input
flabel metal3 s 49200 48228 49800 48468 0 FreeSans 960 0 0 0 io_in[5]
port 34 nsew signal input
flabel metal3 s 200 30548 800 30788 0 FreeSans 960 0 0 0 io_in[6]
port 35 nsew signal input
flabel metal3 s 200 21028 800 21268 0 FreeSans 960 0 0 0 io_in[7]
port 36 nsew signal input
flabel metal3 s 49200 33268 49800 33508 0 FreeSans 960 0 0 0 io_in[8]
port 37 nsew signal input
flabel metal2 s 8362 49200 8474 49800 0 FreeSans 448 90 0 0 io_in[9]
port 38 nsew signal input
flabel metal2 s 26394 200 26506 800 0 FreeSans 448 90 0 0 io_oeb[0]
port 39 nsew signal bidirectional
flabel metal3 s 200 16948 800 17188 0 FreeSans 960 0 0 0 io_oeb[10]
port 40 nsew signal bidirectional
flabel metal3 s 49200 28508 49800 28748 0 FreeSans 960 0 0 0 io_oeb[11]
port 41 nsew signal bidirectional
flabel metal3 s 49200 14908 49800 15148 0 FreeSans 960 0 0 0 io_oeb[12]
port 42 nsew signal bidirectional
flabel metal3 s 49200 13548 49800 13788 0 FreeSans 960 0 0 0 io_oeb[13]
port 43 nsew signal bidirectional
flabel metal3 s 200 4708 800 4948 0 FreeSans 960 0 0 0 io_oeb[14]
port 44 nsew signal bidirectional
flabel metal2 s 14158 49200 14270 49800 0 FreeSans 448 90 0 0 io_oeb[15]
port 45 nsew signal bidirectional
flabel metal3 s 49200 1988 49800 2228 0 FreeSans 960 0 0 0 io_oeb[16]
port 46 nsew signal bidirectional
flabel metal2 s 13514 200 13626 800 0 FreeSans 448 90 0 0 io_oeb[17]
port 47 nsew signal bidirectional
flabel metal2 s 36054 49200 36166 49800 0 FreeSans 448 90 0 0 io_oeb[18]
port 48 nsew signal bidirectional
flabel metal2 s 14802 49200 14914 49800 0 FreeSans 448 90 0 0 io_oeb[19]
port 49 nsew signal bidirectional
flabel metal2 s 39274 200 39386 800 0 FreeSans 448 90 0 0 io_oeb[1]
port 50 nsew signal bidirectional
flabel metal3 s 49200 21708 49800 21948 0 FreeSans 960 0 0 0 io_oeb[20]
port 51 nsew signal bidirectional
flabel metal2 s 1922 49200 2034 49800 0 FreeSans 448 90 0 0 io_oeb[21]
port 52 nsew signal bidirectional
flabel metal2 s 5142 200 5254 800 0 FreeSans 448 90 0 0 io_oeb[22]
port 53 nsew signal bidirectional
flabel metal2 s 25106 49200 25218 49800 0 FreeSans 448 90 0 0 io_oeb[23]
port 54 nsew signal bidirectional
flabel metal2 s 25750 49200 25862 49800 0 FreeSans 448 90 0 0 io_oeb[24]
port 55 nsew signal bidirectional
flabel metal2 s 47646 200 47758 800 0 FreeSans 448 90 0 0 io_oeb[25]
port 56 nsew signal bidirectional
flabel metal3 s 49200 39388 49800 39628 0 FreeSans 960 0 0 0 io_oeb[26]
port 57 nsew signal bidirectional
flabel metal2 s 29614 49200 29726 49800 0 FreeSans 448 90 0 0 io_oeb[27]
port 58 nsew signal bidirectional
flabel metal2 s 41850 200 41962 800 0 FreeSans 448 90 0 0 io_oeb[28]
port 59 nsew signal bidirectional
flabel metal3 s 49200 32588 49800 32828 0 FreeSans 960 0 0 0 io_oeb[29]
port 60 nsew signal bidirectional
flabel metal2 s 41850 49200 41962 49800 0 FreeSans 448 90 0 0 io_oeb[2]
port 61 nsew signal bidirectional
flabel metal2 s 2566 49200 2678 49800 0 FreeSans 448 90 0 0 io_oeb[30]
port 62 nsew signal bidirectional
flabel metal2 s 41206 200 41318 800 0 FreeSans 448 90 0 0 io_oeb[31]
port 63 nsew signal bidirectional
flabel metal3 s 200 25108 800 25348 0 FreeSans 960 0 0 0 io_oeb[32]
port 64 nsew signal bidirectional
flabel metal2 s 48934 200 49046 800 0 FreeSans 448 90 0 0 io_oeb[33]
port 65 nsew signal bidirectional
flabel metal2 s 10938 49200 11050 49800 0 FreeSans 448 90 0 0 io_oeb[34]
port 66 nsew signal bidirectional
flabel metal3 s 200 21708 800 21948 0 FreeSans 960 0 0 0 io_oeb[35]
port 67 nsew signal bidirectional
flabel metal3 s 200 11508 800 11748 0 FreeSans 960 0 0 0 io_oeb[36]
port 68 nsew signal bidirectional
flabel metal3 s 200 18308 800 18548 0 FreeSans 960 0 0 0 io_oeb[37]
port 69 nsew signal bidirectional
flabel metal2 s 25750 200 25862 800 0 FreeSans 448 90 0 0 io_oeb[3]
port 70 nsew signal bidirectional
flabel metal3 s 49200 -52 49800 188 0 FreeSans 960 0 0 0 io_oeb[4]
port 71 nsew signal bidirectional
flabel metal3 s 200 32588 800 32828 0 FreeSans 960 0 0 0 io_oeb[5]
port 72 nsew signal bidirectional
flabel metal3 s 49200 17628 49800 17868 0 FreeSans 960 0 0 0 io_oeb[6]
port 73 nsew signal bidirectional
flabel metal2 s 12870 49200 12982 49800 0 FreeSans 448 90 0 0 io_oeb[7]
port 74 nsew signal bidirectional
flabel metal2 s 4498 200 4610 800 0 FreeSans 448 90 0 0 io_oeb[8]
port 75 nsew signal bidirectional
flabel metal2 s 10938 200 11050 800 0 FreeSans 448 90 0 0 io_oeb[9]
port 76 nsew signal bidirectional
flabel metal3 s 49200 46868 49800 47108 0 FreeSans 960 0 0 0 io_out[0]
port 77 nsew signal bidirectional
flabel metal3 s 49200 27828 49800 28068 0 FreeSans 960 0 0 0 io_out[10]
port 78 nsew signal bidirectional
flabel metal3 s 200 2668 800 2908 0 FreeSans 960 0 0 0 io_out[11]
port 79 nsew signal bidirectional
flabel metal3 s 200 7428 800 7668 0 FreeSans 960 0 0 0 io_out[12]
port 80 nsew signal bidirectional
flabel metal2 s 40562 200 40674 800 0 FreeSans 448 90 0 0 io_out[13]
port 81 nsew signal bidirectional
flabel metal3 s 49200 40068 49800 40308 0 FreeSans 960 0 0 0 io_out[14]
port 82 nsew signal bidirectional
flabel metal3 s 200 41428 800 41668 0 FreeSans 960 0 0 0 io_out[15]
port 83 nsew signal bidirectional
flabel metal3 s 49200 26468 49800 26708 0 FreeSans 960 0 0 0 io_out[16]
port 84 nsew signal bidirectional
flabel metal2 s 46358 49200 46470 49800 0 FreeSans 448 90 0 0 io_out[17]
port 85 nsew signal bidirectional
flabel metal2 s 47002 200 47114 800 0 FreeSans 448 90 0 0 io_out[18]
port 86 nsew signal bidirectional
flabel metal3 s 200 23748 800 23988 0 FreeSans 960 0 0 0 io_out[19]
port 87 nsew signal bidirectional
flabel metal2 s 33478 49200 33590 49800 0 FreeSans 448 90 0 0 io_out[1]
port 88 nsew signal bidirectional
flabel metal2 s 40562 49200 40674 49800 0 FreeSans 448 90 0 0 io_out[20]
port 89 nsew signal bidirectional
flabel metal3 s 200 40748 800 40988 0 FreeSans 960 0 0 0 io_out[21]
port 90 nsew signal bidirectional
flabel metal2 s 32190 200 32302 800 0 FreeSans 448 90 0 0 io_out[22]
port 91 nsew signal bidirectional
flabel metal3 s 49200 22388 49800 22628 0 FreeSans 960 0 0 0 io_out[23]
port 92 nsew signal bidirectional
flabel metal2 s 27682 200 27794 800 0 FreeSans 448 90 0 0 io_out[24]
port 93 nsew signal bidirectional
flabel metal2 s 36698 49200 36810 49800 0 FreeSans 448 90 0 0 io_out[25]
port 94 nsew signal bidirectional
flabel metal3 s 200 5388 800 5628 0 FreeSans 960 0 0 0 io_out[26]
port 95 nsew signal bidirectional
flabel metal2 s 38630 49200 38742 49800 0 FreeSans 448 90 0 0 io_out[27]
port 96 nsew signal bidirectional
flabel metal2 s 17378 200 17490 800 0 FreeSans 448 90 0 0 io_out[28]
port 97 nsew signal bidirectional
flabel metal3 s 49200 1308 49800 1548 0 FreeSans 960 0 0 0 io_out[29]
port 98 nsew signal bidirectional
flabel metal2 s 7074 200 7186 800 0 FreeSans 448 90 0 0 io_out[2]
port 99 nsew signal bidirectional
flabel metal3 s 200 6748 800 6988 0 FreeSans 960 0 0 0 io_out[30]
port 100 nsew signal bidirectional
flabel metal3 s 200 14228 800 14468 0 FreeSans 960 0 0 0 io_out[31]
port 101 nsew signal bidirectional
flabel metal3 s 200 47548 800 47788 0 FreeSans 960 0 0 0 io_out[32]
port 102 nsew signal bidirectional
flabel metal3 s 49200 6748 49800 6988 0 FreeSans 960 0 0 0 io_out[33]
port 103 nsew signal bidirectional
flabel metal3 s 49200 41428 49800 41668 0 FreeSans 960 0 0 0 io_out[34]
port 104 nsew signal bidirectional
flabel metal3 s 49200 38028 49800 38268 0 FreeSans 960 0 0 0 io_out[35]
port 105 nsew signal bidirectional
flabel metal2 s 15446 49200 15558 49800 0 FreeSans 448 90 0 0 io_out[36]
port 106 nsew signal bidirectional
flabel metal3 s 49200 44828 49800 45068 0 FreeSans 960 0 0 0 io_out[37]
port 107 nsew signal bidirectional
flabel metal3 s 200 43468 800 43708 0 FreeSans 960 0 0 0 io_out[3]
port 108 nsew signal bidirectional
flabel metal3 s 49200 29188 49800 29428 0 FreeSans 960 0 0 0 io_out[4]
port 109 nsew signal bidirectional
flabel metal2 s 23174 49200 23286 49800 0 FreeSans 448 90 0 0 io_out[5]
port 110 nsew signal bidirectional
flabel metal2 s 48290 49200 48402 49800 0 FreeSans 448 90 0 0 io_out[6]
port 111 nsew signal bidirectional
flabel metal3 s 200 20348 800 20588 0 FreeSans 960 0 0 0 io_out[7]
port 112 nsew signal bidirectional
flabel metal2 s 19310 200 19422 800 0 FreeSans 448 90 0 0 io_out[8]
port 113 nsew signal bidirectional
flabel metal3 s 200 14908 800 15148 0 FreeSans 960 0 0 0 io_out[9]
port 114 nsew signal bidirectional
flabel metal3 s 49200 8108 49800 8348 0 FreeSans 960 0 0 0 la1_data_in[0]
port 115 nsew signal input
flabel metal2 s 21886 200 21998 800 0 FreeSans 448 90 0 0 la1_data_in[10]
port 116 nsew signal input
flabel metal3 s 49200 6068 49800 6308 0 FreeSans 960 0 0 0 la1_data_in[11]
port 117 nsew signal input
flabel metal3 s 200 37348 800 37588 0 FreeSans 960 0 0 0 la1_data_in[12]
port 118 nsew signal input
flabel metal2 s 34122 200 34234 800 0 FreeSans 448 90 0 0 la1_data_in[13]
port 119 nsew signal input
flabel metal3 s 200 13548 800 13788 0 FreeSans 960 0 0 0 la1_data_in[14]
port 120 nsew signal input
flabel metal2 s 16734 49200 16846 49800 0 FreeSans 448 90 0 0 la1_data_in[15]
port 121 nsew signal input
flabel metal2 s 31546 49200 31658 49800 0 FreeSans 448 90 0 0 la1_data_in[16]
port 122 nsew signal input
flabel metal2 s 23818 49200 23930 49800 0 FreeSans 448 90 0 0 la1_data_in[17]
port 123 nsew signal input
flabel metal2 s 43782 200 43894 800 0 FreeSans 448 90 0 0 la1_data_in[18]
port 124 nsew signal input
flabel metal2 s 17378 49200 17490 49800 0 FreeSans 448 90 0 0 la1_data_in[19]
port 125 nsew signal input
flabel metal2 s 19954 200 20066 800 0 FreeSans 448 90 0 0 la1_data_in[1]
port 126 nsew signal input
flabel metal3 s 200 36668 800 36908 0 FreeSans 960 0 0 0 la1_data_in[20]
port 127 nsew signal input
flabel metal2 s 48934 49200 49046 49800 0 FreeSans 448 90 0 0 la1_data_in[21]
port 128 nsew signal input
flabel metal3 s 49200 8788 49800 9028 0 FreeSans 960 0 0 0 la1_data_in[22]
port 129 nsew signal input
flabel metal3 s 200 628 800 868 0 FreeSans 960 0 0 0 la1_data_in[23]
port 130 nsew signal input
flabel metal2 s 14158 200 14270 800 0 FreeSans 448 90 0 0 la1_data_in[24]
port 131 nsew signal input
flabel metal3 s 200 38708 800 38948 0 FreeSans 960 0 0 0 la1_data_in[25]
port 132 nsew signal input
flabel metal3 s 49200 3348 49800 3588 0 FreeSans 960 0 0 0 la1_data_in[26]
port 133 nsew signal input
flabel metal2 s 28970 200 29082 800 0 FreeSans 448 90 0 0 la1_data_in[27]
port 134 nsew signal input
flabel metal3 s 200 33948 800 34188 0 FreeSans 960 0 0 0 la1_data_in[28]
port 135 nsew signal input
flabel metal2 s 1278 49200 1390 49800 0 FreeSans 448 90 0 0 la1_data_in[29]
port 136 nsew signal input
flabel metal2 s 11582 200 11694 800 0 FreeSans 448 90 0 0 la1_data_in[2]
port 137 nsew signal input
flabel metal2 s 1278 200 1390 800 0 FreeSans 448 90 0 0 la1_data_in[30]
port 138 nsew signal input
flabel metal2 s 38630 200 38742 800 0 FreeSans 448 90 0 0 la1_data_in[31]
port 139 nsew signal input
flabel metal3 s 200 31908 800 32148 0 FreeSans 960 0 0 0 la1_data_in[3]
port 140 nsew signal input
flabel metal2 s 42494 49200 42606 49800 0 FreeSans 448 90 0 0 la1_data_in[4]
port 141 nsew signal input
flabel metal3 s 49200 24428 49800 24668 0 FreeSans 960 0 0 0 la1_data_in[5]
port 142 nsew signal input
flabel metal2 s 19310 49200 19422 49800 0 FreeSans 448 90 0 0 la1_data_in[6]
port 143 nsew signal input
flabel metal3 s 200 23068 800 23308 0 FreeSans 960 0 0 0 la1_data_in[7]
port 144 nsew signal input
flabel metal2 s 20598 49200 20710 49800 0 FreeSans 448 90 0 0 la1_data_in[8]
port 145 nsew signal input
flabel metal3 s 200 34628 800 34868 0 FreeSans 960 0 0 0 la1_data_in[9]
port 146 nsew signal input
flabel metal2 s 7718 200 7830 800 0 FreeSans 448 90 0 0 la1_data_out[0]
port 147 nsew signal bidirectional
flabel metal3 s 49200 12188 49800 12428 0 FreeSans 960 0 0 0 la1_data_out[10]
port 148 nsew signal bidirectional
flabel metal2 s 22530 200 22642 800 0 FreeSans 448 90 0 0 la1_data_out[11]
port 149 nsew signal bidirectional
flabel metal3 s 49200 46188 49800 46428 0 FreeSans 960 0 0 0 la1_data_out[12]
port 150 nsew signal bidirectional
flabel metal2 s 4498 49200 4610 49800 0 FreeSans 448 90 0 0 la1_data_out[13]
port 151 nsew signal bidirectional
flabel metal2 s 27038 49200 27150 49800 0 FreeSans 448 90 0 0 la1_data_out[14]
port 152 nsew signal bidirectional
flabel metal3 s 200 1308 800 1548 0 FreeSans 960 0 0 0 la1_data_out[15]
port 153 nsew signal bidirectional
flabel metal3 s 49200 16948 49800 17188 0 FreeSans 960 0 0 0 la1_data_out[16]
port 154 nsew signal bidirectional
flabel metal3 s 49200 35988 49800 36228 0 FreeSans 960 0 0 0 la1_data_out[17]
port 155 nsew signal bidirectional
flabel metal2 s 5786 49200 5898 49800 0 FreeSans 448 90 0 0 la1_data_out[18]
port 156 nsew signal bidirectional
flabel metal3 s 49200 25788 49800 26028 0 FreeSans 960 0 0 0 la1_data_out[19]
port 157 nsew signal bidirectional
flabel metal3 s 200 45508 800 45748 0 FreeSans 960 0 0 0 la1_data_out[1]
port 158 nsew signal bidirectional
flabel metal3 s 200 10148 800 10388 0 FreeSans 960 0 0 0 la1_data_out[20]
port 159 nsew signal bidirectional
flabel metal3 s 49200 42788 49800 43028 0 FreeSans 960 0 0 0 la1_data_out[21]
port 160 nsew signal bidirectional
flabel metal2 s 30258 49200 30370 49800 0 FreeSans 448 90 0 0 la1_data_out[22]
port 161 nsew signal bidirectional
flabel metal2 s 12870 200 12982 800 0 FreeSans 448 90 0 0 la1_data_out[23]
port 162 nsew signal bidirectional
flabel metal3 s 49200 18988 49800 19228 0 FreeSans 960 0 0 0 la1_data_out[24]
port 163 nsew signal bidirectional
flabel metal3 s 200 3348 800 3588 0 FreeSans 960 0 0 0 la1_data_out[25]
port 164 nsew signal bidirectional
flabel metal3 s 49200 5388 49800 5628 0 FreeSans 960 0 0 0 la1_data_out[26]
port 165 nsew signal bidirectional
flabel metal3 s 200 48228 800 48468 0 FreeSans 960 0 0 0 la1_data_out[27]
port 166 nsew signal bidirectional
flabel metal2 s 45070 200 45182 800 0 FreeSans 448 90 0 0 la1_data_out[28]
port 167 nsew signal bidirectional
flabel metal2 s 6430 200 6542 800 0 FreeSans 448 90 0 0 la1_data_out[29]
port 168 nsew signal bidirectional
flabel metal2 s 20598 200 20710 800 0 FreeSans 448 90 0 0 la1_data_out[2]
port 169 nsew signal bidirectional
flabel metal3 s 49200 12868 49800 13108 0 FreeSans 960 0 0 0 la1_data_out[30]
port 170 nsew signal bidirectional
flabel metal3 s 49200 48908 49800 49148 0 FreeSans 960 0 0 0 la1_data_out[31]
port 171 nsew signal bidirectional
flabel metal3 s 200 9468 800 9708 0 FreeSans 960 0 0 0 la1_data_out[3]
port 172 nsew signal bidirectional
flabel metal2 s 45714 200 45826 800 0 FreeSans 448 90 0 0 la1_data_out[4]
port 173 nsew signal bidirectional
flabel metal2 s 3210 200 3322 800 0 FreeSans 448 90 0 0 la1_data_out[5]
port 174 nsew signal bidirectional
flabel metal3 s 49200 20348 49800 20588 0 FreeSans 960 0 0 0 la1_data_out[6]
port 175 nsew signal bidirectional
flabel metal2 s 634 200 746 800 0 FreeSans 448 90 0 0 la1_data_out[7]
port 176 nsew signal bidirectional
flabel metal3 s 49200 37348 49800 37588 0 FreeSans 960 0 0 0 la1_data_out[8]
port 177 nsew signal bidirectional
flabel metal2 s 47002 49200 47114 49800 0 FreeSans 448 90 0 0 la1_data_out[9]
port 178 nsew signal bidirectional
flabel metal2 s 49578 200 49690 800 0 FreeSans 448 90 0 0 la1_oenb[0]
port 179 nsew signal input
flabel metal2 s 45070 49200 45182 49800 0 FreeSans 448 90 0 0 la1_oenb[10]
port 180 nsew signal input
flabel metal3 s 200 27828 800 28068 0 FreeSans 960 0 0 0 la1_oenb[11]
port 181 nsew signal input
flabel metal3 s 200 29868 800 30108 0 FreeSans 960 0 0 0 la1_oenb[12]
port 182 nsew signal input
flabel metal2 s 30258 200 30370 800 0 FreeSans 448 90 0 0 la1_oenb[13]
port 183 nsew signal input
flabel metal2 s -10 200 102 800 0 FreeSans 448 90 0 0 la1_oenb[14]
port 184 nsew signal input
flabel metal2 s 35410 200 35522 800 0 FreeSans 448 90 0 0 la1_oenb[15]
port 185 nsew signal input
flabel metal3 s 200 35988 800 36228 0 FreeSans 960 0 0 0 la1_oenb[16]
port 186 nsew signal input
flabel metal2 s 3854 49200 3966 49800 0 FreeSans 448 90 0 0 la1_oenb[17]
port 187 nsew signal input
flabel metal2 s 21886 49200 21998 49800 0 FreeSans 448 90 0 0 la1_oenb[18]
port 188 nsew signal input
flabel metal3 s 200 27148 800 27388 0 FreeSans 960 0 0 0 la1_oenb[19]
port 189 nsew signal input
flabel metal2 s 9006 200 9118 800 0 FreeSans 448 90 0 0 la1_oenb[1]
port 190 nsew signal input
flabel metal2 s 2566 200 2678 800 0 FreeSans 448 90 0 0 la1_oenb[20]
port 191 nsew signal input
flabel metal2 s 32190 49200 32302 49800 0 FreeSans 448 90 0 0 la1_oenb[21]
port 192 nsew signal input
flabel metal2 s 21242 49200 21354 49800 0 FreeSans 448 90 0 0 la1_oenb[22]
port 193 nsew signal input
flabel metal2 s 24462 200 24574 800 0 FreeSans 448 90 0 0 la1_oenb[23]
port 194 nsew signal input
flabel metal2 s 39918 49200 40030 49800 0 FreeSans 448 90 0 0 la1_oenb[24]
port 195 nsew signal input
flabel metal3 s 49200 10148 49800 10388 0 FreeSans 960 0 0 0 la1_oenb[25]
port 196 nsew signal input
flabel metal3 s 200 39388 800 39628 0 FreeSans 960 0 0 0 la1_oenb[26]
port 197 nsew signal input
flabel metal3 s 49200 35308 49800 35548 0 FreeSans 960 0 0 0 la1_oenb[27]
port 198 nsew signal input
flabel metal2 s 9650 200 9762 800 0 FreeSans 448 90 0 0 la1_oenb[28]
port 199 nsew signal input
flabel metal2 s 18022 200 18134 800 0 FreeSans 448 90 0 0 la1_oenb[29]
port 200 nsew signal input
flabel metal3 s 200 8108 800 8348 0 FreeSans 960 0 0 0 la1_oenb[2]
port 201 nsew signal input
flabel metal3 s 49200 34628 49800 34868 0 FreeSans 960 0 0 0 la1_oenb[30]
port 202 nsew signal input
flabel metal2 s 28326 200 28438 800 0 FreeSans 448 90 0 0 la1_oenb[31]
port 203 nsew signal input
flabel metal2 s 35410 49200 35522 49800 0 FreeSans 448 90 0 0 la1_oenb[3]
port 204 nsew signal input
flabel metal2 s 34122 49200 34234 49800 0 FreeSans 448 90 0 0 la1_oenb[4]
port 205 nsew signal input
flabel metal3 s 200 49588 800 49828 0 FreeSans 960 0 0 0 la1_oenb[5]
port 206 nsew signal input
flabel metal2 s 7718 49200 7830 49800 0 FreeSans 448 90 0 0 la1_oenb[6]
port 207 nsew signal input
flabel metal2 s 34766 200 34878 800 0 FreeSans 448 90 0 0 la1_oenb[7]
port 208 nsew signal input
flabel metal3 s 200 12188 800 12428 0 FreeSans 960 0 0 0 la1_oenb[8]
port 209 nsew signal input
flabel metal3 s 200 42788 800 43028 0 FreeSans 960 0 0 0 la1_oenb[9]
port 210 nsew signal input
flabel metal4 s 4208 2128 4528 47376 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 34928 2128 35248 47376 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 19568 2128 19888 47376 0 FreeSans 1920 90 0 0 vssd1
port 212 nsew ground bidirectional
flabel metal3 s 49200 23748 49800 23988 0 FreeSans 960 0 0 0 wb_clk_i
port 213 nsew signal input
rlabel metal1 24978 47328 24978 47328 0 vccd1
rlabel metal1 24978 46784 24978 46784 0 vssd1
rlabel metal2 12926 30498 12926 30498 0 _0000_
rlabel via1 10805 30702 10805 30702 0 _0001_
rlabel metal1 10023 30294 10023 30294 0 _0002_
rlabel metal1 10023 32470 10023 32470 0 _0003_
rlabel via1 8413 29206 8413 29206 0 _0004_
rlabel via1 9057 26962 9057 26962 0 _0005_
rlabel metal1 10207 24106 10207 24106 0 _0006_
rlabel metal2 8878 24310 8878 24310 0 _0007_
rlabel metal2 7130 25670 7130 25670 0 _0008_
rlabel metal1 6072 27098 6072 27098 0 _0009_
rlabel metal2 12374 32300 12374 32300 0 _0010_
rlabel metal1 10212 30702 10212 30702 0 _0011_
rlabel metal1 9338 30226 9338 30226 0 _0012_
rlabel metal1 9108 31994 9108 31994 0 _0013_
rlabel metal2 8142 28900 8142 28900 0 _0014_
rlabel metal1 8556 26894 8556 26894 0 _0015_
rlabel metal1 8878 24242 8878 24242 0 _0016_
rlabel metal1 7912 24718 7912 24718 0 _0017_
rlabel metal2 6486 25636 6486 25636 0 _0018_
rlabel metal1 5842 27404 5842 27404 0 _0019_
rlabel metal2 6026 32708 6026 32708 0 _0020_
rlabel metal2 7406 33660 7406 33660 0 _0021_
rlabel metal2 9430 34204 9430 34204 0 _0022_
rlabel metal2 4186 33796 4186 33796 0 _0023_
rlabel metal2 4370 34884 4370 34884 0 _0024_
rlabel metal1 4232 36346 4232 36346 0 _0025_
rlabel metal2 4830 37468 4830 37468 0 _0026_
rlabel metal2 6578 38012 6578 38012 0 _0027_
rlabel metal1 8188 36754 8188 36754 0 _0028_
rlabel metal1 9016 36074 9016 36074 0 _0029_
rlabel metal2 28934 31110 28934 31110 0 _0030_
rlabel viali 32342 28458 32342 28458 0 _0031_
rlabel metal1 35548 31790 35548 31790 0 _0032_
rlabel metal2 32798 33762 32798 33762 0 _0033_
rlabel metal2 38318 32198 38318 32198 0 _0034_
rlabel metal1 38900 29546 38900 29546 0 _0035_
rlabel metal1 40066 25806 40066 25806 0 _0036_
rlabel metal1 35277 26282 35277 26282 0 _0037_
rlabel metal1 36156 23834 36156 23834 0 _0038_
rlabel metal2 33350 21794 33350 21794 0 _0039_
rlabel metal2 32338 19618 32338 19618 0 _0040_
rlabel metal1 37770 18258 37770 18258 0 _0041_
rlabel metal1 33948 15674 33948 15674 0 _0042_
rlabel metal2 32614 14790 32614 14790 0 _0043_
rlabel metal1 38092 12886 38092 12886 0 _0044_
rlabel via1 33437 10642 33437 10642 0 _0045_
rlabel metal2 22126 32198 22126 32198 0 _0046_
rlabel metal2 20194 31586 20194 31586 0 _0047_
rlabel metal1 16463 33898 16463 33898 0 _0048_
rlabel metal2 16882 34850 16882 34850 0 _0049_
rlabel via1 25249 32878 25249 32878 0 _0050_
rlabel metal2 28014 36550 28014 36550 0 _0051_
rlabel metal1 27569 37162 27569 37162 0 _0052_
rlabel metal2 23690 34850 23690 34850 0 _0053_
rlabel metal2 20930 37026 20930 37026 0 _0054_
rlabel metal2 18722 38114 18722 38114 0 _0055_
rlabel via1 24881 38318 24881 38318 0 _0056_
rlabel via1 23409 37842 23409 37842 0 _0057_
rlabel via1 13197 36822 13197 36822 0 _0058_
rlabel metal1 12880 37978 12880 37978 0 _0059_
rlabel metal1 15778 37978 15778 37978 0 _0060_
rlabel via1 14034 34578 14034 34578 0 _0061_
rlabel metal2 23322 29988 23322 29988 0 _0062_
rlabel via1 26261 29614 26261 29614 0 _0063_
rlabel metal2 22586 22406 22586 22406 0 _0064_
rlabel metal2 20010 26078 20010 26078 0 _0065_
rlabel metal2 17434 27846 17434 27846 0 _0066_
rlabel metal1 14761 24854 14761 24854 0 _0067_
rlabel metal2 16882 21692 16882 21692 0 _0068_
rlabel via1 14577 19754 14577 19754 0 _0069_
rlabel metal2 18538 17442 18538 17442 0 _0070_
rlabel via1 13473 13906 13473 13906 0 _0071_
rlabel metal2 25254 19142 25254 19142 0 _0072_
rlabel metal1 24881 15062 24881 15062 0 _0073_
rlabel metal2 20286 16354 20286 16354 0 _0074_
rlabel via1 16233 11050 16233 11050 0 _0075_
rlabel via1 19453 10710 19453 10710 0 _0076_
rlabel metal2 24886 10404 24886 10404 0 _0077_
rlabel metal1 29527 29138 29527 29138 0 _0078_
rlabel metal1 29435 28118 29435 28118 0 _0079_
rlabel metal1 33948 29750 33948 29750 0 _0080_
rlabel metal1 32057 29546 32057 29546 0 _0081_
rlabel metal1 34536 29138 34536 29138 0 _0082_
rlabel metal2 35006 28322 35006 28322 0 _0083_
rlabel metal2 31234 25670 31234 25670 0 _0084_
rlabel metal1 32292 25466 32292 25466 0 _0085_
rlabel metal1 33120 23290 33120 23290 0 _0086_
rlabel via1 29849 21522 29849 21522 0 _0087_
rlabel via1 28745 19414 28745 19414 0 _0088_
rlabel metal1 29113 17238 29113 17238 0 _0089_
rlabel metal1 28704 15674 28704 15674 0 _0090_
rlabel metal1 30912 14586 30912 14586 0 _0091_
rlabel via1 28009 12818 28009 12818 0 _0092_
rlabel metal1 30355 12886 30355 12886 0 _0093_
rlabel metal1 6573 32878 6573 32878 0 _0094_
rlabel metal1 7298 33558 7298 33558 0 _0095_
rlabel via1 9701 33966 9701 33966 0 _0096_
rlabel metal1 4825 33966 4825 33966 0 _0097_
rlabel metal2 5750 34850 5750 34850 0 _0098_
rlabel metal2 6026 36550 6026 36550 0 _0099_
rlabel metal1 4722 37162 4722 37162 0 _0100_
rlabel metal1 6424 37910 6424 37910 0 _0101_
rlabel metal1 8643 36822 8643 36822 0 _0102_
rlabel metal1 9721 35734 9721 35734 0 _0103_
rlabel metal1 43649 14314 43649 14314 0 _0104_
rlabel metal2 46690 16354 46690 16354 0 _0105_
rlabel metal1 45075 18326 45075 18326 0 _0106_
rlabel metal2 43746 20706 43746 20706 0 _0107_
rlabel metal1 39233 16490 39233 16490 0 _0108_
rlabel metal2 40526 14178 40526 14178 0 _0109_
rlabel metal1 38819 19346 38819 19346 0 _0110_
rlabel metal1 40066 19720 40066 19720 0 _0111_
rlabel via1 42462 21998 42462 21998 0 _0112_
rlabel via1 41625 24106 41625 24106 0 _0113_
rlabel metal1 44528 23834 44528 23834 0 _0114_
rlabel metal2 44206 26758 44206 26758 0 _0115_
rlabel metal1 45208 30702 45208 30702 0 _0116_
rlabel metal2 42642 31110 42642 31110 0 _0117_
rlabel metal1 44620 27642 44620 27642 0 _0118_
rlabel metal2 41814 27914 41814 27914 0 _0119_
rlabel metal1 15359 29546 15359 29546 0 _0120_
rlabel metal2 15686 31314 15686 31314 0 _0121_
rlabel metal1 17812 30702 17812 30702 0 _0122_
rlabel metal1 13519 32470 13519 32470 0 _0123_
rlabel metal2 12282 33694 12282 33694 0 _0124_
rlabel via1 14494 29206 14494 29206 0 _0125_
rlabel metal2 11822 24582 11822 24582 0 _0126_
rlabel metal1 12010 22678 12010 22678 0 _0127_
rlabel metal2 12098 26078 12098 26078 0 _0128_
rlabel via1 12930 28118 12930 28118 0 _0129_
rlabel metal1 26261 25262 26261 25262 0 _0130_
rlabel metal1 30237 23766 30237 23766 0 _0131_
rlabel metal2 29394 34850 29394 34850 0 _0132_
rlabel via1 30033 32878 30033 32878 0 _0133_
rlabel metal2 36938 34850 36938 34850 0 _0134_
rlabel metal2 33074 35462 33074 35462 0 _0135_
rlabel metal2 38778 34340 38778 34340 0 _0136_
rlabel metal1 40240 31790 40240 31790 0 _0137_
rlabel via1 39242 24106 39242 24106 0 _0138_
rlabel metal1 32655 27030 32655 27030 0 _0139_
rlabel metal1 34868 23290 34868 23290 0 _0140_
rlabel via1 31229 21998 31229 21998 0 _0141_
rlabel via1 30493 18666 30493 18666 0 _0142_
rlabel metal1 31974 17578 31974 17578 0 _0143_
rlabel metal2 32430 15878 32430 15878 0 _0144_
rlabel metal1 32379 13226 32379 13226 0 _0145_
rlabel metal2 29578 10914 29578 10914 0 _0146_
rlabel metal1 32149 11118 32149 11118 0 _0147_
rlabel metal2 39054 22406 39054 22406 0 _0148_
rlabel metal1 25203 27370 25203 27370 0 _0149_
rlabel metal1 27135 27370 27135 27370 0 _0150_
rlabel metal1 24513 22678 24513 22678 0 _0151_
rlabel metal1 23317 25942 23317 25942 0 _0152_
rlabel via1 14393 26962 14393 26962 0 _0153_
rlabel metal2 14306 23494 14306 23494 0 _0154_
rlabel metal1 13933 21590 13933 21590 0 _0155_
rlabel via1 12185 19754 12185 19754 0 _0156_
rlabel metal2 12558 17884 12558 17884 0 _0157_
rlabel metal1 12088 17170 12088 17170 0 _0158_
rlabel metal1 26465 19414 26465 19414 0 _0159_
rlabel metal1 26454 14382 26454 14382 0 _0160_
rlabel metal1 17843 15062 17843 15062 0 _0161_
rlabel metal2 17066 13090 17066 13090 0 _0162_
rlabel metal1 17705 10710 17705 10710 0 _0163_
rlabel via1 28294 10642 28294 10642 0 _0164_
rlabel metal1 27360 32402 27360 32402 0 _0165_
rlabel via1 22305 28050 22305 28050 0 _0166_
rlabel via1 21569 29546 21569 29546 0 _0167_
rlabel metal1 23797 21590 23797 21590 0 _0168_
rlabel metal2 20102 28662 20102 28662 0 _0169_
rlabel metal2 19458 28968 19458 28968 0 _0170_
rlabel metal1 19448 23698 19448 23698 0 _0171_
rlabel metal1 20485 22678 20485 22678 0 _0172_
rlabel metal1 19448 20434 19448 20434 0 _0173_
rlabel metal2 22034 18938 22034 18938 0 _0174_
rlabel via1 19729 18734 19729 18734 0 _0175_
rlabel metal1 27937 18666 27937 18666 0 _0176_
rlabel metal1 26250 15402 26250 15402 0 _0177_
rlabel metal1 20270 17578 20270 17578 0 _0178_
rlabel metal1 20649 13906 20649 13906 0 _0179_
rlabel metal1 23087 13294 23087 13294 0 _0180_
rlabel metal1 26266 12410 26266 12410 0 _0181_
rlabel metal1 16330 14450 16330 14450 0 _0182_
rlabel metal1 15456 14314 15456 14314 0 _0183_
rlabel metal1 14076 14382 14076 14382 0 _0184_
rlabel metal2 23230 16456 23230 16456 0 _0185_
rlabel metal1 23506 17850 23506 17850 0 _0186_
rlabel metal2 23966 18564 23966 18564 0 _0187_
rlabel metal2 24058 16490 24058 16490 0 _0188_
rlabel metal1 24748 16082 24748 16082 0 _0189_
rlabel metal2 25254 16252 25254 16252 0 _0190_
rlabel metal1 21206 15130 21206 15130 0 _0191_
rlabel metal2 21482 15878 21482 15878 0 _0192_
rlabel metal2 20470 16252 20470 16252 0 _0193_
rlabel metal1 20102 13430 20102 13430 0 _0194_
rlabel metal1 20424 12750 20424 12750 0 _0195_
rlabel metal1 19044 12614 19044 12614 0 _0196_
rlabel metal2 17066 11900 17066 11900 0 _0197_
rlabel metal2 22494 11356 22494 11356 0 _0198_
rlabel metal2 22954 11730 22954 11730 0 _0199_
rlabel metal1 20562 9962 20562 9962 0 _0200_
rlabel metal1 19964 10234 19964 10234 0 _0201_
rlabel metal1 23322 10098 23322 10098 0 _0202_
rlabel metal2 23874 10302 23874 10302 0 _0203_
rlabel metal2 24978 11322 24978 11322 0 _0204_
rlabel metal2 24702 10506 24702 10506 0 _0205_
rlabel metal1 27554 23630 27554 23630 0 _0206_
rlabel metal1 28612 23086 28612 23086 0 _0207_
rlabel metal1 28704 21590 28704 21590 0 _0208_
rlabel metal1 29026 20026 29026 20026 0 _0209_
rlabel metal1 32614 25228 32614 25228 0 _0210_
rlabel metal1 30682 12172 30682 12172 0 _0211_
rlabel metal2 33994 25058 33994 25058 0 _0212_
rlabel metal1 13754 24854 13754 24854 0 _0213_
rlabel metal2 30498 29308 30498 29308 0 _0214_
rlabel metal1 29854 27642 29854 27642 0 _0215_
rlabel metal2 34086 29818 34086 29818 0 _0216_
rlabel metal1 32430 28934 32430 28934 0 _0217_
rlabel metal1 33718 29070 33718 29070 0 _0218_
rlabel metal1 34776 28050 34776 28050 0 _0219_
rlabel metal1 22218 19822 22218 19822 0 _0220_
rlabel metal1 30360 12206 30360 12206 0 _0221_
rlabel metal1 31096 25262 31096 25262 0 _0222_
rlabel metal1 32430 25296 32430 25296 0 _0223_
rlabel metal2 33258 23290 33258 23290 0 _0224_
rlabel metal1 29992 21114 29992 21114 0 _0225_
rlabel metal1 28934 19856 28934 19856 0 _0226_
rlabel metal1 29394 17646 29394 17646 0 _0227_
rlabel metal1 28934 15436 28934 15436 0 _0228_
rlabel metal1 31142 14416 31142 14416 0 _0229_
rlabel metal1 28428 12410 28428 12410 0 _0230_
rlabel metal2 30222 13158 30222 13158 0 _0231_
rlabel metal1 6486 25228 6486 25228 0 _0232_
rlabel metal1 36616 13498 36616 13498 0 _0233_
rlabel metal1 37812 15130 37812 15130 0 _0234_
rlabel metal2 42274 16252 42274 16252 0 _0235_
rlabel metal1 36064 12614 36064 12614 0 _0236_
rlabel metal1 36754 12682 36754 12682 0 _0237_
rlabel metal1 35558 12920 35558 12920 0 _0238_
rlabel metal2 43286 15266 43286 15266 0 _0239_
rlabel metal1 41101 21930 41101 21930 0 _0240_
rlabel metal1 44712 15402 44712 15402 0 _0241_
rlabel metal1 44574 14858 44574 14858 0 _0242_
rlabel metal1 43792 14994 43792 14994 0 _0243_
rlabel metal2 44666 15776 44666 15776 0 _0244_
rlabel metal2 40986 20604 40986 20604 0 _0245_
rlabel metal2 45402 15844 45402 15844 0 _0246_
rlabel metal1 45678 16184 45678 16184 0 _0247_
rlabel metal2 44298 17816 44298 17816 0 _0248_
rlabel metal2 45494 17952 45494 17952 0 _0249_
rlabel metal2 44298 19074 44298 19074 0 _0250_
rlabel metal1 43976 18734 43976 18734 0 _0251_
rlabel metal2 43930 18156 43930 18156 0 _0252_
rlabel metal2 44390 18870 44390 18870 0 _0253_
rlabel metal2 45402 18292 45402 18292 0 _0254_
rlabel metal1 44160 19890 44160 19890 0 _0255_
rlabel metal1 44071 19482 44071 19482 0 _0256_
rlabel metal2 44114 20230 44114 20230 0 _0257_
rlabel metal1 41400 17170 41400 17170 0 _0258_
rlabel via1 44198 15402 44198 15402 0 _0259_
rlabel metal2 43286 16116 43286 16116 0 _0260_
rlabel metal1 41331 17034 41331 17034 0 _0261_
rlabel metal1 40756 17170 40756 17170 0 _0262_
rlabel metal1 40204 16558 40204 16558 0 _0263_
rlabel metal2 41814 16796 41814 16796 0 _0264_
rlabel metal1 40572 14994 40572 14994 0 _0265_
rlabel metal1 40388 15606 40388 15606 0 _0266_
rlabel metal2 40894 14382 40894 14382 0 _0267_
rlabel metal2 40802 19108 40802 19108 0 _0268_
rlabel metal1 39376 19822 39376 19822 0 _0269_
rlabel metal2 40250 18496 40250 18496 0 _0270_
rlabel metal1 40296 17646 40296 17646 0 _0271_
rlabel metal2 40066 18530 40066 18530 0 _0272_
rlabel metal2 40434 18904 40434 18904 0 _0273_
rlabel metal1 39790 19278 39790 19278 0 _0274_
rlabel metal2 41354 19669 41354 19669 0 _0275_
rlabel metal1 40250 19924 40250 19924 0 _0276_
rlabel metal1 40342 19856 40342 19856 0 _0277_
rlabel metal2 41262 18938 41262 18938 0 _0278_
rlabel metal2 42918 20162 42918 20162 0 _0279_
rlabel metal2 41354 17850 41354 17850 0 _0280_
rlabel metal1 41906 16592 41906 16592 0 _0281_
rlabel metal2 42826 18870 42826 18870 0 _0282_
rlabel metal1 42504 22474 42504 22474 0 _0283_
rlabel metal2 43470 22610 43470 22610 0 _0284_
rlabel metal2 43654 21692 43654 21692 0 _0285_
rlabel metal2 44206 22440 44206 22440 0 _0286_
rlabel metal1 42734 21658 42734 21658 0 _0287_
rlabel metal1 43378 24140 43378 24140 0 _0288_
rlabel metal1 44737 25126 44737 25126 0 _0289_
rlabel metal2 41814 25092 41814 25092 0 _0290_
rlabel metal2 43102 25636 43102 25636 0 _0291_
rlabel metal2 44206 24378 44206 24378 0 _0292_
rlabel metal2 44298 23868 44298 23868 0 _0293_
rlabel metal2 45218 25670 45218 25670 0 _0294_
rlabel metal1 43930 26010 43930 26010 0 _0295_
rlabel metal1 43470 27982 43470 27982 0 _0296_
rlabel metal1 43654 29682 43654 29682 0 _0297_
rlabel metal2 43930 29818 43930 29818 0 _0298_
rlabel metal1 44436 29818 44436 29818 0 _0299_
rlabel metal2 44206 30498 44206 30498 0 _0300_
rlabel metal1 42780 30702 42780 30702 0 _0301_
rlabel metal2 43746 29852 43746 29852 0 _0302_
rlabel metal1 44068 27370 44068 27370 0 _0303_
rlabel metal2 43378 28220 43378 28220 0 _0304_
rlabel metal1 43930 28186 43930 28186 0 _0305_
rlabel metal2 42826 28356 42826 28356 0 _0306_
rlabel metal1 19918 23052 19918 23052 0 _0307_
rlabel metal1 17940 29682 17940 29682 0 _0308_
rlabel metal2 16882 28934 16882 28934 0 _0309_
rlabel metal2 15502 29750 15502 29750 0 _0310_
rlabel metal1 11868 28458 11868 28458 0 _0311_
rlabel metal2 17066 31416 17066 31416 0 _0312_
rlabel metal1 15916 30702 15916 30702 0 _0313_
rlabel metal2 17526 30464 17526 30464 0 _0314_
rlabel metal1 18078 31280 18078 31280 0 _0315_
rlabel metal1 14766 31926 14766 31926 0 _0316_
rlabel metal2 14306 32436 14306 32436 0 _0317_
rlabel metal2 12190 32504 12190 32504 0 _0318_
rlabel metal1 12190 32538 12190 32538 0 _0319_
rlabel metal1 13754 28424 13754 28424 0 _0320_
rlabel metal1 13846 28730 13846 28730 0 _0321_
rlabel metal2 13018 24582 13018 24582 0 _0322_
rlabel metal1 12788 24174 12788 24174 0 _0323_
rlabel metal2 11638 22542 11638 22542 0 _0324_
rlabel metal1 11224 22610 11224 22610 0 _0325_
rlabel metal1 12052 25194 12052 25194 0 _0326_
rlabel metal1 11868 25466 11868 25466 0 _0327_
rlabel metal2 12190 28152 12190 28152 0 _0328_
rlabel metal1 12742 28560 12742 28560 0 _0329_
rlabel metal1 27646 21556 27646 21556 0 _0330_
rlabel metal1 27324 24378 27324 24378 0 _0331_
rlabel metal2 26450 21692 26450 21692 0 _0332_
rlabel metal2 21298 17680 21298 17680 0 _0333_
rlabel metal2 20102 24276 20102 24276 0 _0334_
rlabel metal2 27186 25262 27186 25262 0 _0335_
rlabel metal1 29026 24276 29026 24276 0 _0336_
rlabel metal1 29072 21998 29072 21998 0 _0337_
rlabel metal2 31602 11084 31602 11084 0 _0338_
rlabel metal1 39790 33966 39790 33966 0 _0339_
rlabel metal2 28106 21386 28106 21386 0 _0340_
rlabel metal1 30866 11696 30866 11696 0 _0341_
rlabel metal1 38134 34034 38134 34034 0 _0342_
rlabel metal2 39238 34612 39238 34612 0 _0343_
rlabel metal1 29946 34578 29946 34578 0 _0344_
rlabel metal1 30360 33626 30360 33626 0 _0345_
rlabel metal1 37628 34170 37628 34170 0 _0346_
rlabel metal1 32936 35054 32936 35054 0 _0347_
rlabel metal2 38962 34442 38962 34442 0 _0348_
rlabel metal1 40388 32538 40388 32538 0 _0349_
rlabel metal2 38870 24310 38870 24310 0 _0350_
rlabel metal1 32982 26010 32982 26010 0 _0351_
rlabel metal1 34914 23086 34914 23086 0 _0352_
rlabel metal2 31326 22780 31326 22780 0 _0353_
rlabel metal1 31096 11730 31096 11730 0 _0354_
rlabel metal1 30820 18394 30820 18394 0 _0355_
rlabel metal1 30774 16762 30774 16762 0 _0356_
rlabel metal1 31372 15130 31372 15130 0 _0357_
rlabel metal1 31970 13294 31970 13294 0 _0358_
rlabel metal2 29762 10812 29762 10812 0 _0359_
rlabel metal1 31924 11730 31924 11730 0 _0360_
rlabel metal1 26542 23800 26542 23800 0 _0361_
rlabel metal1 26220 11288 26220 11288 0 _0362_
rlabel metal1 14858 23086 14858 23086 0 _0363_
rlabel metal1 25530 10166 25530 10166 0 _0364_
rlabel metal1 14904 24174 14904 24174 0 _0365_
rlabel metal1 25392 27098 25392 27098 0 _0366_
rlabel metal2 27830 27574 27830 27574 0 _0367_
rlabel metal1 24702 22202 24702 22202 0 _0368_
rlabel metal1 23598 26384 23598 26384 0 _0369_
rlabel metal2 20286 23936 20286 23936 0 _0370_
rlabel metal2 14582 26996 14582 26996 0 _0371_
rlabel metal2 14490 23562 14490 23562 0 _0372_
rlabel metal1 14398 21114 14398 21114 0 _0373_
rlabel metal1 12696 19482 12696 19482 0 _0374_
rlabel metal1 12742 18258 12742 18258 0 _0375_
rlabel metal1 12742 17544 12742 17544 0 _0376_
rlabel metal2 27370 19516 27370 19516 0 _0377_
rlabel metal2 25806 14518 25806 14518 0 _0378_
rlabel metal1 18124 14586 18124 14586 0 _0379_
rlabel metal1 17664 12818 17664 12818 0 _0380_
rlabel metal2 19826 24106 19826 24106 0 _0381_
rlabel metal1 18124 10234 18124 10234 0 _0382_
rlabel metal1 26496 10234 26496 10234 0 _0383_
rlabel metal1 27692 20910 27692 20910 0 _0384_
rlabel metal1 26588 12410 26588 12410 0 _0385_
rlabel metal1 20194 24582 20194 24582 0 _0386_
rlabel metal1 22540 27642 22540 27642 0 _0387_
rlabel metal2 22126 29682 22126 29682 0 _0388_
rlabel metal1 23966 21114 23966 21114 0 _0389_
rlabel metal2 20286 28220 20286 28220 0 _0390_
rlabel metal1 19642 28560 19642 28560 0 _0391_
rlabel metal2 19642 24582 19642 24582 0 _0392_
rlabel metal1 20562 22066 20562 22066 0 _0393_
rlabel metal1 19596 20026 19596 20026 0 _0394_
rlabel metal2 22218 19516 22218 19516 0 _0395_
rlabel metal2 20010 18870 20010 18870 0 _0396_
rlabel metal1 28152 18394 28152 18394 0 _0397_
rlabel metal1 26772 16082 26772 16082 0 _0398_
rlabel metal1 20562 17306 20562 17306 0 _0399_
rlabel metal1 21068 13498 21068 13498 0 _0400_
rlabel metal1 23368 12954 23368 12954 0 _0401_
rlabel metal1 26404 12206 26404 12206 0 _0402_
rlabel metal1 5566 36108 5566 36108 0 _0403_
rlabel metal1 9936 36142 9936 36142 0 _0404_
rlabel metal1 8740 37230 8740 37230 0 _0405_
rlabel metal1 6256 37366 6256 37366 0 _0406_
rlabel metal1 5014 36346 5014 36346 0 _0407_
rlabel metal1 5934 35802 5934 35802 0 _0408_
rlabel metal1 5704 33626 5704 33626 0 _0409_
rlabel metal1 5290 34612 5290 34612 0 _0410_
rlabel metal1 9752 33626 9752 33626 0 _0411_
rlabel metal1 7544 33014 7544 33014 0 _0412_
rlabel metal2 7038 34170 7038 34170 0 _0413_
rlabel metal1 2392 44846 2392 44846 0 _0414_
rlabel metal2 24886 4318 24886 4318 0 _0415_
rlabel metal1 6348 41106 6348 41106 0 _0416_
rlabel metal2 2530 6052 2530 6052 0 _0417_
rlabel metal1 41124 45458 41124 45458 0 _0418_
rlabel metal1 4876 4114 4876 4114 0 _0419_
rlabel metal1 4876 3502 4876 3502 0 _0420_
rlabel metal2 2622 23698 2622 23698 0 _0421_
rlabel metal1 4186 4556 4186 4556 0 _0422_
rlabel metal1 19918 24752 19918 24752 0 _0423_
rlabel metal1 3818 10642 3818 10642 0 _0424_
rlabel metal1 6256 4114 6256 4114 0 _0425_
rlabel metal1 8740 27574 8740 27574 0 _0426_
rlabel metal2 10258 28458 10258 28458 0 _0427_
rlabel metal2 9982 27030 9982 27030 0 _0428_
rlabel metal2 10626 27778 10626 27778 0 _0429_
rlabel metal1 11868 28186 11868 28186 0 _0430_
rlabel metal1 9706 25364 9706 25364 0 _0431_
rlabel metal2 13110 29988 13110 29988 0 _0432_
rlabel metal1 12880 31314 12880 31314 0 _0433_
rlabel metal2 11730 30838 11730 30838 0 _0434_
rlabel metal2 11086 32198 11086 32198 0 _0435_
rlabel metal1 8602 30736 8602 30736 0 _0436_
rlabel metal2 9154 28220 9154 28220 0 _0437_
rlabel metal2 11178 24378 11178 24378 0 _0438_
rlabel metal1 9384 23698 9384 23698 0 _0439_
rlabel metal1 7774 25262 7774 25262 0 _0440_
rlabel metal1 6302 26962 6302 26962 0 _0441_
rlabel metal2 7130 33354 7130 33354 0 _0442_
rlabel metal1 7084 27982 7084 27982 0 _0443_
rlabel metal1 29992 30158 29992 30158 0 _0444_
rlabel metal1 30084 30362 30084 30362 0 _0445_
rlabel metal1 34270 32300 34270 32300 0 _0446_
rlabel metal1 35052 32334 35052 32334 0 _0447_
rlabel metal1 29440 30702 29440 30702 0 _0448_
rlabel metal1 31602 24140 31602 24140 0 _0449_
rlabel metal1 33350 12818 33350 12818 0 _0450_
rlabel metal1 33074 19414 33074 19414 0 _0451_
rlabel metal2 31786 32096 31786 32096 0 _0452_
rlabel metal1 31234 31926 31234 31926 0 _0453_
rlabel metal1 33488 31790 33488 31790 0 _0454_
rlabel metal2 31602 31484 31602 31484 0 _0455_
rlabel metal2 33074 29818 33074 29818 0 _0456_
rlabel metal1 33718 12954 33718 12954 0 _0457_
rlabel metal1 33442 21454 33442 21454 0 _0458_
rlabel metal2 33074 32572 33074 32572 0 _0459_
rlabel metal2 36386 32640 36386 32640 0 _0460_
rlabel metal2 36018 34884 36018 34884 0 _0461_
rlabel metal1 36800 34034 36800 34034 0 _0462_
rlabel metal1 36340 34170 36340 34170 0 _0463_
rlabel metal1 35926 31382 35926 31382 0 _0464_
rlabel metal1 35512 32742 35512 32742 0 _0465_
rlabel metal1 35880 32402 35880 32402 0 _0466_
rlabel metal1 35098 34986 35098 34986 0 _0467_
rlabel metal1 35006 33966 35006 33966 0 _0468_
rlabel metal2 35466 34782 35466 34782 0 _0469_
rlabel metal2 36570 33626 36570 33626 0 _0470_
rlabel metal1 34362 32538 34362 32538 0 _0471_
rlabel metal2 33626 32640 33626 32640 0 _0472_
rlabel metal1 33028 33082 33028 33082 0 _0473_
rlabel metal2 38962 32309 38962 32309 0 _0474_
rlabel metal1 39054 31994 39054 31994 0 _0475_
rlabel metal2 37858 32028 37858 32028 0 _0476_
rlabel metal1 35374 34000 35374 34000 0 _0477_
rlabel metal1 37536 33830 37536 33830 0 _0478_
rlabel metal1 37720 31790 37720 31790 0 _0479_
rlabel metal1 37030 30906 37030 30906 0 _0480_
rlabel metal1 39790 29478 39790 29478 0 _0481_
rlabel metal1 40066 30158 40066 30158 0 _0482_
rlabel metal2 40710 29716 40710 29716 0 _0483_
rlabel metal1 39100 28934 39100 28934 0 _0484_
rlabel metal1 37950 28118 37950 28118 0 _0485_
rlabel metal1 39284 30158 39284 30158 0 _0486_
rlabel metal1 38916 29614 38916 29614 0 _0487_
rlabel metal1 38456 29614 38456 29614 0 _0488_
rlabel metal1 39284 27302 39284 27302 0 _0489_
rlabel metal1 40158 27438 40158 27438 0 _0490_
rlabel metal1 40388 26010 40388 26010 0 _0491_
rlabel metal2 40342 26724 40342 26724 0 _0492_
rlabel metal1 39744 25874 39744 25874 0 _0493_
rlabel metal1 37812 27098 37812 27098 0 _0494_
rlabel metal2 38410 28322 38410 28322 0 _0495_
rlabel metal1 37122 26384 37122 26384 0 _0496_
rlabel metal1 37030 26486 37030 26486 0 _0497_
rlabel metal1 36524 26554 36524 26554 0 _0498_
rlabel metal1 35880 26010 35880 26010 0 _0499_
rlabel metal2 35466 26486 35466 26486 0 _0500_
rlabel metal2 39928 19346 39928 19346 0 _0501_
rlabel metal2 38318 21828 38318 21828 0 _0502_
rlabel metal1 39192 28526 39192 28526 0 _0503_
rlabel metal2 38318 28866 38318 28866 0 _0504_
rlabel metal1 39422 28560 39422 28560 0 _0505_
rlabel metal1 38640 29138 38640 29138 0 _0506_
rlabel metal1 38502 22032 38502 22032 0 _0507_
rlabel metal1 36984 21998 36984 21998 0 _0508_
rlabel metal1 36708 21522 36708 21522 0 _0509_
rlabel metal1 37674 22644 37674 22644 0 _0510_
rlabel metal2 37398 21488 37398 21488 0 _0511_
rlabel metal1 37812 22202 37812 22202 0 _0512_
rlabel metal2 37674 23494 37674 23494 0 _0513_
rlabel metal2 35558 21692 35558 21692 0 _0514_
rlabel metal1 35236 20434 35236 20434 0 _0515_
rlabel metal2 35282 21828 35282 21828 0 _0516_
rlabel metal2 35650 21284 35650 21284 0 _0517_
rlabel metal1 32798 21454 32798 21454 0 _0518_
rlabel metal1 32200 21522 32200 21522 0 _0519_
rlabel metal1 34776 20230 34776 20230 0 _0520_
rlabel metal2 33718 19788 33718 19788 0 _0521_
rlabel metal2 33810 20094 33810 20094 0 _0522_
rlabel metal2 33902 20026 33902 20026 0 _0523_
rlabel metal1 33074 19346 33074 19346 0 _0524_
rlabel metal2 40710 14076 40710 14076 0 _0525_
rlabel metal1 34454 17170 34454 17170 0 _0526_
rlabel metal1 35328 17850 35328 17850 0 _0527_
rlabel metal1 35328 18734 35328 18734 0 _0528_
rlabel metal1 34960 18802 34960 18802 0 _0529_
rlabel metal1 35972 18734 35972 18734 0 _0530_
rlabel metal2 36570 18462 36570 18462 0 _0531_
rlabel metal1 36524 17850 36524 17850 0 _0532_
rlabel metal1 36294 20434 36294 20434 0 _0533_
rlabel metal2 36938 21318 36938 21318 0 _0534_
rlabel metal2 37582 18768 37582 18768 0 _0535_
rlabel metal2 36018 20774 36018 20774 0 _0536_
rlabel metal1 35742 18088 35742 18088 0 _0537_
rlabel metal1 35328 18326 35328 18326 0 _0538_
rlabel metal2 36110 17306 36110 17306 0 _0539_
rlabel metal2 36478 15980 36478 15980 0 _0540_
rlabel metal2 36846 14076 36846 14076 0 _0541_
rlabel metal2 36386 15708 36386 15708 0 _0542_
rlabel metal1 37168 14926 37168 14926 0 _0543_
rlabel metal1 38088 15470 38088 15470 0 _0544_
rlabel metal1 34362 15436 34362 15436 0 _0545_
rlabel metal1 35834 14994 35834 14994 0 _0546_
rlabel metal1 34546 14586 34546 14586 0 _0547_
rlabel metal2 35006 14212 35006 14212 0 _0548_
rlabel metal1 35558 14892 35558 14892 0 _0549_
rlabel metal1 33166 14416 33166 14416 0 _0550_
rlabel metal2 33350 14858 33350 14858 0 _0551_
rlabel metal2 36386 13158 36386 13158 0 _0552_
rlabel metal1 36800 11118 36800 11118 0 _0553_
rlabel metal2 35558 11526 35558 11526 0 _0554_
rlabel metal1 36524 12818 36524 12818 0 _0555_
rlabel metal2 37674 13804 37674 13804 0 _0556_
rlabel metal2 36754 13124 36754 13124 0 _0557_
rlabel metal1 37950 12410 37950 12410 0 _0558_
rlabel metal1 34776 12818 34776 12818 0 _0559_
rlabel metal1 35098 12784 35098 12784 0 _0560_
rlabel metal1 35282 12614 35282 12614 0 _0561_
rlabel metal2 35374 11900 35374 11900 0 _0562_
rlabel metal1 35190 12240 35190 12240 0 _0563_
rlabel metal1 34684 12070 34684 12070 0 _0564_
rlabel metal2 33534 11900 33534 11900 0 _0565_
rlabel metal1 24150 15674 24150 15674 0 _0566_
rlabel metal2 23966 17850 23966 17850 0 _0567_
rlabel metal1 23782 15436 23782 15436 0 _0568_
rlabel metal2 23322 16082 23322 16082 0 _0569_
rlabel metal2 23782 18122 23782 18122 0 _0570_
rlabel metal1 22954 17612 22954 17612 0 _0571_
rlabel metal1 23092 16762 23092 16762 0 _0572_
rlabel metal1 14582 15504 14582 15504 0 _0573_
rlabel metal1 14582 16116 14582 16116 0 _0574_
rlabel metal1 14490 15674 14490 15674 0 _0575_
rlabel metal1 16146 16048 16146 16048 0 _0576_
rlabel metal2 20838 15674 20838 15674 0 _0577_
rlabel metal2 19550 25602 19550 25602 0 _0578_
rlabel metal2 23598 24310 23598 24310 0 _0579_
rlabel metal1 25576 29138 25576 29138 0 _0580_
rlabel metal2 25438 29852 25438 29852 0 _0581_
rlabel metal1 23828 25330 23828 25330 0 _0582_
rlabel metal2 23138 24276 23138 24276 0 _0583_
rlabel metal2 20654 25092 20654 25092 0 _0584_
rlabel metal1 17848 25874 17848 25874 0 _0585_
rlabel metal2 18630 25568 18630 25568 0 _0586_
rlabel metal1 20148 25874 20148 25874 0 _0587_
rlabel metal1 17894 24752 17894 24752 0 _0588_
rlabel metal1 17250 24378 17250 24378 0 _0589_
rlabel metal2 17894 25092 17894 25092 0 _0590_
rlabel metal2 18170 23603 18170 23603 0 _0591_
rlabel metal1 17043 19346 17043 19346 0 _0592_
rlabel metal1 18032 20434 18032 20434 0 _0593_
rlabel metal2 17342 24888 17342 24888 0 _0594_
rlabel metal1 18170 24582 18170 24582 0 _0595_
rlabel metal1 16422 18666 16422 18666 0 _0596_
rlabel metal2 16698 18530 16698 18530 0 _0597_
rlabel metal1 16928 22406 16928 22406 0 _0598_
rlabel metal1 16422 17680 16422 17680 0 _0599_
rlabel metal1 15364 15470 15364 15470 0 _0600_
rlabel metal2 15134 17476 15134 17476 0 _0601_
rlabel metal1 15824 17850 15824 17850 0 _0602_
rlabel metal1 16698 16762 16698 16762 0 _0603_
rlabel metal2 21022 16252 21022 16252 0 _0604_
rlabel metal1 19504 14042 19504 14042 0 _0605_
rlabel metal2 20194 14790 20194 14790 0 _0606_
rlabel metal1 20386 15130 20386 15130 0 _0607_
rlabel metal1 22126 11832 22126 11832 0 _0608_
rlabel metal1 23874 9520 23874 9520 0 _0609_
rlabel metal1 22908 9894 22908 9894 0 _0610_
rlabel metal1 23782 10030 23782 10030 0 _0611_
rlabel metal2 22218 9996 22218 9996 0 _0612_
rlabel metal1 21758 9554 21758 9554 0 _0613_
rlabel metal1 22494 11118 22494 11118 0 _0614_
rlabel metal1 23138 10710 23138 10710 0 _0615_
rlabel metal2 18998 11934 18998 11934 0 _0616_
rlabel metal1 18768 11594 18768 11594 0 _0617_
rlabel metal1 21206 11764 21206 11764 0 _0618_
rlabel viali 22126 10642 22126 10642 0 _0619_
rlabel metal2 21850 10438 21850 10438 0 _0620_
rlabel metal1 22632 10778 22632 10778 0 _0621_
rlabel metal2 20838 34850 20838 34850 0 _0622_
rlabel metal1 19550 37842 19550 37842 0 _0623_
rlabel metal1 20700 33082 20700 33082 0 _0624_
rlabel metal1 21206 32946 21206 32946 0 _0625_
rlabel metal2 21206 33762 21206 33762 0 _0626_
rlabel metal1 22126 31892 22126 31892 0 _0627_
rlabel metal1 25530 25874 25530 25874 0 _0628_
rlabel metal1 24794 32368 24794 32368 0 _0629_
rlabel metal2 25070 32096 25070 32096 0 _0630_
rlabel metal1 25438 36720 25438 36720 0 _0631_
rlabel metal2 22218 32266 22218 32266 0 _0632_
rlabel metal1 23506 10132 23506 10132 0 _0633_
rlabel metal1 23874 38828 23874 38828 0 _0634_
rlabel metal1 17664 27506 17664 27506 0 _0635_
rlabel metal1 20608 32402 20608 32402 0 _0636_
rlabel metal1 20608 31382 20608 31382 0 _0637_
rlabel metal1 20194 32198 20194 32198 0 _0638_
rlabel metal2 18722 33592 18722 33592 0 _0639_
rlabel metal1 23414 40018 23414 40018 0 _0640_
rlabel metal2 18814 33796 18814 33796 0 _0641_
rlabel metal2 17250 32844 17250 32844 0 _0642_
rlabel metal2 18170 32844 18170 32844 0 _0643_
rlabel metal1 18400 33490 18400 33490 0 _0644_
rlabel metal2 17526 34306 17526 34306 0 _0645_
rlabel metal1 17434 34000 17434 34000 0 _0646_
rlabel metal1 25773 33490 25773 33490 0 _0647_
rlabel metal2 17710 34238 17710 34238 0 _0648_
rlabel metal1 16698 34510 16698 34510 0 _0649_
rlabel metal1 24012 39406 24012 39406 0 _0650_
rlabel metal2 17158 34748 17158 34748 0 _0651_
rlabel metal2 27554 33082 27554 33082 0 _0652_
rlabel metal1 27784 33626 27784 33626 0 _0653_
rlabel metal1 25990 34986 25990 34986 0 _0654_
rlabel metal1 18814 33524 18814 33524 0 _0655_
rlabel metal1 22126 34476 22126 34476 0 _0656_
rlabel metal2 22034 34238 22034 34238 0 _0657_
rlabel metal2 23506 34340 23506 34340 0 _0658_
rlabel metal2 25622 33694 25622 33694 0 _0659_
rlabel metal1 25622 33422 25622 33422 0 _0660_
rlabel metal1 27738 35122 27738 35122 0 _0661_
rlabel metal2 27646 34646 27646 34646 0 _0662_
rlabel metal1 27416 35258 27416 35258 0 _0663_
rlabel metal1 24702 36720 24702 36720 0 _0664_
rlabel metal1 25392 36142 25392 36142 0 _0665_
rlabel metal2 26174 35394 26174 35394 0 _0666_
rlabel metal1 26450 36346 26450 36346 0 _0667_
rlabel via1 26550 36006 26550 36006 0 _0668_
rlabel metal1 26726 36312 26726 36312 0 _0669_
rlabel metal1 25208 36822 25208 36822 0 _0670_
rlabel metal2 28198 37060 28198 37060 0 _0671_
rlabel metal2 24794 35054 24794 35054 0 _0672_
rlabel metal1 25530 35530 25530 35530 0 _0673_
rlabel metal1 24334 36550 24334 36550 0 _0674_
rlabel metal1 23828 34578 23828 34578 0 _0675_
rlabel metal2 21758 36516 21758 36516 0 _0676_
rlabel metal2 25806 35496 25806 35496 0 _0677_
rlabel metal2 21482 35292 21482 35292 0 _0678_
rlabel metal1 23782 35020 23782 35020 0 _0679_
rlabel metal2 21574 35700 21574 35700 0 _0680_
rlabel metal2 19550 36550 19550 36550 0 _0681_
rlabel metal1 20056 37638 20056 37638 0 _0682_
rlabel metal1 19918 36720 19918 36720 0 _0683_
rlabel metal1 18860 37298 18860 37298 0 _0684_
rlabel metal2 18630 37502 18630 37502 0 _0685_
rlabel metal1 17986 37910 17986 37910 0 _0686_
rlabel metal2 18262 37638 18262 37638 0 _0687_
rlabel metal2 22310 37196 22310 37196 0 _0688_
rlabel metal1 22172 38930 22172 38930 0 _0689_
rlabel metal1 22034 38896 22034 38896 0 _0690_
rlabel metal1 24242 39610 24242 39610 0 _0691_
rlabel via1 23690 40477 23690 40477 0 _0692_
rlabel metal1 22264 39950 22264 39950 0 _0693_
rlabel metal2 23598 38556 23598 38556 0 _0694_
rlabel metal2 24426 39542 24426 39542 0 _0695_
rlabel metal2 23690 39610 23690 39610 0 _0696_
rlabel metal2 23506 38692 23506 38692 0 _0697_
rlabel metal2 23598 39100 23598 39100 0 _0698_
rlabel metal1 22356 38522 22356 38522 0 _0699_
rlabel metal2 23046 39678 23046 39678 0 _0700_
rlabel metal2 16054 39202 16054 39202 0 _0701_
rlabel metal1 13800 37298 13800 37298 0 _0702_
rlabel metal1 13570 37196 13570 37196 0 _0703_
rlabel metal1 13064 37230 13064 37230 0 _0704_
rlabel metal1 14444 37978 14444 37978 0 _0705_
rlabel metal1 13386 37842 13386 37842 0 _0706_
rlabel metal1 14950 38318 14950 38318 0 _0707_
rlabel metal1 15502 37842 15502 37842 0 _0708_
rlabel metal2 15962 36788 15962 36788 0 _0709_
rlabel metal1 14306 34170 14306 34170 0 _0710_
rlabel metal2 14582 36482 14582 36482 0 _0711_
rlabel metal2 4830 38080 4830 38080 0 _0712_
rlabel metal2 24426 28900 24426 28900 0 _0713_
rlabel metal2 23782 28798 23782 28798 0 _0714_
rlabel metal1 23460 12274 23460 12274 0 _0715_
rlabel metal1 23414 28730 23414 28730 0 _0716_
rlabel metal2 25622 30158 25622 30158 0 _0717_
rlabel metal2 25438 30906 25438 30906 0 _0718_
rlabel metal1 23874 23834 23874 23834 0 _0719_
rlabel metal2 23690 21971 23690 21971 0 _0720_
rlabel metal1 22954 22202 22954 22202 0 _0721_
rlabel metal1 22862 22950 22862 22950 0 _0722_
rlabel metal1 20102 25330 20102 25330 0 _0723_
rlabel metal1 21114 26894 21114 26894 0 _0724_
rlabel metal2 20838 26554 20838 26554 0 _0725_
rlabel metal1 20148 26350 20148 26350 0 _0726_
rlabel metal1 18308 25738 18308 25738 0 _0727_
rlabel metal1 17710 26418 17710 26418 0 _0728_
rlabel metal1 17756 27098 17756 27098 0 _0729_
rlabel metal1 17986 27506 17986 27506 0 _0730_
rlabel metal1 17020 26214 17020 26214 0 _0731_
rlabel metal1 17664 24242 17664 24242 0 _0732_
rlabel metal1 17342 24072 17342 24072 0 _0733_
rlabel metal1 15502 24072 15502 24072 0 _0734_
rlabel metal1 17112 21590 17112 21590 0 _0735_
rlabel metal1 17158 21420 17158 21420 0 _0736_
rlabel metal1 17204 21046 17204 21046 0 _0737_
rlabel metal1 17894 21862 17894 21862 0 _0738_
rlabel metal1 16974 19482 16974 19482 0 _0739_
rlabel metal1 17526 20026 17526 20026 0 _0740_
rlabel metal1 15962 20366 15962 20366 0 _0741_
rlabel metal1 16054 20400 16054 20400 0 _0742_
rlabel metal1 15410 19482 15410 19482 0 _0743_
rlabel metal2 14674 19958 14674 19958 0 _0744_
rlabel metal1 16284 17850 16284 17850 0 _0745_
rlabel metal1 16422 16626 16422 16626 0 _0746_
rlabel metal1 16698 16592 16698 16592 0 _0747_
rlabel metal1 17480 16694 17480 16694 0 _0748_
rlabel metal2 18354 17612 18354 17612 0 _0749_
rlabel metal1 16376 15538 16376 15538 0 _0750_
rlabel metal2 7682 3502 7682 3502 0 _0751_
rlabel metal2 3082 43520 3082 43520 0 _0752_
rlabel metal1 19642 3094 19642 3094 0 _0753_
rlabel metal2 2898 9316 2898 9316 0 _0754_
rlabel metal2 47886 3604 47886 3604 0 _0755_
rlabel metal2 3542 3774 3542 3774 0 _0756_
rlabel metal1 46690 19924 46690 19924 0 _0757_
rlabel metal2 6946 29410 6946 29410 0 _0758_
rlabel metal2 46046 32028 46046 32028 0 _0759_
rlabel metal2 45586 32606 45586 32606 0 _0760_
rlabel metal2 46690 26588 46690 26588 0 _0761_
rlabel metal2 22034 24412 22034 24412 0 _0762_
rlabel metal2 16054 40290 16054 40290 0 _0763_
rlabel metal1 13938 39610 13938 39610 0 _0764_
rlabel metal2 17802 40222 17802 40222 0 _0765_
rlabel metal2 6946 28798 6946 28798 0 _0766_
rlabel metal2 47886 23970 47886 23970 0 _0767_
rlabel metal1 48024 35802 48024 35802 0 _0768_
rlabel metal2 5934 43554 5934 43554 0 _0769_
rlabel metal1 46782 24786 46782 24786 0 _0770_
rlabel metal2 3266 10268 3266 10268 0 _0771_
rlabel metal1 47288 42602 47288 42602 0 _0772_
rlabel metal2 29946 45696 29946 45696 0 _0773_
rlabel metal1 12328 2346 12328 2346 0 _0774_
rlabel metal1 46920 18802 46920 18802 0 _0775_
rlabel metal1 3266 3604 3266 3604 0 _0776_
rlabel metal2 48162 5372 48162 5372 0 _0777_
rlabel metal1 5382 45526 5382 45526 0 _0778_
rlabel metal2 45402 4012 45402 4012 0 _0779_
rlabel metal2 6118 3740 6118 3740 0 _0780_
rlabel metal1 46598 12614 46598 12614 0 _0781_
rlabel metal1 47104 45526 47104 45526 0 _0782_
rlabel metal1 39100 45798 39100 45798 0 _0783_
rlabel metal2 33258 46308 33258 46308 0 _0784_
rlabel metal2 6854 3196 6854 3196 0 _0785_
rlabel metal1 2346 42874 2346 42874 0 _0786_
rlabel metal1 47288 29682 47288 29682 0 _0787_
rlabel metal2 22678 46308 22678 46308 0 _0788_
rlabel metal2 46690 46172 46690 46172 0 _0789_
rlabel metal2 2438 20196 2438 20196 0 _0790_
rlabel metal1 19918 2346 19918 2346 0 _0791_
rlabel metal2 5106 14756 5106 14756 0 _0792_
rlabel metal2 48162 27676 48162 27676 0 _0793_
rlabel metal1 3266 2312 3266 2312 0 _0794_
rlabel metal2 2898 7650 2898 7650 0 _0795_
rlabel metal2 38226 3842 38226 3842 0 _0796_
rlabel metal2 47150 40222 47150 40222 0 _0797_
rlabel metal1 6900 41242 6900 41242 0 _0798_
rlabel metal2 48162 26044 48162 26044 0 _0799_
rlabel metal2 45954 46308 45954 46308 0 _0800_
rlabel metal2 46322 6188 46322 6188 0 _0801_
rlabel metal2 6670 23970 6670 23970 0 _0802_
rlabel metal1 40388 45050 40388 45050 0 _0803_
rlabel metal1 6348 31382 6348 31382 0 _0804_
rlabel metal2 32430 6562 32430 6562 0 _0805_
rlabel metal2 47886 21794 47886 21794 0 _0806_
rlabel metal2 27370 3502 27370 3502 0 _0807_
rlabel metal1 36984 45526 36984 45526 0 _0808_
rlabel metal1 3680 5610 3680 5610 0 _0809_
rlabel metal1 39192 46138 39192 46138 0 _0810_
rlabel metal2 17066 3230 17066 3230 0 _0811_
rlabel metal2 45126 3774 45126 3774 0 _0812_
rlabel metal2 2438 6562 2438 6562 0 _0813_
rlabel metal2 2438 14178 2438 14178 0 _0814_
rlabel metal1 4554 44506 4554 44506 0 _0815_
rlabel metal2 43102 6562 43102 6562 0 _0816_
rlabel metal2 47150 41378 47150 41378 0 _0817_
rlabel metal2 48162 37468 48162 37468 0 _0818_
rlabel metal2 16698 45662 16698 45662 0 _0819_
rlabel metal2 47886 44642 47886 44642 0 _0820_
rlabel metal2 25990 3740 25990 3740 0 _0821_
rlabel metal2 38962 3502 38962 3502 0 _0822_
rlabel metal1 42228 45526 42228 45526 0 _0823_
rlabel metal1 25208 2618 25208 2618 0 _0824_
rlabel metal2 47058 5678 47058 5678 0 _0825_
rlabel metal1 4278 31994 4278 31994 0 _0826_
rlabel metal2 47886 17442 47886 17442 0 _0827_
rlabel metal2 12926 46308 12926 46308 0 _0828_
rlabel metal1 4462 2346 4462 2346 0 _0829_
rlabel metal2 10718 3740 10718 3740 0 _0830_
rlabel metal1 2852 16558 2852 16558 0 _0831_
rlabel metal1 46920 28594 46920 28594 0 _0832_
rlabel metal2 48162 14620 48162 14620 0 _0833_
rlabel metal2 47886 13090 47886 13090 0 _0834_
rlabel metal2 3082 4964 3082 4964 0 _0835_
rlabel metal1 13754 46138 13754 46138 0 _0836_
rlabel metal1 44390 4182 44390 4182 0 _0837_
rlabel metal2 13386 3502 13386 3502 0 _0838_
rlabel metal1 35604 45866 35604 45866 0 _0839_
rlabel metal1 14536 46138 14536 46138 0 _0840_
rlabel metal2 46690 21148 46690 21148 0 _0841_
rlabel metal1 6072 46138 6072 46138 0 _0842_
rlabel metal2 4370 3230 4370 3230 0 _0843_
rlabel metal1 24380 45866 24380 45866 0 _0844_
rlabel metal1 25116 45594 25116 45594 0 _0845_
rlabel metal1 47012 2346 47012 2346 0 _0846_
rlabel metal2 47886 39202 47886 39202 0 _0847_
rlabel metal1 29256 46138 29256 46138 0 _0848_
rlabel metal2 42826 3230 42826 3230 0 _0849_
rlabel metal1 46874 32946 46874 32946 0 _0850_
rlabel metal2 3542 46750 3542 46750 0 _0851_
rlabel metal2 40802 3740 40802 3740 0 _0852_
rlabel metal1 2898 24718 2898 24718 0 _0853_
rlabel metal1 45034 2346 45034 2346 0 _0854_
rlabel metal1 10672 45594 10672 45594 0 _0855_
rlabel metal1 2898 22406 2898 22406 0 _0856_
rlabel metal2 2254 11934 2254 11934 0 _0857_
rlabel metal1 2300 17850 2300 17850 0 _0858_
rlabel metal2 4094 46359 4094 46359 0 active
rlabel metal1 18032 30294 18032 30294 0 clknet_0_wb_clk_i
rlabel metal1 17342 19754 17342 19754 0 clknet_4_0_0_wb_clk_i
rlabel metal1 39652 12818 39652 12818 0 clknet_4_10_0_wb_clk_i
rlabel metal2 37766 18496 37766 18496 0 clknet_4_11_0_wb_clk_i
rlabel metal2 34270 23936 34270 23936 0 clknet_4_12_0_wb_clk_i
rlabel metal2 35374 33490 35374 33490 0 clknet_4_13_0_wb_clk_i
rlabel metal1 39238 24174 39238 24174 0 clknet_4_14_0_wb_clk_i
rlabel metal2 38042 33456 38042 33456 0 clknet_4_15_0_wb_clk_i
rlabel metal1 13570 23630 13570 23630 0 clknet_4_1_0_wb_clk_i
rlabel metal1 19734 13838 19734 13838 0 clknet_4_2_0_wb_clk_i
rlabel metal1 20378 22508 20378 22508 0 clknet_4_3_0_wb_clk_i
rlabel metal2 18446 29886 18446 29886 0 clknet_4_4_0_wb_clk_i
rlabel metal1 16560 38318 16560 38318 0 clknet_4_5_0_wb_clk_i
rlabel metal1 21666 29614 21666 29614 0 clknet_4_6_0_wb_clk_i
rlabel metal2 24610 37774 24610 37774 0 clknet_4_7_0_wb_clk_i
rlabel metal1 26105 10642 26105 10642 0 clknet_4_8_0_wb_clk_i
rlabel metal1 32798 21930 32798 21930 0 clknet_4_9_0_wb_clk_i
rlabel metal1 8234 35054 8234 35054 0 gps_channel0.ca_gen.g1\[10\]
rlabel metal1 7728 33082 7728 33082 0 gps_channel0.ca_gen.g1\[1\]
rlabel metal1 9062 33286 9062 33286 0 gps_channel0.ca_gen.g1\[2\]
rlabel metal2 10350 33660 10350 33660 0 gps_channel0.ca_gen.g1\[3\]
rlabel metal2 5290 33558 5290 33558 0 gps_channel0.ca_gen.g1\[4\]
rlabel metal2 5474 35360 5474 35360 0 gps_channel0.ca_gen.g1\[5\]
rlabel metal2 5474 36448 5474 36448 0 gps_channel0.ca_gen.g1\[6\]
rlabel metal1 6578 37434 6578 37434 0 gps_channel0.ca_gen.g1\[7\]
rlabel metal2 7958 37536 7958 37536 0 gps_channel0.ca_gen.g1\[8\]
rlabel metal2 9246 36448 9246 36448 0 gps_channel0.ca_gen.g1\[9\]
rlabel metal2 7222 27812 7222 27812 0 gps_channel0.ca_gen.g2\[10\]
rlabel metal1 13662 30906 13662 30906 0 gps_channel0.ca_gen.g2\[1\]
rlabel metal2 12190 29920 12190 29920 0 gps_channel0.ca_gen.g2\[2\]
rlabel metal1 10718 30090 10718 30090 0 gps_channel0.ca_gen.g2\[3\]
rlabel metal2 10350 32640 10350 32640 0 gps_channel0.ca_gen.g2\[4\]
rlabel metal1 9568 28594 9568 28594 0 gps_channel0.ca_gen.g2\[5\]
rlabel metal2 10258 25503 10258 25503 0 gps_channel0.ca_gen.g2\[6\]
rlabel metal2 10166 23936 10166 23936 0 gps_channel0.ca_gen.g2\[7\]
rlabel metal1 9568 24922 9568 24922 0 gps_channel0.ca_gen.g2\[8\]
rlabel metal1 7590 26962 7590 26962 0 gps_channel0.ca_gen.g2\[9\]
rlabel metal2 11822 27472 11822 27472 0 gps_channel0.ca_gen.g2_init\[10\]
rlabel metal2 17250 29002 17250 29002 0 gps_channel0.ca_gen.g2_init\[1\]
rlabel metal1 16606 31688 16606 31688 0 gps_channel0.ca_gen.g2_init\[2\]
rlabel metal2 17894 29852 17894 29852 0 gps_channel0.ca_gen.g2_init\[3\]
rlabel metal1 12650 31722 12650 31722 0 gps_channel0.ca_gen.g2_init\[4\]
rlabel metal2 11730 33082 11730 33082 0 gps_channel0.ca_gen.g2_init\[5\]
rlabel metal1 13064 29002 13064 29002 0 gps_channel0.ca_gen.g2_init\[6\]
rlabel via1 12374 24582 12374 24582 0 gps_channel0.ca_gen.g2_init\[7\]
rlabel metal2 11730 23222 11730 23222 0 gps_channel0.ca_gen.g2_init\[8\]
rlabel metal1 11086 25262 11086 25262 0 gps_channel0.ca_gen.g2_init\[9\]
rlabel metal1 24610 30022 24610 30022 0 gps_channel0.ca_nco.accumulator\[0\]
rlabel metal1 24748 18734 24748 18734 0 gps_channel0.ca_nco.accumulator\[10\]
rlabel metal1 25530 15470 25530 15470 0 gps_channel0.ca_nco.accumulator\[11\]
rlabel metal1 19780 16422 19780 16422 0 gps_channel0.ca_nco.accumulator\[12\]
rlabel metal2 17342 11696 17342 11696 0 gps_channel0.ca_nco.accumulator\[13\]
rlabel metal1 20562 10030 20562 10030 0 gps_channel0.ca_nco.accumulator\[14\]
rlabel metal1 24840 10778 24840 10778 0 gps_channel0.ca_nco.accumulator\[15\]
rlabel metal1 23000 31858 23000 31858 0 gps_channel0.ca_nco.accumulator\[16\]
rlabel metal1 19458 31314 19458 31314 0 gps_channel0.ca_nco.accumulator\[17\]
rlabel metal2 17802 33694 17802 33694 0 gps_channel0.ca_nco.accumulator\[18\]
rlabel metal1 18216 34510 18216 34510 0 gps_channel0.ca_nco.accumulator\[19\]
rlabel metal2 27370 30498 27370 30498 0 gps_channel0.ca_nco.accumulator\[1\]
rlabel metal2 25898 34833 25898 34833 0 gps_channel0.ca_nco.accumulator\[20\]
rlabel metal2 25162 35360 25162 35360 0 gps_channel0.ca_nco.accumulator\[21\]
rlabel metal1 24794 36040 24794 36040 0 gps_channel0.ca_nco.accumulator\[22\]
rlabel metal2 23230 35428 23230 35428 0 gps_channel0.ca_nco.accumulator\[23\]
rlabel metal2 20654 38148 20654 38148 0 gps_channel0.ca_nco.accumulator\[24\]
rlabel metal2 18906 38726 18906 38726 0 gps_channel0.ca_nco.accumulator\[25\]
rlabel metal2 25622 38964 25622 38964 0 gps_channel0.ca_nco.accumulator\[26\]
rlabel metal1 24242 38862 24242 38862 0 gps_channel0.ca_nco.accumulator\[27\]
rlabel metal2 14766 39712 14766 39712 0 gps_channel0.ca_nco.accumulator\[28\]
rlabel metal2 14950 39440 14950 39440 0 gps_channel0.ca_nco.accumulator\[29\]
rlabel metal2 23230 23222 23230 23222 0 gps_channel0.ca_nco.accumulator\[2\]
rlabel metal2 16974 39236 16974 39236 0 gps_channel0.ca_nco.accumulator\[30\]
rlabel metal2 7130 29648 7130 29648 0 gps_channel0.ca_nco.accumulator\[31\]
rlabel metal2 21482 26112 21482 26112 0 gps_channel0.ca_nco.accumulator\[3\]
rlabel metal1 18446 28186 18446 28186 0 gps_channel0.ca_nco.accumulator\[4\]
rlabel metal1 16721 24786 16721 24786 0 gps_channel0.ca_nco.accumulator\[5\]
rlabel metal1 17526 21896 17526 21896 0 gps_channel0.ca_nco.accumulator\[6\]
rlabel metal1 15502 20026 15502 20026 0 gps_channel0.ca_nco.accumulator\[7\]
rlabel metal2 17158 18054 17158 18054 0 gps_channel0.ca_nco.accumulator\[8\]
rlabel metal2 14398 15232 14398 15232 0 gps_channel0.ca_nco.accumulator\[9\]
rlabel metal2 23414 28288 23414 28288 0 gps_channel0.ca_nco.phase_in\[0\]
rlabel metal1 26450 18632 26450 18632 0 gps_channel0.ca_nco.phase_in\[10\]
rlabel metal2 27830 16252 27830 16252 0 gps_channel0.ca_nco.phase_in\[11\]
rlabel metal1 21620 17170 21620 17170 0 gps_channel0.ca_nco.phase_in\[12\]
rlabel metal2 21666 13124 21666 13124 0 gps_channel0.ca_nco.phase_in\[13\]
rlabel metal1 23736 12206 23736 12206 0 gps_channel0.ca_nco.phase_in\[14\]
rlabel metal1 25668 12954 25668 12954 0 gps_channel0.ca_nco.phase_in\[15\]
rlabel metal1 23138 29478 23138 29478 0 gps_channel0.ca_nco.phase_in\[1\]
rlabel metal1 22356 21658 22356 21658 0 gps_channel0.ca_nco.phase_in\[2\]
rlabel metal1 21114 28526 21114 28526 0 gps_channel0.ca_nco.phase_in\[3\]
rlabel metal1 18308 28934 18308 28934 0 gps_channel0.ca_nco.phase_in\[4\]
rlabel metal1 20286 24140 20286 24140 0 gps_channel0.ca_nco.phase_in\[5\]
rlabel metal1 19458 22032 19458 22032 0 gps_channel0.ca_nco.phase_in\[6\]
rlabel metal2 20378 20026 20378 20026 0 gps_channel0.ca_nco.phase_in\[7\]
rlabel metal2 21482 18462 21482 18462 0 gps_channel0.ca_nco.phase_in\[8\]
rlabel metal1 20608 18258 20608 18258 0 gps_channel0.ca_nco.phase_in\[9\]
rlabel metal2 26266 24956 26266 24956 0 gps_channel0.ca_nco.phase_sync
rlabel metal1 24840 28526 24840 28526 0 gps_channel0.ca_nco.step\[0\]
rlabel metal2 25254 19652 25254 19652 0 gps_channel0.ca_nco.step\[10\]
rlabel metal2 25530 14110 25530 14110 0 gps_channel0.ca_nco.step\[11\]
rlabel metal2 18814 14586 18814 14586 0 gps_channel0.ca_nco.step\[12\]
rlabel metal1 18722 13260 18722 13260 0 gps_channel0.ca_nco.step\[13\]
rlabel metal2 18906 10234 18906 10234 0 gps_channel0.ca_nco.step\[14\]
rlabel metal2 23230 9758 23230 9758 0 gps_channel0.ca_nco.step\[15\]
rlabel metal1 23690 36142 23690 36142 0 gps_channel0.ca_nco.step\[16\]
rlabel metal2 27554 29648 27554 29648 0 gps_channel0.ca_nco.step\[1\]
rlabel metal1 25392 21998 25392 21998 0 gps_channel0.ca_nco.step\[2\]
rlabel metal2 21666 25534 21666 25534 0 gps_channel0.ca_nco.step\[3\]
rlabel metal1 16905 26418 16905 26418 0 gps_channel0.ca_nco.step\[4\]
rlabel metal1 16882 24242 16882 24242 0 gps_channel0.ca_nco.step\[5\]
rlabel metal1 16652 22610 16652 22610 0 gps_channel0.ca_nco.step\[6\]
rlabel metal2 13478 19516 13478 19516 0 gps_channel0.ca_nco.step\[7\]
rlabel metal1 13708 17850 13708 17850 0 gps_channel0.ca_nco.step\[8\]
rlabel metal2 13294 17408 13294 17408 0 gps_channel0.ca_nco.step\[9\]
rlabel metal1 21850 24276 21850 24276 0 gps_channel0.lo_i
rlabel metal1 31786 31790 31786 31790 0 gps_channel0.lo_nco.accumulator\[0\]
rlabel metal1 34086 19346 34086 19346 0 gps_channel0.lo_nco.accumulator\[10\]
rlabel metal1 35098 17612 35098 17612 0 gps_channel0.lo_nco.accumulator\[11\]
rlabel metal1 35512 15878 35512 15878 0 gps_channel0.lo_nco.accumulator\[12\]
rlabel metal2 33994 14620 33994 14620 0 gps_channel0.lo_nco.accumulator\[13\]
rlabel metal1 37582 12614 37582 12614 0 gps_channel0.lo_nco.accumulator\[14\]
rlabel metal2 34730 11934 34730 11934 0 gps_channel0.lo_nco.accumulator\[15\]
rlabel metal2 44390 14858 44390 14858 0 gps_channel0.lo_nco.accumulator\[16\]
rlabel metal2 44482 17442 44482 17442 0 gps_channel0.lo_nco.accumulator\[17\]
rlabel metal2 44574 18258 44574 18258 0 gps_channel0.lo_nco.accumulator\[18\]
rlabel metal1 44436 20366 44436 20366 0 gps_channel0.lo_nco.accumulator\[19\]
rlabel metal1 31556 32334 31556 32334 0 gps_channel0.lo_nco.accumulator\[1\]
rlabel metal2 39974 16218 39974 16218 0 gps_channel0.lo_nco.accumulator\[20\]
rlabel metal2 40986 15402 40986 15402 0 gps_channel0.lo_nco.accumulator\[21\]
rlabel metal2 40250 19380 40250 19380 0 gps_channel0.lo_nco.accumulator\[22\]
rlabel metal1 40756 19822 40756 19822 0 gps_channel0.lo_nco.accumulator\[23\]
rlabel metal1 41860 22610 41860 22610 0 gps_channel0.lo_nco.accumulator\[24\]
rlabel metal1 42412 24378 42412 24378 0 gps_channel0.lo_nco.accumulator\[25\]
rlabel metal2 45586 25058 45586 25058 0 gps_channel0.lo_nco.accumulator\[26\]
rlabel metal1 44896 25806 44896 25806 0 gps_channel0.lo_nco.accumulator\[27\]
rlabel metal1 46230 30906 46230 30906 0 gps_channel0.lo_nco.accumulator\[28\]
rlabel metal1 44850 31450 44850 31450 0 gps_channel0.lo_nco.accumulator\[29\]
rlabel metal2 36846 34782 36846 34782 0 gps_channel0.lo_nco.accumulator\[2\]
rlabel metal1 18446 30260 18446 30260 0 gps_channel0.lo_nco.accumulator\[30\]
rlabel metal1 33626 33830 33626 33830 0 gps_channel0.lo_nco.accumulator\[3\]
rlabel metal1 39376 31790 39376 31790 0 gps_channel0.lo_nco.accumulator\[4\]
rlabel metal1 39882 29648 39882 29648 0 gps_channel0.lo_nco.accumulator\[5\]
rlabel metal1 38548 25874 38548 25874 0 gps_channel0.lo_nco.accumulator\[6\]
rlabel metal2 36386 27234 36386 27234 0 gps_channel0.lo_nco.accumulator\[7\]
rlabel metal1 36662 23630 36662 23630 0 gps_channel0.lo_nco.accumulator\[8\]
rlabel metal1 33994 21556 33994 21556 0 gps_channel0.lo_nco.accumulator\[9\]
rlabel metal1 29808 29614 29808 29614 0 gps_channel0.lo_nco.phase_in\[0\]
rlabel metal1 32177 19414 32177 19414 0 gps_channel0.lo_nco.phase_in\[10\]
rlabel metal1 36202 17578 36202 17578 0 gps_channel0.lo_nco.phase_in\[11\]
rlabel metal1 33810 15504 33810 15504 0 gps_channel0.lo_nco.phase_in\[12\]
rlabel metal1 32062 15436 32062 15436 0 gps_channel0.lo_nco.phase_in\[13\]
rlabel metal2 29118 12274 29118 12274 0 gps_channel0.lo_nco.phase_in\[14\]
rlabel metal1 31142 12206 31142 12206 0 gps_channel0.lo_nco.phase_in\[15\]
rlabel metal2 33442 28322 33442 28322 0 gps_channel0.lo_nco.phase_in\[1\]
rlabel metal1 34960 31450 34960 31450 0 gps_channel0.lo_nco.phase_in\[2\]
rlabel metal1 33442 32470 33442 32470 0 gps_channel0.lo_nco.phase_in\[3\]
rlabel metal1 36846 29104 36846 29104 0 gps_channel0.lo_nco.phase_in\[4\]
rlabel metal2 36478 29478 36478 29478 0 gps_channel0.lo_nco.phase_in\[5\]
rlabel metal2 38410 25602 38410 25602 0 gps_channel0.lo_nco.phase_in\[6\]
rlabel metal2 33442 26792 33442 26792 0 gps_channel0.lo_nco.phase_in\[7\]
rlabel metal1 34592 24038 34592 24038 0 gps_channel0.lo_nco.phase_in\[8\]
rlabel metal1 31280 21386 31280 21386 0 gps_channel0.lo_nco.phase_in\[9\]
rlabel metal1 31234 24174 31234 24174 0 gps_channel0.lo_nco.phase_sync
rlabel metal2 31234 34714 31234 34714 0 gps_channel0.lo_nco.step\[0\]
rlabel metal1 34086 19482 34086 19482 0 gps_channel0.lo_nco.step\[10\]
rlabel metal2 33810 17952 33810 17952 0 gps_channel0.lo_nco.step\[11\]
rlabel metal1 32752 15878 32752 15878 0 gps_channel0.lo_nco.step\[12\]
rlabel metal1 33350 13906 33350 13906 0 gps_channel0.lo_nco.step\[13\]
rlabel metal2 31142 10812 31142 10812 0 gps_channel0.lo_nco.step\[14\]
rlabel metal2 33074 11492 33074 11492 0 gps_channel0.lo_nco.step\[15\]
rlabel metal1 40388 21998 40388 21998 0 gps_channel0.lo_nco.step\[16\]
rlabel metal1 30774 33082 30774 33082 0 gps_channel0.lo_nco.step\[1\]
rlabel metal2 37674 34748 37674 34748 0 gps_channel0.lo_nco.step\[2\]
rlabel metal2 33534 35292 33534 35292 0 gps_channel0.lo_nco.step\[3\]
rlabel metal1 39468 34034 39468 34034 0 gps_channel0.lo_nco.step\[4\]
rlabel metal1 41400 31994 41400 31994 0 gps_channel0.lo_nco.step\[5\]
rlabel metal1 38456 24718 38456 24718 0 gps_channel0.lo_nco.step\[6\]
rlabel metal2 36570 27200 36570 27200 0 gps_channel0.lo_nco.step\[7\]
rlabel metal1 35512 23154 35512 23154 0 gps_channel0.lo_nco.step\[8\]
rlabel metal1 33074 22202 33074 22202 0 gps_channel0.lo_nco.step\[9\]
rlabel metal2 6578 31484 6578 31484 0 gps_channel0.prompt_i
rlabel metal2 6762 29852 6762 29852 0 gps_channel0.prompt_q
rlabel metal1 9200 47022 9200 47022 0 io_in[23]
rlabel metal2 26450 2166 26450 2166 0 io_oeb[0]
rlabel via2 2898 17085 2898 17085 0 io_oeb[10]
rlabel metal3 48814 28628 48814 28628 0 io_oeb[11]
rlabel metal2 46874 14739 46874 14739 0 io_oeb[12]
rlabel metal2 46874 13515 46874 13515 0 io_oeb[13]
rlabel metal3 1740 4828 1740 4828 0 io_oeb[14]
rlabel metal1 14490 47090 14490 47090 0 io_oeb[15]
rlabel via2 46874 2091 46874 2091 0 io_oeb[16]
rlabel metal1 13616 2958 13616 2958 0 io_oeb[17]
rlabel metal2 36110 47644 36110 47644 0 io_oeb[18]
rlabel metal2 14858 47882 14858 47882 0 io_oeb[19]
rlabel metal2 39330 1860 39330 1860 0 io_oeb[1]
rlabel metal3 48814 21828 48814 21828 0 io_oeb[20]
rlabel metal2 1978 47984 1978 47984 0 io_oeb[21]
rlabel metal2 5198 1860 5198 1860 0 io_oeb[22]
rlabel metal2 25162 47644 25162 47644 0 io_oeb[23]
rlabel metal2 25806 47882 25806 47882 0 io_oeb[24]
rlabel metal1 47242 2482 47242 2482 0 io_oeb[25]
rlabel via2 46874 39491 46874 39491 0 io_oeb[26]
rlabel metal2 29670 47882 29670 47882 0 io_oeb[27]
rlabel metal1 42504 2822 42504 2822 0 io_oeb[28]
rlabel metal3 48860 32708 48860 32708 0 io_oeb[29]
rlabel metal1 43102 46444 43102 46444 0 io_oeb[2]
rlabel metal2 2622 47882 2622 47882 0 io_oeb[30]
rlabel metal2 41262 2166 41262 2166 0 io_oeb[31]
rlabel metal3 1142 25228 1142 25228 0 io_oeb[32]
rlabel metal1 44114 2516 44114 2516 0 io_oeb[33]
rlabel metal1 11040 46002 11040 46002 0 io_oeb[34]
rlabel metal3 1142 21828 1142 21828 0 io_oeb[35]
rlabel metal3 1740 11628 1740 11628 0 io_oeb[36]
rlabel metal2 2806 18309 2806 18309 0 io_oeb[37]
rlabel metal2 25806 1860 25806 1860 0 io_oeb[3]
rlabel metal3 48906 68 48906 68 0 io_oeb[4]
rlabel metal1 4186 32334 4186 32334 0 io_oeb[5]
rlabel via2 46874 17731 46874 17731 0 io_oeb[6]
rlabel metal2 13018 46529 13018 46529 0 io_oeb[7]
rlabel metal2 4554 1622 4554 1622 0 io_oeb[8]
rlabel metal2 10994 2166 10994 2166 0 io_oeb[9]
rlabel metal1 43562 45390 43562 45390 0 io_out[0]
rlabel metal2 46874 27727 46874 27727 0 io_out[10]
rlabel metal3 1142 2788 1142 2788 0 io_out[11]
rlabel metal3 1142 7548 1142 7548 0 io_out[12]
rlabel metal2 40618 1503 40618 1503 0 io_out[13]
rlabel metal3 48860 40188 48860 40188 0 io_out[14]
rlabel via2 3082 41531 3082 41531 0 io_out[15]
rlabel metal2 46874 25959 46874 25959 0 io_out[16]
rlabel metal2 46414 47882 46414 47882 0 io_out[17]
rlabel metal2 47058 1761 47058 1761 0 io_out[18]
rlabel metal3 2016 23868 2016 23868 0 io_out[19]
rlabel metal2 33534 47882 33534 47882 0 io_out[1]
rlabel metal2 40618 47644 40618 47644 0 io_out[20]
rlabel metal3 1970 40868 1970 40868 0 io_out[21]
rlabel metal1 32292 6834 32292 6834 0 io_out[22]
rlabel metal3 48124 22508 48124 22508 0 io_out[23]
rlabel metal2 27738 1860 27738 1860 0 io_out[24]
rlabel metal1 37950 46444 37950 46444 0 io_out[25]
rlabel metal3 1142 5508 1142 5508 0 io_out[26]
rlabel metal1 40250 46444 40250 46444 0 io_out[27]
rlabel metal2 17434 1860 17434 1860 0 io_out[28]
rlabel metal3 48078 1428 48078 1428 0 io_out[29]
rlabel metal2 7130 1622 7130 1622 0 io_out[2]
rlabel metal3 1142 6868 1142 6868 0 io_out[30]
rlabel metal3 1142 14348 1142 14348 0 io_out[31]
rlabel metal2 2806 46835 2806 46835 0 io_out[32]
rlabel metal3 48124 6868 48124 6868 0 io_out[33]
rlabel metal3 48814 41548 48814 41548 0 io_out[34]
rlabel metal2 46506 37689 46506 37689 0 io_out[35]
rlabel metal2 15502 47644 15502 47644 0 io_out[36]
rlabel via2 46874 44931 46874 44931 0 io_out[37]
rlabel metal2 2806 43401 2806 43401 0 io_out[3]
rlabel metal3 48860 29308 48860 29308 0 io_out[4]
rlabel metal2 23230 47882 23230 47882 0 io_out[5]
rlabel metal2 48346 47644 48346 47644 0 io_out[6]
rlabel metal2 2806 20417 2806 20417 0 io_out[7]
rlabel metal2 19366 1571 19366 1571 0 io_out[8]
rlabel via2 3450 15045 3450 15045 0 io_out[9]
rlabel metal1 48300 8466 48300 8466 0 la1_data_in[0]
rlabel metal1 32062 47022 32062 47022 0 la1_data_in[16]
rlabel metal1 24242 47022 24242 47022 0 la1_data_in[17]
rlabel metal1 43930 3434 43930 3434 0 la1_data_in[18]
rlabel metal2 17526 47617 17526 47617 0 la1_data_in[19]
rlabel metal1 20056 3502 20056 3502 0 la1_data_in[1]
rlabel metal3 1188 36788 1188 36788 0 la1_data_in[20]
rlabel metal1 48622 47022 48622 47022 0 la1_data_in[21]
rlabel via2 48254 8891 48254 8891 0 la1_data_in[22]
rlabel metal3 1740 748 1740 748 0 la1_data_in[23]
rlabel metal2 14214 1588 14214 1588 0 la1_data_in[24]
rlabel metal3 1188 38828 1188 38828 0 la1_data_in[25]
rlabel via2 48346 3485 48346 3485 0 la1_data_in[26]
rlabel metal2 29026 1554 29026 1554 0 la1_data_in[27]
rlabel metal3 1142 34068 1142 34068 0 la1_data_in[28]
rlabel metal2 1334 48086 1334 48086 0 la1_data_in[29]
rlabel metal2 11638 1894 11638 1894 0 la1_data_in[2]
rlabel metal2 1334 2676 1334 2676 0 la1_data_in[30]
rlabel metal2 38686 1554 38686 1554 0 la1_data_in[31]
rlabel metal3 1142 32028 1142 32028 0 la1_data_in[3]
rlabel metal1 42596 47022 42596 47022 0 la1_data_in[4]
rlabel metal2 48254 24667 48254 24667 0 la1_data_in[5]
rlabel metal1 19412 47022 19412 47022 0 la1_data_in[6]
rlabel metal2 7774 1860 7774 1860 0 la1_data_out[0]
rlabel metal3 48676 12308 48676 12308 0 la1_data_out[10]
rlabel metal2 22586 823 22586 823 0 la1_data_out[11]
rlabel metal3 47480 46308 47480 46308 0 la1_data_out[12]
rlabel metal1 13018 46376 13018 46376 0 la1_data_out[13]
rlabel metal2 27094 47814 27094 47814 0 la1_data_out[14]
rlabel metal3 1786 1428 1786 1428 0 la1_data_out[15]
rlabel metal3 48768 17068 48768 17068 0 la1_data_out[16]
rlabel metal2 46874 36159 46874 36159 0 la1_data_out[17]
rlabel metal2 5842 47933 5842 47933 0 la1_data_out[18]
rlabel metal2 46782 25857 46782 25857 0 la1_data_out[19]
rlabel metal2 3174 44965 3174 44965 0 la1_data_out[1]
rlabel metal3 1142 10268 1142 10268 0 la1_data_out[20]
rlabel metal3 48814 42908 48814 42908 0 la1_data_out[21]
rlabel metal1 30360 46002 30360 46002 0 la1_data_out[22]
rlabel metal2 12926 1622 12926 1622 0 la1_data_out[23]
rlabel metal3 48814 19108 48814 19108 0 la1_data_out[24]
rlabel metal3 1142 3468 1142 3468 0 la1_data_out[25]
rlabel metal2 46874 5083 46874 5083 0 la1_data_out[26]
rlabel metal2 2898 46869 2898 46869 0 la1_data_out[27]
rlabel metal2 45126 1367 45126 1367 0 la1_data_out[28]
rlabel metal2 6486 2166 6486 2166 0 la1_data_out[29]
rlabel metal2 20654 1860 20654 1860 0 la1_data_out[2]
rlabel metal3 48814 12988 48814 12988 0 la1_data_out[30]
rlabel metal2 46782 48059 46782 48059 0 la1_data_out[31]
rlabel metal3 1832 9588 1832 9588 0 la1_data_out[3]
rlabel metal2 45770 2404 45770 2404 0 la1_data_out[4]
rlabel metal2 3266 1860 3266 1860 0 la1_data_out[5]
rlabel metal3 48814 20468 48814 20468 0 la1_data_out[6]
rlabel metal2 460 16560 460 16560 0 la1_data_out[7]
rlabel metal3 48676 37468 48676 37468 0 la1_data_out[8]
rlabel metal1 47288 32470 47288 32470 0 la1_data_out[9]
rlabel metal1 2714 47124 2714 47124 0 net1
rlabel metal2 20010 23936 20010 23936 0 net10
rlabel metal1 14030 47022 14030 47022 0 net100
rlabel metal1 44482 3978 44482 3978 0 net101
rlabel metal2 13202 3264 13202 3264 0 net102
rlabel metal2 35374 46172 35374 46172 0 net103
rlabel metal1 14444 45458 14444 45458 0 net104
rlabel metal1 46506 21012 46506 21012 0 net105
rlabel metal2 6026 46818 6026 46818 0 net106
rlabel metal1 4600 2958 4600 2958 0 net107
rlabel metal1 24656 45458 24656 45458 0 net108
rlabel metal1 24794 46580 24794 46580 0 net109
rlabel metal2 21298 22950 21298 22950 0 net11
rlabel metal1 47518 2414 47518 2414 0 net110
rlabel metal2 48346 39644 48346 39644 0 net111
rlabel metal1 28980 46478 28980 46478 0 net112
rlabel metal1 42274 2958 42274 2958 0 net113
rlabel metal1 47472 32402 47472 32402 0 net114
rlabel metal1 4140 46546 4140 46546 0 net115
rlabel metal1 40848 3026 40848 3026 0 net116
rlabel metal2 3450 25500 3450 25500 0 net117
rlabel metal1 44712 2482 44712 2482 0 net118
rlabel metal2 10534 46172 10534 46172 0 net119
rlabel metal2 7222 3842 7222 3842 0 net12
rlabel metal2 3450 21760 3450 21760 0 net120
rlabel metal2 2070 11492 2070 11492 0 net121
rlabel metal2 2070 18496 2070 18496 0 net122
rlabel metal1 13570 2618 13570 2618 0 net13
rlabel metal2 1886 33048 1886 33048 0 net14
rlabel metal2 30314 5269 30314 5269 0 net15
rlabel metal1 29808 2618 29808 2618 0 net16
rlabel metal1 1886 34714 1886 34714 0 net17
rlabel metal2 21390 13634 21390 13634 0 net18
rlabel metal2 17986 31484 17986 31484 0 net19
rlabel metal1 8326 35156 8326 35156 0 net2
rlabel metal1 4347 4726 4347 4726 0 net20
rlabel metal1 34776 2278 34776 2278 0 net21
rlabel metal2 5474 32674 5474 32674 0 net22
rlabel metal1 43240 47158 43240 47158 0 net23
rlabel metal2 32246 22712 32246 22712 0 net24
rlabel metal1 20056 47158 20056 47158 0 net25
rlabel metal2 7498 3264 7498 3264 0 net26
rlabel metal2 2070 44608 2070 44608 0 net27
rlabel metal1 19872 2958 19872 2958 0 net28
rlabel metal1 2116 9146 2116 9146 0 net29
rlabel metal1 25668 12206 25668 12206 0 net3
rlabel metal2 46782 4352 46782 4352 0 net30
rlabel metal2 3726 3468 3726 3468 0 net31
rlabel metal2 46506 20060 46506 20060 0 net32
rlabel metal1 46782 23698 46782 23698 0 net33
rlabel metal2 48346 36380 48346 36380 0 net34
rlabel metal2 7314 43996 7314 43996 0 net35
rlabel metal2 47242 25296 47242 25296 0 net36
rlabel metal1 3450 10132 3450 10132 0 net37
rlabel metal1 46782 42738 46782 42738 0 net38
rlabel metal2 29762 46512 29762 46512 0 net39
rlabel metal1 17342 28628 17342 28628 0 net4
rlabel metal1 12190 2482 12190 2482 0 net40
rlabel metal1 46506 18836 46506 18836 0 net41
rlabel metal1 4094 3570 4094 3570 0 net42
rlabel metal2 48346 4828 48346 4828 0 net43
rlabel metal1 4462 45390 4462 45390 0 net44
rlabel metal1 44896 3570 44896 3570 0 net45
rlabel metal1 5704 3502 5704 3502 0 net46
rlabel metal1 46782 12342 46782 12342 0 net47
rlabel metal2 47242 45696 47242 45696 0 net48
rlabel metal2 38962 46240 38962 46240 0 net49
rlabel metal1 25070 33354 25070 33354 0 net5
rlabel metal1 33074 46580 33074 46580 0 net50
rlabel metal2 6670 2652 6670 2652 0 net51
rlabel metal2 2070 43520 2070 43520 0 net52
rlabel metal2 46506 29852 46506 29852 0 net53
rlabel metal2 22494 46784 22494 46784 0 net54
rlabel metal1 45954 46002 45954 46002 0 net55
rlabel metal2 2070 20672 2070 20672 0 net56
rlabel metal1 19412 2482 19412 2482 0 net57
rlabel metal2 6026 15232 6026 15232 0 net58
rlabel metal2 48346 28254 48346 28254 0 net59
rlabel metal1 21390 29512 21390 29512 0 net6
rlabel metal1 3220 2482 3220 2482 0 net60
rlabel metal1 2346 7412 2346 7412 0 net61
rlabel metal2 39054 4352 39054 4352 0 net62
rlabel metal2 46506 40732 46506 40732 0 net63
rlabel metal2 7314 41820 7314 41820 0 net64
rlabel metal2 48346 25500 48346 25500 0 net65
rlabel metal1 45402 46444 45402 46444 0 net66
rlabel metal2 46138 6256 46138 6256 0 net67
rlabel metal2 40158 46512 40158 46512 0 net68
rlabel metal1 31648 6766 31648 6766 0 net69
rlabel metal1 20470 27982 20470 27982 0 net7
rlabel metal1 48162 22406 48162 22406 0 net70
rlabel metal2 27186 3264 27186 3264 0 net71
rlabel metal1 36892 46478 36892 46478 0 net72
rlabel metal2 3450 5916 3450 5916 0 net73
rlabel metal2 39790 46818 39790 46818 0 net74
rlabel metal2 16882 3264 16882 3264 0 net75
rlabel metal1 44666 3026 44666 3026 0 net76
rlabel metal2 3450 7004 3450 7004 0 net77
rlabel metal2 3450 14620 3450 14620 0 net78
rlabel metal1 4140 45934 4140 45934 0 net79
rlabel metal1 35282 13430 35282 13430 0 net8
rlabel metal1 43056 6834 43056 6834 0 net80
rlabel metal2 46506 41820 46506 41820 0 net81
rlabel metal2 48346 37774 48346 37774 0 net82
rlabel metal2 16882 46172 16882 46172 0 net83
rlabel metal2 48346 45084 48346 45084 0 net84
rlabel metal1 25576 3502 25576 3502 0 net85
rlabel metal2 38778 3264 38778 3264 0 net86
rlabel metal1 42090 46546 42090 46546 0 net87
rlabel metal2 24794 3468 24794 3468 0 net88
rlabel metal1 47518 4114 47518 4114 0 net89
rlabel metal1 2346 37298 2346 37298 0 net9
rlabel metal2 3818 32640 3818 32640 0 net90
rlabel metal2 48346 17884 48346 17884 0 net91
rlabel metal2 12466 46818 12466 46818 0 net92
rlabel metal2 4094 2703 4094 2703 0 net93
rlabel metal2 10534 3264 10534 3264 0 net94
rlabel metal1 2116 16762 2116 16762 0 net95
rlabel metal2 46506 28764 46506 28764 0 net96
rlabel metal2 48346 14960 48346 14960 0 net97
rlabel metal2 48346 13600 48346 13600 0 net98
rlabel metal2 2530 4930 2530 4930 0 net99
rlabel metal1 30314 24718 30314 24718 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
