// This is the unpowered netlist.
module wrapped_channel (active,
    wb_clk_i,
    io_in,
    io_oeb,
    io_out,
    la1_data_in,
    la1_data_out,
    la1_oenb);
 input active;
 input wb_clk_i;
 input [37:0] io_in;
 inout [37:0] io_oeb;
 inout [37:0] io_out;
 input [31:0] la1_data_in;
 inout [31:0] la1_data_out;
 input [31:0] la1_oenb;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire clknet_0_wb_clk_i;
 wire \gps_channel0.ca_gen.g1[10] ;
 wire \gps_channel0.ca_gen.g1[1] ;
 wire \gps_channel0.ca_gen.g1[2] ;
 wire \gps_channel0.ca_gen.g1[3] ;
 wire \gps_channel0.ca_gen.g1[4] ;
 wire \gps_channel0.ca_gen.g1[5] ;
 wire \gps_channel0.ca_gen.g1[6] ;
 wire \gps_channel0.ca_gen.g1[7] ;
 wire \gps_channel0.ca_gen.g1[8] ;
 wire \gps_channel0.ca_gen.g1[9] ;
 wire \gps_channel0.ca_gen.g2[10] ;
 wire \gps_channel0.ca_gen.g2[1] ;
 wire \gps_channel0.ca_gen.g2[2] ;
 wire \gps_channel0.ca_gen.g2[3] ;
 wire \gps_channel0.ca_gen.g2[4] ;
 wire \gps_channel0.ca_gen.g2[5] ;
 wire \gps_channel0.ca_gen.g2[6] ;
 wire \gps_channel0.ca_gen.g2[7] ;
 wire \gps_channel0.ca_gen.g2[8] ;
 wire \gps_channel0.ca_gen.g2[9] ;
 wire \gps_channel0.ca_gen.g2_init[10] ;
 wire \gps_channel0.ca_gen.g2_init[1] ;
 wire \gps_channel0.ca_gen.g2_init[2] ;
 wire \gps_channel0.ca_gen.g2_init[3] ;
 wire \gps_channel0.ca_gen.g2_init[4] ;
 wire \gps_channel0.ca_gen.g2_init[5] ;
 wire \gps_channel0.ca_gen.g2_init[6] ;
 wire \gps_channel0.ca_gen.g2_init[7] ;
 wire \gps_channel0.ca_gen.g2_init[8] ;
 wire \gps_channel0.ca_gen.g2_init[9] ;
 wire \gps_channel0.ca_nco.accumulator[0] ;
 wire \gps_channel0.ca_nco.accumulator[10] ;
 wire \gps_channel0.ca_nco.accumulator[11] ;
 wire \gps_channel0.ca_nco.accumulator[12] ;
 wire \gps_channel0.ca_nco.accumulator[13] ;
 wire \gps_channel0.ca_nco.accumulator[14] ;
 wire \gps_channel0.ca_nco.accumulator[15] ;
 wire \gps_channel0.ca_nco.accumulator[16] ;
 wire \gps_channel0.ca_nco.accumulator[17] ;
 wire \gps_channel0.ca_nco.accumulator[18] ;
 wire \gps_channel0.ca_nco.accumulator[19] ;
 wire \gps_channel0.ca_nco.accumulator[1] ;
 wire \gps_channel0.ca_nco.accumulator[20] ;
 wire \gps_channel0.ca_nco.accumulator[21] ;
 wire \gps_channel0.ca_nco.accumulator[22] ;
 wire \gps_channel0.ca_nco.accumulator[23] ;
 wire \gps_channel0.ca_nco.accumulator[24] ;
 wire \gps_channel0.ca_nco.accumulator[25] ;
 wire \gps_channel0.ca_nco.accumulator[26] ;
 wire \gps_channel0.ca_nco.accumulator[27] ;
 wire \gps_channel0.ca_nco.accumulator[28] ;
 wire \gps_channel0.ca_nco.accumulator[29] ;
 wire \gps_channel0.ca_nco.accumulator[2] ;
 wire \gps_channel0.ca_nco.accumulator[30] ;
 wire \gps_channel0.ca_nco.accumulator[31] ;
 wire \gps_channel0.ca_nco.accumulator[3] ;
 wire \gps_channel0.ca_nco.accumulator[4] ;
 wire \gps_channel0.ca_nco.accumulator[5] ;
 wire \gps_channel0.ca_nco.accumulator[6] ;
 wire \gps_channel0.ca_nco.accumulator[7] ;
 wire \gps_channel0.ca_nco.accumulator[8] ;
 wire \gps_channel0.ca_nco.accumulator[9] ;
 wire \gps_channel0.ca_nco.phase_in[0] ;
 wire \gps_channel0.ca_nco.phase_in[10] ;
 wire \gps_channel0.ca_nco.phase_in[11] ;
 wire \gps_channel0.ca_nco.phase_in[12] ;
 wire \gps_channel0.ca_nco.phase_in[13] ;
 wire \gps_channel0.ca_nco.phase_in[14] ;
 wire \gps_channel0.ca_nco.phase_in[15] ;
 wire \gps_channel0.ca_nco.phase_in[1] ;
 wire \gps_channel0.ca_nco.phase_in[2] ;
 wire \gps_channel0.ca_nco.phase_in[3] ;
 wire \gps_channel0.ca_nco.phase_in[4] ;
 wire \gps_channel0.ca_nco.phase_in[5] ;
 wire \gps_channel0.ca_nco.phase_in[6] ;
 wire \gps_channel0.ca_nco.phase_in[7] ;
 wire \gps_channel0.ca_nco.phase_in[8] ;
 wire \gps_channel0.ca_nco.phase_in[9] ;
 wire \gps_channel0.ca_nco.phase_sync ;
 wire \gps_channel0.ca_nco.step[0] ;
 wire \gps_channel0.ca_nco.step[10] ;
 wire \gps_channel0.ca_nco.step[11] ;
 wire \gps_channel0.ca_nco.step[12] ;
 wire \gps_channel0.ca_nco.step[13] ;
 wire \gps_channel0.ca_nco.step[14] ;
 wire \gps_channel0.ca_nco.step[15] ;
 wire \gps_channel0.ca_nco.step[16] ;
 wire \gps_channel0.ca_nco.step[1] ;
 wire \gps_channel0.ca_nco.step[2] ;
 wire \gps_channel0.ca_nco.step[3] ;
 wire \gps_channel0.ca_nco.step[4] ;
 wire \gps_channel0.ca_nco.step[5] ;
 wire \gps_channel0.ca_nco.step[6] ;
 wire \gps_channel0.ca_nco.step[7] ;
 wire \gps_channel0.ca_nco.step[8] ;
 wire \gps_channel0.ca_nco.step[9] ;
 wire \gps_channel0.lo_i ;
 wire \gps_channel0.lo_nco.accumulator[0] ;
 wire \gps_channel0.lo_nco.accumulator[10] ;
 wire \gps_channel0.lo_nco.accumulator[11] ;
 wire \gps_channel0.lo_nco.accumulator[12] ;
 wire \gps_channel0.lo_nco.accumulator[13] ;
 wire \gps_channel0.lo_nco.accumulator[14] ;
 wire \gps_channel0.lo_nco.accumulator[15] ;
 wire \gps_channel0.lo_nco.accumulator[16] ;
 wire \gps_channel0.lo_nco.accumulator[17] ;
 wire \gps_channel0.lo_nco.accumulator[18] ;
 wire \gps_channel0.lo_nco.accumulator[19] ;
 wire \gps_channel0.lo_nco.accumulator[1] ;
 wire \gps_channel0.lo_nco.accumulator[20] ;
 wire \gps_channel0.lo_nco.accumulator[21] ;
 wire \gps_channel0.lo_nco.accumulator[22] ;
 wire \gps_channel0.lo_nco.accumulator[23] ;
 wire \gps_channel0.lo_nco.accumulator[24] ;
 wire \gps_channel0.lo_nco.accumulator[25] ;
 wire \gps_channel0.lo_nco.accumulator[26] ;
 wire \gps_channel0.lo_nco.accumulator[27] ;
 wire \gps_channel0.lo_nco.accumulator[28] ;
 wire \gps_channel0.lo_nco.accumulator[29] ;
 wire \gps_channel0.lo_nco.accumulator[2] ;
 wire \gps_channel0.lo_nco.accumulator[30] ;
 wire \gps_channel0.lo_nco.accumulator[3] ;
 wire \gps_channel0.lo_nco.accumulator[4] ;
 wire \gps_channel0.lo_nco.accumulator[5] ;
 wire \gps_channel0.lo_nco.accumulator[6] ;
 wire \gps_channel0.lo_nco.accumulator[7] ;
 wire \gps_channel0.lo_nco.accumulator[8] ;
 wire \gps_channel0.lo_nco.accumulator[9] ;
 wire \gps_channel0.lo_nco.phase_in[0] ;
 wire \gps_channel0.lo_nco.phase_in[10] ;
 wire \gps_channel0.lo_nco.phase_in[11] ;
 wire \gps_channel0.lo_nco.phase_in[12] ;
 wire \gps_channel0.lo_nco.phase_in[13] ;
 wire \gps_channel0.lo_nco.phase_in[14] ;
 wire \gps_channel0.lo_nco.phase_in[15] ;
 wire \gps_channel0.lo_nco.phase_in[1] ;
 wire \gps_channel0.lo_nco.phase_in[2] ;
 wire \gps_channel0.lo_nco.phase_in[3] ;
 wire \gps_channel0.lo_nco.phase_in[4] ;
 wire \gps_channel0.lo_nco.phase_in[5] ;
 wire \gps_channel0.lo_nco.phase_in[6] ;
 wire \gps_channel0.lo_nco.phase_in[7] ;
 wire \gps_channel0.lo_nco.phase_in[8] ;
 wire \gps_channel0.lo_nco.phase_in[9] ;
 wire \gps_channel0.lo_nco.phase_sync ;
 wire \gps_channel0.lo_nco.step[0] ;
 wire \gps_channel0.lo_nco.step[10] ;
 wire \gps_channel0.lo_nco.step[11] ;
 wire \gps_channel0.lo_nco.step[12] ;
 wire \gps_channel0.lo_nco.step[13] ;
 wire \gps_channel0.lo_nco.step[14] ;
 wire \gps_channel0.lo_nco.step[15] ;
 wire \gps_channel0.lo_nco.step[16] ;
 wire \gps_channel0.lo_nco.step[1] ;
 wire \gps_channel0.lo_nco.step[2] ;
 wire \gps_channel0.lo_nco.step[3] ;
 wire \gps_channel0.lo_nco.step[4] ;
 wire \gps_channel0.lo_nco.step[5] ;
 wire \gps_channel0.lo_nco.step[6] ;
 wire \gps_channel0.lo_nco.step[7] ;
 wire \gps_channel0.lo_nco.step[8] ;
 wire \gps_channel0.lo_nco.step[9] ;
 wire \gps_channel0.prompt_i ;
 wire \gps_channel0.prompt_q ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire clknet_4_0_0_wb_clk_i;
 wire clknet_4_1_0_wb_clk_i;
 wire clknet_4_2_0_wb_clk_i;
 wire clknet_4_3_0_wb_clk_i;
 wire clknet_4_4_0_wb_clk_i;
 wire clknet_4_5_0_wb_clk_i;
 wire clknet_4_6_0_wb_clk_i;
 wire clknet_4_7_0_wb_clk_i;
 wire clknet_4_8_0_wb_clk_i;
 wire clknet_4_9_0_wb_clk_i;
 wire clknet_4_10_0_wb_clk_i;
 wire clknet_4_11_0_wb_clk_i;
 wire clknet_4_12_0_wb_clk_i;
 wire clknet_4_13_0_wb_clk_i;
 wire clknet_4_14_0_wb_clk_i;
 wire clknet_4_15_0_wb_clk_i;

 sky130_fd_sc_hd__clkbuf_2 _0956_ (.A(net22),
    .X(_0403_));
 sky130_fd_sc_hd__or2b_1 _0957_ (.A(\gps_channel0.ca_gen.g1[9] ),
    .B_N(_0403_),
    .X(_0404_));
 sky130_fd_sc_hd__clkbuf_1 _0958_ (.A(_0404_),
    .X(_0103_));
 sky130_fd_sc_hd__or2b_1 _0959_ (.A(\gps_channel0.ca_gen.g1[8] ),
    .B_N(_0403_),
    .X(_0405_));
 sky130_fd_sc_hd__clkbuf_1 _0960_ (.A(_0405_),
    .X(_0102_));
 sky130_fd_sc_hd__or2b_1 _0961_ (.A(\gps_channel0.ca_gen.g1[7] ),
    .B_N(_0403_),
    .X(_0406_));
 sky130_fd_sc_hd__clkbuf_1 _0962_ (.A(_0406_),
    .X(_0101_));
 sky130_fd_sc_hd__or2b_1 _0963_ (.A(\gps_channel0.ca_gen.g1[6] ),
    .B_N(_0403_),
    .X(_0407_));
 sky130_fd_sc_hd__clkbuf_1 _0964_ (.A(_0407_),
    .X(_0100_));
 sky130_fd_sc_hd__or2b_1 _0965_ (.A(\gps_channel0.ca_gen.g1[5] ),
    .B_N(_0403_),
    .X(_0408_));
 sky130_fd_sc_hd__clkbuf_1 _0966_ (.A(_0408_),
    .X(_0099_));
 sky130_fd_sc_hd__or2b_1 _0967_ (.A(\gps_channel0.ca_gen.g1[4] ),
    .B_N(_0403_),
    .X(_0409_));
 sky130_fd_sc_hd__clkbuf_1 _0968_ (.A(_0409_),
    .X(_0098_));
 sky130_fd_sc_hd__inv_2 _0969_ (.A(\gps_channel0.ca_gen.g1[3] ),
    .Y(_0410_));
 sky130_fd_sc_hd__nand2_1 _0970_ (.A(_0403_),
    .B(_0410_),
    .Y(_0097_));
 sky130_fd_sc_hd__or2b_1 _0971_ (.A(\gps_channel0.ca_gen.g1[2] ),
    .B_N(_0403_),
    .X(_0411_));
 sky130_fd_sc_hd__clkbuf_1 _0972_ (.A(_0411_),
    .X(_0096_));
 sky130_fd_sc_hd__or2b_1 _0973_ (.A(\gps_channel0.ca_gen.g1[1] ),
    .B_N(_0403_),
    .X(_0412_));
 sky130_fd_sc_hd__clkbuf_1 _0974_ (.A(_0412_),
    .X(_0095_));
 sky130_fd_sc_hd__o21ai_1 _0975_ (.A1(_0410_),
    .A2(\gps_channel0.ca_gen.g1[10] ),
    .B1(_0403_),
    .Y(_0413_));
 sky130_fd_sc_hd__a21o_1 _0976_ (.A1(_0410_),
    .A2(\gps_channel0.ca_gen.g1[10] ),
    .B1(_0413_),
    .X(_0094_));
 sky130_fd_sc_hd__buf_6 _0977_ (.A(net1),
    .X(_0414_));
 sky130_fd_sc_hd__buf_8 _0978_ (.A(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__buf_8 _0979_ (.A(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__inv_2 _0980_ (.A(_0416_),
    .Y(_0797_));
 sky130_fd_sc_hd__inv_2 _0981_ (.A(_0416_),
    .Y(_0798_));
 sky130_fd_sc_hd__inv_2 _0982_ (.A(_0416_),
    .Y(_0799_));
 sky130_fd_sc_hd__inv_2 _0983_ (.A(_0416_),
    .Y(_0800_));
 sky130_fd_sc_hd__inv_2 _0984_ (.A(_0416_),
    .Y(_0801_));
 sky130_fd_sc_hd__inv_2 _0985_ (.A(_0416_),
    .Y(_0802_));
 sky130_fd_sc_hd__inv_2 _0986_ (.A(_0416_),
    .Y(_0803_));
 sky130_fd_sc_hd__inv_2 _0987_ (.A(_0416_),
    .Y(_0804_));
 sky130_fd_sc_hd__inv_2 _0988_ (.A(_0416_),
    .Y(_0805_));
 sky130_fd_sc_hd__inv_2 _0989_ (.A(_0416_),
    .Y(_0806_));
 sky130_fd_sc_hd__buf_8 _0990_ (.A(_0415_),
    .X(_0417_));
 sky130_fd_sc_hd__inv_2 _0991_ (.A(_0417_),
    .Y(_0807_));
 sky130_fd_sc_hd__inv_2 _0992_ (.A(_0417_),
    .Y(_0808_));
 sky130_fd_sc_hd__inv_2 _0993_ (.A(_0417_),
    .Y(_0809_));
 sky130_fd_sc_hd__inv_2 _0994_ (.A(_0417_),
    .Y(_0810_));
 sky130_fd_sc_hd__inv_2 _0995_ (.A(_0417_),
    .Y(_0811_));
 sky130_fd_sc_hd__inv_2 _0996_ (.A(_0417_),
    .Y(_0812_));
 sky130_fd_sc_hd__inv_2 _0997_ (.A(_0417_),
    .Y(_0813_));
 sky130_fd_sc_hd__inv_2 _0998_ (.A(_0417_),
    .Y(_0814_));
 sky130_fd_sc_hd__inv_2 _0999_ (.A(_0417_),
    .Y(_0815_));
 sky130_fd_sc_hd__inv_2 _1000_ (.A(_0417_),
    .Y(_0816_));
 sky130_fd_sc_hd__buf_8 _1001_ (.A(_0414_),
    .X(_0418_));
 sky130_fd_sc_hd__inv_2 _1002_ (.A(_0418_),
    .Y(_0817_));
 sky130_fd_sc_hd__inv_2 _1003_ (.A(_0418_),
    .Y(_0818_));
 sky130_fd_sc_hd__inv_2 _1004_ (.A(_0418_),
    .Y(_0819_));
 sky130_fd_sc_hd__inv_2 _1005_ (.A(_0418_),
    .Y(_0820_));
 sky130_fd_sc_hd__inv_2 _1006_ (.A(_0418_),
    .Y(_0822_));
 sky130_fd_sc_hd__inv_2 _1007_ (.A(_0418_),
    .Y(_0823_));
 sky130_fd_sc_hd__inv_2 _1008_ (.A(_0418_),
    .Y(_0824_));
 sky130_fd_sc_hd__inv_2 _1009_ (.A(_0418_),
    .Y(_0825_));
 sky130_fd_sc_hd__inv_2 _1010_ (.A(_0418_),
    .Y(_0826_));
 sky130_fd_sc_hd__inv_2 _1011_ (.A(_0418_),
    .Y(_0827_));
 sky130_fd_sc_hd__buf_8 _1012_ (.A(_0414_),
    .X(_0419_));
 sky130_fd_sc_hd__inv_2 _1013_ (.A(_0419_),
    .Y(_0828_));
 sky130_fd_sc_hd__inv_2 _1014_ (.A(_0419_),
    .Y(_0829_));
 sky130_fd_sc_hd__inv_2 _1015_ (.A(_0419_),
    .Y(_0830_));
 sky130_fd_sc_hd__inv_2 _1016_ (.A(_0419_),
    .Y(_0831_));
 sky130_fd_sc_hd__inv_2 _1017_ (.A(_0419_),
    .Y(_0832_));
 sky130_fd_sc_hd__inv_2 _1018_ (.A(_0419_),
    .Y(_0833_));
 sky130_fd_sc_hd__inv_2 _1019_ (.A(_0419_),
    .Y(_0834_));
 sky130_fd_sc_hd__inv_2 _1020_ (.A(_0419_),
    .Y(_0835_));
 sky130_fd_sc_hd__inv_2 _1021_ (.A(_0419_),
    .Y(_0836_));
 sky130_fd_sc_hd__inv_2 _1022_ (.A(_0419_),
    .Y(_0837_));
 sky130_fd_sc_hd__buf_8 _1023_ (.A(_0414_),
    .X(_0420_));
 sky130_fd_sc_hd__inv_2 _1024_ (.A(_0420_),
    .Y(_0838_));
 sky130_fd_sc_hd__inv_2 _1025_ (.A(_0420_),
    .Y(_0839_));
 sky130_fd_sc_hd__inv_2 _1026_ (.A(_0420_),
    .Y(_0840_));
 sky130_fd_sc_hd__inv_2 _1027_ (.A(_0420_),
    .Y(_0841_));
 sky130_fd_sc_hd__inv_2 _1028_ (.A(_0420_),
    .Y(_0842_));
 sky130_fd_sc_hd__inv_2 _1029_ (.A(_0420_),
    .Y(_0843_));
 sky130_fd_sc_hd__inv_2 _1030_ (.A(_0420_),
    .Y(_0844_));
 sky130_fd_sc_hd__inv_2 _1031_ (.A(_0420_),
    .Y(_0845_));
 sky130_fd_sc_hd__inv_2 _1032_ (.A(_0420_),
    .Y(_0846_));
 sky130_fd_sc_hd__inv_2 _1033_ (.A(_0420_),
    .Y(_0847_));
 sky130_fd_sc_hd__clkbuf_16 _1034_ (.A(_0414_),
    .X(_0421_));
 sky130_fd_sc_hd__inv_2 _1035_ (.A(_0421_),
    .Y(_0848_));
 sky130_fd_sc_hd__inv_2 _1036_ (.A(_0421_),
    .Y(_0849_));
 sky130_fd_sc_hd__inv_2 _1037_ (.A(_0421_),
    .Y(_0850_));
 sky130_fd_sc_hd__inv_2 _1038_ (.A(_0421_),
    .Y(_0851_));
 sky130_fd_sc_hd__inv_2 _1039_ (.A(_0421_),
    .Y(_0852_));
 sky130_fd_sc_hd__inv_2 _1040_ (.A(_0421_),
    .Y(_0853_));
 sky130_fd_sc_hd__inv_2 _1041_ (.A(_0421_),
    .Y(_0854_));
 sky130_fd_sc_hd__inv_2 _1042_ (.A(_0421_),
    .Y(_0855_));
 sky130_fd_sc_hd__inv_2 _1043_ (.A(_0421_),
    .Y(_0856_));
 sky130_fd_sc_hd__inv_2 _1044_ (.A(_0421_),
    .Y(_0751_));
 sky130_fd_sc_hd__buf_8 _1045_ (.A(_0414_),
    .X(_0422_));
 sky130_fd_sc_hd__inv_2 _1046_ (.A(_0422_),
    .Y(_0857_));
 sky130_fd_sc_hd__inv_2 _1047_ (.A(_0422_),
    .Y(_0752_));
 sky130_fd_sc_hd__inv_2 _1048_ (.A(_0422_),
    .Y(_0858_));
 sky130_fd_sc_hd__inv_2 _1049_ (.A(_0422_),
    .Y(_0753_));
 sky130_fd_sc_hd__inv_2 _1050_ (.A(_0422_),
    .Y(_0754_));
 sky130_fd_sc_hd__inv_2 _1051_ (.A(_0422_),
    .Y(_0755_));
 sky130_fd_sc_hd__inv_2 _1052_ (.A(_0422_),
    .Y(_0756_));
 sky130_fd_sc_hd__inv_2 _1053_ (.A(_0422_),
    .Y(_0757_));
 sky130_fd_sc_hd__inv_2 _1054_ (.A(_0422_),
    .Y(_0758_));
 sky130_fd_sc_hd__inv_2 _1055_ (.A(_0422_),
    .Y(_0759_));
 sky130_fd_sc_hd__buf_6 _1056_ (.A(_0414_),
    .X(_0423_));
 sky130_fd_sc_hd__inv_2 _1057_ (.A(_0423_),
    .Y(_0760_));
 sky130_fd_sc_hd__inv_2 _1058_ (.A(_0423_),
    .Y(_0761_));
 sky130_fd_sc_hd__inv_2 _1059_ (.A(_0423_),
    .Y(_0762_));
 sky130_fd_sc_hd__inv_2 _1060_ (.A(_0423_),
    .Y(_0763_));
 sky130_fd_sc_hd__inv_2 _1061_ (.A(_0423_),
    .Y(_0764_));
 sky130_fd_sc_hd__inv_2 _1062_ (.A(_0423_),
    .Y(_0765_));
 sky130_fd_sc_hd__inv_2 _1063_ (.A(_0423_),
    .Y(_0766_));
 sky130_fd_sc_hd__inv_2 _1064_ (.A(_0423_),
    .Y(_0767_));
 sky130_fd_sc_hd__inv_2 _1065_ (.A(_0423_),
    .Y(_0768_));
 sky130_fd_sc_hd__inv_2 _1066_ (.A(_0423_),
    .Y(_0769_));
 sky130_fd_sc_hd__clkbuf_16 _1067_ (.A(_0414_),
    .X(_0424_));
 sky130_fd_sc_hd__inv_2 _1068_ (.A(_0424_),
    .Y(_0770_));
 sky130_fd_sc_hd__inv_2 _1069_ (.A(_0424_),
    .Y(_0771_));
 sky130_fd_sc_hd__inv_2 _1070_ (.A(_0424_),
    .Y(_0772_));
 sky130_fd_sc_hd__inv_2 _1071_ (.A(_0424_),
    .Y(_0773_));
 sky130_fd_sc_hd__inv_2 _1072_ (.A(_0424_),
    .Y(_0774_));
 sky130_fd_sc_hd__inv_2 _1073_ (.A(_0424_),
    .Y(_0775_));
 sky130_fd_sc_hd__inv_2 _1074_ (.A(_0424_),
    .Y(_0776_));
 sky130_fd_sc_hd__inv_2 _1075_ (.A(_0424_),
    .Y(_0777_));
 sky130_fd_sc_hd__inv_2 _1076_ (.A(_0424_),
    .Y(_0778_));
 sky130_fd_sc_hd__inv_2 _1077_ (.A(_0424_),
    .Y(_0779_));
 sky130_fd_sc_hd__buf_8 _1078_ (.A(_0414_),
    .X(_0425_));
 sky130_fd_sc_hd__inv_2 _1079_ (.A(_0425_),
    .Y(_0780_));
 sky130_fd_sc_hd__inv_2 _1080_ (.A(_0425_),
    .Y(_0781_));
 sky130_fd_sc_hd__inv_2 _1081_ (.A(_0425_),
    .Y(_0787_));
 sky130_fd_sc_hd__inv_2 _1082_ (.A(_0425_),
    .Y(_0784_));
 sky130_fd_sc_hd__inv_2 _1083_ (.A(_0425_),
    .Y(_0782_));
 sky130_fd_sc_hd__inv_2 _1084_ (.A(_0425_),
    .Y(_0785_));
 sky130_fd_sc_hd__inv_2 _1085_ (.A(_0425_),
    .Y(_0791_));
 sky130_fd_sc_hd__inv_2 _1086_ (.A(_0425_),
    .Y(_0792_));
 sky130_fd_sc_hd__inv_2 _1087_ (.A(_0425_),
    .Y(_0793_));
 sky130_fd_sc_hd__inv_2 _1088_ (.A(_0425_),
    .Y(_0789_));
 sky130_fd_sc_hd__inv_2 _1089_ (.A(_0415_),
    .Y(_0790_));
 sky130_fd_sc_hd__inv_2 _1090_ (.A(_0415_),
    .Y(_0788_));
 sky130_fd_sc_hd__inv_2 _1091_ (.A(_0415_),
    .Y(_0786_));
 sky130_fd_sc_hd__inv_2 _1092_ (.A(_0415_),
    .Y(_0794_));
 sky130_fd_sc_hd__inv_2 _1093_ (.A(_0415_),
    .Y(_0795_));
 sky130_fd_sc_hd__inv_2 _1094_ (.A(_0415_),
    .Y(_0796_));
 sky130_fd_sc_hd__inv_2 _1095_ (.A(_0415_),
    .Y(_0821_));
 sky130_fd_sc_hd__inv_2 _1096_ (.A(_0415_),
    .Y(_0783_));
 sky130_fd_sc_hd__xnor2_1 _1097_ (.A(\gps_channel0.ca_gen.g2[10] ),
    .B(\gps_channel0.ca_gen.g2[9] ),
    .Y(_0426_));
 sky130_fd_sc_hd__xnor2_1 _1098_ (.A(\gps_channel0.ca_gen.g2[3] ),
    .B(\gps_channel0.ca_gen.g2[2] ),
    .Y(_0427_));
 sky130_fd_sc_hd__xor2_1 _1099_ (.A(\gps_channel0.ca_gen.g2[8] ),
    .B(\gps_channel0.ca_gen.g2[6] ),
    .X(_0428_));
 sky130_fd_sc_hd__xnor2_1 _1100_ (.A(_0427_),
    .B(_0428_),
    .Y(_0429_));
 sky130_fd_sc_hd__xnor2_1 _1101_ (.A(_0426_),
    .B(_0429_),
    .Y(_0430_));
 sky130_fd_sc_hd__clkbuf_4 _1102_ (.A(net22),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _1103_ (.A0(\gps_channel0.ca_gen.g2_init[1] ),
    .A1(_0430_),
    .S(_0431_),
    .X(_0432_));
 sky130_fd_sc_hd__clkbuf_1 _1104_ (.A(_0432_),
    .X(_0000_));
 sky130_fd_sc_hd__mux2_1 _1105_ (.A0(\gps_channel0.ca_gen.g2_init[2] ),
    .A1(\gps_channel0.ca_gen.g2[1] ),
    .S(_0431_),
    .X(_0433_));
 sky130_fd_sc_hd__clkbuf_1 _1106_ (.A(_0433_),
    .X(_0001_));
 sky130_fd_sc_hd__mux2_1 _1107_ (.A0(\gps_channel0.ca_gen.g2_init[3] ),
    .A1(\gps_channel0.ca_gen.g2[2] ),
    .S(_0431_),
    .X(_0434_));
 sky130_fd_sc_hd__clkbuf_1 _1108_ (.A(_0434_),
    .X(_0002_));
 sky130_fd_sc_hd__mux2_1 _1109_ (.A0(\gps_channel0.ca_gen.g2_init[4] ),
    .A1(\gps_channel0.ca_gen.g2[3] ),
    .S(_0431_),
    .X(_0435_));
 sky130_fd_sc_hd__clkbuf_1 _1110_ (.A(_0435_),
    .X(_0003_));
 sky130_fd_sc_hd__mux2_1 _1111_ (.A0(\gps_channel0.ca_gen.g2_init[5] ),
    .A1(\gps_channel0.ca_gen.g2[4] ),
    .S(_0431_),
    .X(_0436_));
 sky130_fd_sc_hd__clkbuf_1 _1112_ (.A(_0436_),
    .X(_0004_));
 sky130_fd_sc_hd__mux2_1 _1113_ (.A0(\gps_channel0.ca_gen.g2_init[6] ),
    .A1(\gps_channel0.ca_gen.g2[5] ),
    .S(_0431_),
    .X(_0437_));
 sky130_fd_sc_hd__clkbuf_1 _1114_ (.A(_0437_),
    .X(_0005_));
 sky130_fd_sc_hd__mux2_1 _1115_ (.A0(\gps_channel0.ca_gen.g2_init[7] ),
    .A1(\gps_channel0.ca_gen.g2[6] ),
    .S(_0431_),
    .X(_0438_));
 sky130_fd_sc_hd__clkbuf_1 _1116_ (.A(_0438_),
    .X(_0006_));
 sky130_fd_sc_hd__mux2_1 _1117_ (.A0(\gps_channel0.ca_gen.g2_init[8] ),
    .A1(\gps_channel0.ca_gen.g2[7] ),
    .S(_0431_),
    .X(_0439_));
 sky130_fd_sc_hd__clkbuf_1 _1118_ (.A(_0439_),
    .X(_0007_));
 sky130_fd_sc_hd__mux2_1 _1119_ (.A0(\gps_channel0.ca_gen.g2_init[9] ),
    .A1(\gps_channel0.ca_gen.g2[8] ),
    .S(_0431_),
    .X(_0440_));
 sky130_fd_sc_hd__clkbuf_1 _1120_ (.A(_0440_),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_1 _1121_ (.A0(\gps_channel0.ca_gen.g2_init[10] ),
    .A1(\gps_channel0.ca_gen.g2[9] ),
    .S(_0431_),
    .X(_0441_));
 sky130_fd_sc_hd__clkbuf_1 _1122_ (.A(_0441_),
    .X(_0009_));
 sky130_fd_sc_hd__xnor2_1 _1123_ (.A(\gps_channel0.ca_gen.g1[10] ),
    .B(net2),
    .Y(_0442_));
 sky130_fd_sc_hd__xor2_1 _1124_ (.A(\gps_channel0.ca_gen.g2[10] ),
    .B(\gps_channel0.lo_i ),
    .X(_0443_));
 sky130_fd_sc_hd__xnor2_1 _1125_ (.A(_0442_),
    .B(_0443_),
    .Y(\gps_channel0.prompt_i ));
 sky130_fd_sc_hd__xor2_1 _1126_ (.A(\gps_channel0.lo_nco.accumulator[30] ),
    .B(\gps_channel0.prompt_i ),
    .X(\gps_channel0.prompt_q ));
 sky130_fd_sc_hd__nand2_1 _1127_ (.A(\gps_channel0.lo_nco.step[0] ),
    .B(net8),
    .Y(_0444_));
 sky130_fd_sc_hd__xnor2_1 _1128_ (.A(\gps_channel0.lo_nco.accumulator[0] ),
    .B(_0444_),
    .Y(_0445_));
 sky130_fd_sc_hd__nor2_4 _1129_ (.A(\gps_channel0.lo_nco.phase_sync ),
    .B(net3),
    .Y(_0446_));
 sky130_fd_sc_hd__clkbuf_4 _1130_ (.A(_0446_),
    .X(_0447_));
 sky130_fd_sc_hd__mux2_1 _1131_ (.A0(\gps_channel0.lo_nco.phase_in[0] ),
    .A1(_0445_),
    .S(_0447_),
    .X(_0448_));
 sky130_fd_sc_hd__clkbuf_1 _1132_ (.A(_0448_),
    .X(_0030_));
 sky130_fd_sc_hd__or2_1 _1133_ (.A(\gps_channel0.lo_nco.phase_sync ),
    .B(net3),
    .X(_0449_));
 sky130_fd_sc_hd__buf_4 _1134_ (.A(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__nor2_4 _1135_ (.A(net8),
    .B(_0450_),
    .Y(_0451_));
 sky130_fd_sc_hd__xor2_1 _1136_ (.A(\gps_channel0.lo_nco.step[1] ),
    .B(\gps_channel0.lo_nco.accumulator[1] ),
    .X(_0452_));
 sky130_fd_sc_hd__a21oi_1 _1137_ (.A1(\gps_channel0.lo_nco.step[0] ),
    .A2(\gps_channel0.lo_nco.accumulator[0] ),
    .B1(_0452_),
    .Y(_0453_));
 sky130_fd_sc_hd__nand2_4 _1138_ (.A(net8),
    .B(_0446_),
    .Y(_0454_));
 sky130_fd_sc_hd__a31o_1 _1139_ (.A1(\gps_channel0.lo_nco.step[0] ),
    .A2(\gps_channel0.lo_nco.accumulator[0] ),
    .A3(_0452_),
    .B1(_0454_),
    .X(_0455_));
 sky130_fd_sc_hd__nor2_1 _1140_ (.A(_0453_),
    .B(_0455_),
    .Y(_0456_));
 sky130_fd_sc_hd__a221o_1 _1141_ (.A1(\gps_channel0.lo_nco.phase_in[1] ),
    .A2(_0450_),
    .B1(_0451_),
    .B2(\gps_channel0.lo_nco.accumulator[1] ),
    .C1(_0456_),
    .X(_0031_));
 sky130_fd_sc_hd__or2_1 _1142_ (.A(net8),
    .B(_0450_),
    .X(_0457_));
 sky130_fd_sc_hd__clkbuf_4 _1143_ (.A(_0457_),
    .X(_0458_));
 sky130_fd_sc_hd__and2_1 _1144_ (.A(\gps_channel0.lo_nco.step[1] ),
    .B(\gps_channel0.lo_nco.accumulator[1] ),
    .X(_0459_));
 sky130_fd_sc_hd__a31oi_2 _1145_ (.A1(\gps_channel0.lo_nco.step[0] ),
    .A2(\gps_channel0.lo_nco.accumulator[0] ),
    .A3(_0452_),
    .B1(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__or2_1 _1146_ (.A(\gps_channel0.lo_nco.step[2] ),
    .B(\gps_channel0.lo_nco.accumulator[2] ),
    .X(_0461_));
 sky130_fd_sc_hd__nand2_1 _1147_ (.A(\gps_channel0.lo_nco.step[2] ),
    .B(\gps_channel0.lo_nco.accumulator[2] ),
    .Y(_0462_));
 sky130_fd_sc_hd__nand2_1 _1148_ (.A(_0461_),
    .B(_0462_),
    .Y(_0463_));
 sky130_fd_sc_hd__or2_1 _1149_ (.A(_0460_),
    .B(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__nand2_1 _1150_ (.A(_0460_),
    .B(_0463_),
    .Y(_0465_));
 sky130_fd_sc_hd__a21o_1 _1151_ (.A1(_0464_),
    .A2(_0465_),
    .B1(_0454_),
    .X(_0466_));
 sky130_fd_sc_hd__o221a_1 _1152_ (.A1(\gps_channel0.lo_nco.phase_in[2] ),
    .A2(_0447_),
    .B1(_0458_),
    .B2(\gps_channel0.lo_nco.accumulator[2] ),
    .C1(_0466_),
    .X(_0032_));
 sky130_fd_sc_hd__or2_1 _1153_ (.A(\gps_channel0.lo_nco.step[3] ),
    .B(\gps_channel0.lo_nco.accumulator[3] ),
    .X(_0467_));
 sky130_fd_sc_hd__nand2_1 _1154_ (.A(\gps_channel0.lo_nco.step[3] ),
    .B(\gps_channel0.lo_nco.accumulator[3] ),
    .Y(_0468_));
 sky130_fd_sc_hd__nand2_1 _1155_ (.A(_0467_),
    .B(_0468_),
    .Y(_0469_));
 sky130_fd_sc_hd__o21ai_1 _1156_ (.A1(_0460_),
    .A2(_0463_),
    .B1(_0462_),
    .Y(_0470_));
 sky130_fd_sc_hd__xnor2_1 _1157_ (.A(_0469_),
    .B(_0470_),
    .Y(_0471_));
 sky130_fd_sc_hd__mux2_1 _1158_ (.A0(\gps_channel0.lo_nco.phase_in[3] ),
    .A1(_0471_),
    .S(_0446_),
    .X(_0472_));
 sky130_fd_sc_hd__mux2_1 _1159_ (.A0(\gps_channel0.lo_nco.accumulator[3] ),
    .A1(_0472_),
    .S(_0458_),
    .X(_0473_));
 sky130_fd_sc_hd__clkbuf_1 _1160_ (.A(_0473_),
    .X(_0033_));
 sky130_fd_sc_hd__nand2_1 _1161_ (.A(\gps_channel0.lo_nco.step[4] ),
    .B(\gps_channel0.lo_nco.accumulator[4] ),
    .Y(_0474_));
 sky130_fd_sc_hd__or2_1 _1162_ (.A(\gps_channel0.lo_nco.step[4] ),
    .B(\gps_channel0.lo_nco.accumulator[4] ),
    .X(_0475_));
 sky130_fd_sc_hd__nand2_1 _1163_ (.A(_0474_),
    .B(_0475_),
    .Y(_0476_));
 sky130_fd_sc_hd__nand3_1 _1164_ (.A(\gps_channel0.lo_nco.step[2] ),
    .B(\gps_channel0.lo_nco.accumulator[2] ),
    .C(_0467_),
    .Y(_0477_));
 sky130_fd_sc_hd__o311a_1 _1165_ (.A1(_0460_),
    .A2(_0463_),
    .A3(_0469_),
    .B1(_0477_),
    .C1(_0468_),
    .X(_0478_));
 sky130_fd_sc_hd__xor2_1 _1166_ (.A(_0476_),
    .B(_0478_),
    .X(_0479_));
 sky130_fd_sc_hd__or2_1 _1167_ (.A(\gps_channel0.lo_nco.phase_in[4] ),
    .B(_0447_),
    .X(_0480_));
 sky130_fd_sc_hd__o221a_1 _1168_ (.A1(\gps_channel0.lo_nco.accumulator[4] ),
    .A2(_0458_),
    .B1(_0479_),
    .B2(_0454_),
    .C1(_0480_),
    .X(_0034_));
 sky130_fd_sc_hd__o21a_1 _1169_ (.A1(_0476_),
    .A2(_0478_),
    .B1(_0474_),
    .X(_0481_));
 sky130_fd_sc_hd__nor2_1 _1170_ (.A(\gps_channel0.lo_nco.step[5] ),
    .B(\gps_channel0.lo_nco.accumulator[5] ),
    .Y(_0482_));
 sky130_fd_sc_hd__nand2_1 _1171_ (.A(\gps_channel0.lo_nco.step[5] ),
    .B(\gps_channel0.lo_nco.accumulator[5] ),
    .Y(_0483_));
 sky130_fd_sc_hd__and2b_1 _1172_ (.A_N(_0482_),
    .B(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__and2_1 _1173_ (.A(net8),
    .B(_0446_),
    .X(_0485_));
 sky130_fd_sc_hd__clkbuf_2 _1174_ (.A(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__o21ai_1 _1175_ (.A1(_0481_),
    .A2(_0484_),
    .B1(_0486_),
    .Y(_0487_));
 sky130_fd_sc_hd__a21o_1 _1176_ (.A1(_0481_),
    .A2(_0484_),
    .B1(_0487_),
    .X(_0488_));
 sky130_fd_sc_hd__o221a_1 _1177_ (.A1(\gps_channel0.lo_nco.phase_in[5] ),
    .A2(_0447_),
    .B1(_0458_),
    .B2(\gps_channel0.lo_nco.accumulator[5] ),
    .C1(_0488_),
    .X(_0035_));
 sky130_fd_sc_hd__xor2_1 _1178_ (.A(\gps_channel0.lo_nco.step[6] ),
    .B(\gps_channel0.lo_nco.accumulator[6] ),
    .X(_0489_));
 sky130_fd_sc_hd__a21oi_1 _1179_ (.A1(_0481_),
    .A2(_0483_),
    .B1(_0482_),
    .Y(_0490_));
 sky130_fd_sc_hd__or2_1 _1180_ (.A(_0489_),
    .B(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__a21oi_1 _1181_ (.A1(_0489_),
    .A2(_0490_),
    .B1(_0454_),
    .Y(_0492_));
 sky130_fd_sc_hd__a22o_1 _1182_ (.A1(\gps_channel0.lo_nco.phase_in[6] ),
    .A2(_0450_),
    .B1(_0451_),
    .B2(\gps_channel0.lo_nco.accumulator[6] ),
    .X(_0493_));
 sky130_fd_sc_hd__a21o_1 _1183_ (.A1(_0491_),
    .A2(_0492_),
    .B1(_0493_),
    .X(_0036_));
 sky130_fd_sc_hd__nor2_1 _1184_ (.A(\gps_channel0.lo_nco.step[7] ),
    .B(\gps_channel0.lo_nco.accumulator[7] ),
    .Y(_0494_));
 sky130_fd_sc_hd__nand2_1 _1185_ (.A(\gps_channel0.lo_nco.step[7] ),
    .B(\gps_channel0.lo_nco.accumulator[7] ),
    .Y(_0495_));
 sky130_fd_sc_hd__and2b_1 _1186_ (.A_N(_0494_),
    .B(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__a22o_1 _1187_ (.A1(\gps_channel0.lo_nco.step[6] ),
    .A2(\gps_channel0.lo_nco.accumulator[6] ),
    .B1(_0489_),
    .B2(_0490_),
    .X(_0497_));
 sky130_fd_sc_hd__xor2_1 _1188_ (.A(_0496_),
    .B(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _1189_ (.A0(\gps_channel0.lo_nco.phase_in[7] ),
    .A1(_0498_),
    .S(_0446_),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_1 _1190_ (.A0(\gps_channel0.lo_nco.accumulator[7] ),
    .A1(_0499_),
    .S(_0458_),
    .X(_0500_));
 sky130_fd_sc_hd__clkbuf_1 _1191_ (.A(_0500_),
    .X(_0037_));
 sky130_fd_sc_hd__clkbuf_4 _1192_ (.A(_0486_),
    .X(_0501_));
 sky130_fd_sc_hd__nand3b_1 _1193_ (.A_N(_0494_),
    .B(\gps_channel0.lo_nco.accumulator[6] ),
    .C(\gps_channel0.lo_nco.step[6] ),
    .Y(_0502_));
 sky130_fd_sc_hd__and3b_1 _1194_ (.A_N(_0494_),
    .B(_0495_),
    .C(_0489_),
    .X(_0503_));
 sky130_fd_sc_hd__nand3b_1 _1195_ (.A_N(_0476_),
    .B(_0484_),
    .C(_0503_),
    .Y(_0504_));
 sky130_fd_sc_hd__a21oi_1 _1196_ (.A1(_0474_),
    .A2(_0483_),
    .B1(_0482_),
    .Y(_0505_));
 sky130_fd_sc_hd__nand2_1 _1197_ (.A(_0505_),
    .B(_0503_),
    .Y(_0506_));
 sky130_fd_sc_hd__o211a_1 _1198_ (.A1(_0478_),
    .A2(_0504_),
    .B1(_0506_),
    .C1(_0495_),
    .X(_0507_));
 sky130_fd_sc_hd__nand2_1 _1199_ (.A(_0502_),
    .B(_0507_),
    .Y(_0508_));
 sky130_fd_sc_hd__nand2_1 _1200_ (.A(\gps_channel0.lo_nco.step[8] ),
    .B(\gps_channel0.lo_nco.accumulator[8] ),
    .Y(_0509_));
 sky130_fd_sc_hd__or2_1 _1201_ (.A(\gps_channel0.lo_nco.step[8] ),
    .B(\gps_channel0.lo_nco.accumulator[8] ),
    .X(_0510_));
 sky130_fd_sc_hd__nand2_1 _1202_ (.A(_0509_),
    .B(_0510_),
    .Y(_0511_));
 sky130_fd_sc_hd__xor2_1 _1203_ (.A(_0508_),
    .B(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__nand2_1 _1204_ (.A(_0501_),
    .B(_0512_),
    .Y(_0513_));
 sky130_fd_sc_hd__o221a_1 _1205_ (.A1(\gps_channel0.lo_nco.phase_in[8] ),
    .A2(_0447_),
    .B1(_0458_),
    .B2(\gps_channel0.lo_nco.accumulator[8] ),
    .C1(_0513_),
    .X(_0038_));
 sky130_fd_sc_hd__a21bo_1 _1206_ (.A1(_0508_),
    .A2(_0510_),
    .B1_N(_0509_),
    .X(_0514_));
 sky130_fd_sc_hd__or2_1 _1207_ (.A(\gps_channel0.lo_nco.step[9] ),
    .B(\gps_channel0.lo_nco.accumulator[9] ),
    .X(_0515_));
 sky130_fd_sc_hd__nand2_1 _1208_ (.A(\gps_channel0.lo_nco.step[9] ),
    .B(\gps_channel0.lo_nco.accumulator[9] ),
    .Y(_0516_));
 sky130_fd_sc_hd__nand2_1 _1209_ (.A(_0515_),
    .B(_0516_),
    .Y(_0517_));
 sky130_fd_sc_hd__xnor2_1 _1210_ (.A(_0514_),
    .B(_0517_),
    .Y(_0518_));
 sky130_fd_sc_hd__or2_1 _1211_ (.A(\gps_channel0.lo_nco.phase_in[9] ),
    .B(_0447_),
    .X(_0519_));
 sky130_fd_sc_hd__o221a_1 _1212_ (.A1(\gps_channel0.lo_nco.accumulator[9] ),
    .A2(_0458_),
    .B1(_0518_),
    .B2(_0454_),
    .C1(_0519_),
    .X(_0039_));
 sky130_fd_sc_hd__or2b_1 _1213_ (.A(_0514_),
    .B_N(_0516_),
    .X(_0520_));
 sky130_fd_sc_hd__xor2_1 _1214_ (.A(\gps_channel0.lo_nco.step[10] ),
    .B(\gps_channel0.lo_nco.accumulator[10] ),
    .X(_0521_));
 sky130_fd_sc_hd__a21oi_1 _1215_ (.A1(_0515_),
    .A2(_0520_),
    .B1(_0521_),
    .Y(_0522_));
 sky130_fd_sc_hd__and3_1 _1216_ (.A(_0515_),
    .B(_0520_),
    .C(_0521_),
    .X(_0523_));
 sky130_fd_sc_hd__nor3_1 _1217_ (.A(_0454_),
    .B(_0522_),
    .C(_0523_),
    .Y(_0524_));
 sky130_fd_sc_hd__a221o_1 _1218_ (.A1(\gps_channel0.lo_nco.phase_in[10] ),
    .A2(_0450_),
    .B1(_0451_),
    .B2(\gps_channel0.lo_nco.accumulator[10] ),
    .C1(_0524_),
    .X(_0040_));
 sky130_fd_sc_hd__clkbuf_4 _1219_ (.A(_0451_),
    .X(_0525_));
 sky130_fd_sc_hd__nor2_1 _1220_ (.A(\gps_channel0.lo_nco.step[11] ),
    .B(\gps_channel0.lo_nco.accumulator[11] ),
    .Y(_0526_));
 sky130_fd_sc_hd__and2_1 _1221_ (.A(\gps_channel0.lo_nco.step[11] ),
    .B(\gps_channel0.lo_nco.accumulator[11] ),
    .X(_0527_));
 sky130_fd_sc_hd__nor2_1 _1222_ (.A(_0526_),
    .B(_0527_),
    .Y(_0528_));
 sky130_fd_sc_hd__a21o_1 _1223_ (.A1(\gps_channel0.lo_nco.step[10] ),
    .A2(\gps_channel0.lo_nco.accumulator[10] ),
    .B1(_0523_),
    .X(_0529_));
 sky130_fd_sc_hd__xnor2_1 _1224_ (.A(_0528_),
    .B(_0529_),
    .Y(_0530_));
 sky130_fd_sc_hd__nand2_1 _1225_ (.A(_0447_),
    .B(_0530_),
    .Y(_0531_));
 sky130_fd_sc_hd__o21a_1 _1226_ (.A1(\gps_channel0.lo_nco.phase_in[11] ),
    .A2(_0447_),
    .B1(_0458_),
    .X(_0532_));
 sky130_fd_sc_hd__a22o_1 _1227_ (.A1(\gps_channel0.lo_nco.accumulator[11] ),
    .A2(_0525_),
    .B1(_0531_),
    .B2(_0532_),
    .X(_0041_));
 sky130_fd_sc_hd__nand2_1 _1228_ (.A(_0521_),
    .B(_0528_),
    .Y(_0533_));
 sky130_fd_sc_hd__or3_1 _1229_ (.A(_0511_),
    .B(_0517_),
    .C(_0533_),
    .X(_0534_));
 sky130_fd_sc_hd__a21o_1 _1230_ (.A1(_0502_),
    .A2(_0507_),
    .B1(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__and2_1 _1231_ (.A(_0509_),
    .B(_0516_),
    .X(_0536_));
 sky130_fd_sc_hd__or3b_1 _1232_ (.A(_0533_),
    .B(_0536_),
    .C_N(_0515_),
    .X(_0537_));
 sky130_fd_sc_hd__nand3b_1 _1233_ (.A_N(_0526_),
    .B(\gps_channel0.lo_nco.accumulator[10] ),
    .C(\gps_channel0.lo_nco.step[10] ),
    .Y(_0538_));
 sky130_fd_sc_hd__and3b_1 _1234_ (.A_N(_0527_),
    .B(_0537_),
    .C(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__nand2_1 _1235_ (.A(_0535_),
    .B(_0539_),
    .Y(_0540_));
 sky130_fd_sc_hd__nand2_1 _1236_ (.A(\gps_channel0.lo_nco.step[12] ),
    .B(\gps_channel0.lo_nco.accumulator[12] ),
    .Y(_0541_));
 sky130_fd_sc_hd__or2_1 _1237_ (.A(\gps_channel0.lo_nco.step[12] ),
    .B(\gps_channel0.lo_nco.accumulator[12] ),
    .X(_0542_));
 sky130_fd_sc_hd__nand2_1 _1238_ (.A(_0541_),
    .B(_0542_),
    .Y(_0543_));
 sky130_fd_sc_hd__xor2_1 _1239_ (.A(_0540_),
    .B(_0543_),
    .X(_0544_));
 sky130_fd_sc_hd__nand2_1 _1240_ (.A(_0501_),
    .B(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__o221a_1 _1241_ (.A1(\gps_channel0.lo_nco.phase_in[12] ),
    .A2(_0447_),
    .B1(_0458_),
    .B2(\gps_channel0.lo_nco.accumulator[12] ),
    .C1(_0545_),
    .X(_0042_));
 sky130_fd_sc_hd__a21bo_1 _1242_ (.A1(_0540_),
    .A2(_0542_),
    .B1_N(_0541_),
    .X(_0546_));
 sky130_fd_sc_hd__nor2_1 _1243_ (.A(\gps_channel0.lo_nco.step[13] ),
    .B(\gps_channel0.lo_nco.accumulator[13] ),
    .Y(_0547_));
 sky130_fd_sc_hd__nand2_1 _1244_ (.A(\gps_channel0.lo_nco.step[13] ),
    .B(\gps_channel0.lo_nco.accumulator[13] ),
    .Y(_0548_));
 sky130_fd_sc_hd__or2b_1 _1245_ (.A(_0547_),
    .B_N(_0548_),
    .X(_0549_));
 sky130_fd_sc_hd__xnor2_1 _1246_ (.A(_0546_),
    .B(_0549_),
    .Y(_0550_));
 sky130_fd_sc_hd__or2_1 _1247_ (.A(\gps_channel0.lo_nco.phase_in[13] ),
    .B(_0447_),
    .X(_0551_));
 sky130_fd_sc_hd__o221a_1 _1248_ (.A1(\gps_channel0.lo_nco.accumulator[13] ),
    .A2(_0458_),
    .B1(_0550_),
    .B2(_0454_),
    .C1(_0551_),
    .X(_0043_));
 sky130_fd_sc_hd__and2b_1 _1249_ (.A_N(_0546_),
    .B(_0548_),
    .X(_0552_));
 sky130_fd_sc_hd__or2_1 _1250_ (.A(\gps_channel0.lo_nco.step[14] ),
    .B(\gps_channel0.lo_nco.accumulator[14] ),
    .X(_0553_));
 sky130_fd_sc_hd__nand2_1 _1251_ (.A(\gps_channel0.lo_nco.step[14] ),
    .B(\gps_channel0.lo_nco.accumulator[14] ),
    .Y(_0554_));
 sky130_fd_sc_hd__nand2_1 _1252_ (.A(_0553_),
    .B(_0554_),
    .Y(_0555_));
 sky130_fd_sc_hd__o21ai_1 _1253_ (.A1(_0547_),
    .A2(_0552_),
    .B1(_0555_),
    .Y(_0556_));
 sky130_fd_sc_hd__or3_1 _1254_ (.A(_0547_),
    .B(_0552_),
    .C(_0555_),
    .X(_0557_));
 sky130_fd_sc_hd__a22o_1 _1255_ (.A1(\gps_channel0.lo_nco.phase_in[14] ),
    .A2(_0450_),
    .B1(_0451_),
    .B2(\gps_channel0.lo_nco.accumulator[14] ),
    .X(_0558_));
 sky130_fd_sc_hd__a31o_1 _1256_ (.A1(_0501_),
    .A2(_0556_),
    .A3(_0557_),
    .B1(_0558_),
    .X(_0044_));
 sky130_fd_sc_hd__nor2_1 _1257_ (.A(\gps_channel0.lo_nco.step[15] ),
    .B(\gps_channel0.lo_nco.accumulator[15] ),
    .Y(_0559_));
 sky130_fd_sc_hd__and2_1 _1258_ (.A(\gps_channel0.lo_nco.step[15] ),
    .B(\gps_channel0.lo_nco.accumulator[15] ),
    .X(_0560_));
 sky130_fd_sc_hd__nor2_1 _1259_ (.A(_0559_),
    .B(_0560_),
    .Y(_0561_));
 sky130_fd_sc_hd__a21oi_1 _1260_ (.A1(_0554_),
    .A2(_0557_),
    .B1(_0561_),
    .Y(_0562_));
 sky130_fd_sc_hd__a31o_1 _1261_ (.A1(_0554_),
    .A2(_0557_),
    .A3(_0561_),
    .B1(_0450_),
    .X(_0563_));
 sky130_fd_sc_hd__o22a_1 _1262_ (.A1(\gps_channel0.lo_nco.phase_in[15] ),
    .A2(_0446_),
    .B1(_0562_),
    .B2(_0563_),
    .X(_0564_));
 sky130_fd_sc_hd__mux2_1 _1263_ (.A0(\gps_channel0.lo_nco.accumulator[15] ),
    .A1(_0564_),
    .S(_0457_),
    .X(_0565_));
 sky130_fd_sc_hd__clkbuf_1 _1264_ (.A(_0565_),
    .X(_0045_));
 sky130_fd_sc_hd__nor2_1 _1265_ (.A(\gps_channel0.ca_nco.step[11] ),
    .B(\gps_channel0.ca_nco.accumulator[11] ),
    .Y(_0566_));
 sky130_fd_sc_hd__nand2_1 _1266_ (.A(\gps_channel0.ca_nco.step[10] ),
    .B(\gps_channel0.ca_nco.accumulator[10] ),
    .Y(_0567_));
 sky130_fd_sc_hd__nand2_1 _1267_ (.A(\gps_channel0.ca_nco.step[11] ),
    .B(\gps_channel0.ca_nco.accumulator[11] ),
    .Y(_0568_));
 sky130_fd_sc_hd__or2b_1 _1268_ (.A(_0566_),
    .B_N(_0568_),
    .X(_0569_));
 sky130_fd_sc_hd__or2_1 _1269_ (.A(\gps_channel0.ca_nco.step[10] ),
    .B(\gps_channel0.ca_nco.accumulator[10] ),
    .X(_0570_));
 sky130_fd_sc_hd__nand2_1 _1270_ (.A(_0567_),
    .B(_0570_),
    .Y(_0571_));
 sky130_fd_sc_hd__or2_1 _1271_ (.A(_0569_),
    .B(_0571_),
    .X(_0572_));
 sky130_fd_sc_hd__nand2_1 _1272_ (.A(\gps_channel0.ca_nco.step[9] ),
    .B(\gps_channel0.ca_nco.accumulator[9] ),
    .Y(_0573_));
 sky130_fd_sc_hd__nand2_1 _1273_ (.A(\gps_channel0.ca_nco.step[8] ),
    .B(\gps_channel0.ca_nco.accumulator[8] ),
    .Y(_0574_));
 sky130_fd_sc_hd__nor2_1 _1274_ (.A(\gps_channel0.ca_nco.step[9] ),
    .B(\gps_channel0.ca_nco.accumulator[9] ),
    .Y(_0575_));
 sky130_fd_sc_hd__a21o_1 _1275_ (.A1(_0573_),
    .A2(_0574_),
    .B1(_0575_),
    .X(_0576_));
 sky130_fd_sc_hd__o221a_1 _1276_ (.A1(_0566_),
    .A2(_0567_),
    .B1(_0572_),
    .B2(_0576_),
    .C1(_0568_),
    .X(_0577_));
 sky130_fd_sc_hd__nand2_1 _1277_ (.A(\gps_channel0.ca_nco.step[3] ),
    .B(\gps_channel0.ca_nco.accumulator[3] ),
    .Y(_0578_));
 sky130_fd_sc_hd__or2_1 _1278_ (.A(\gps_channel0.ca_nco.step[2] ),
    .B(\gps_channel0.ca_nco.accumulator[2] ),
    .X(_0579_));
 sky130_fd_sc_hd__xor2_1 _1279_ (.A(\gps_channel0.ca_nco.step[1] ),
    .B(\gps_channel0.ca_nco.accumulator[1] ),
    .X(_0580_));
 sky130_fd_sc_hd__and2_1 _1280_ (.A(\gps_channel0.ca_nco.step[1] ),
    .B(\gps_channel0.ca_nco.accumulator[1] ),
    .X(_0581_));
 sky130_fd_sc_hd__a31o_1 _1281_ (.A1(\gps_channel0.ca_nco.step[0] ),
    .A2(\gps_channel0.ca_nco.accumulator[0] ),
    .A3(_0580_),
    .B1(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__nand2_1 _1282_ (.A(\gps_channel0.ca_nco.step[2] ),
    .B(\gps_channel0.ca_nco.accumulator[2] ),
    .Y(_0583_));
 sky130_fd_sc_hd__a21boi_2 _1283_ (.A1(_0579_),
    .A2(_0582_),
    .B1_N(_0583_),
    .Y(_0584_));
 sky130_fd_sc_hd__xor2_1 _1284_ (.A(\gps_channel0.ca_nco.step[4] ),
    .B(\gps_channel0.ca_nco.accumulator[4] ),
    .X(_0585_));
 sky130_fd_sc_hd__inv_2 _1285_ (.A(_0585_),
    .Y(_0586_));
 sky130_fd_sc_hd__nor2_1 _1286_ (.A(\gps_channel0.ca_nco.step[3] ),
    .B(\gps_channel0.ca_nco.accumulator[3] ),
    .Y(_0587_));
 sky130_fd_sc_hd__or2_1 _1287_ (.A(\gps_channel0.ca_nco.step[5] ),
    .B(\gps_channel0.ca_nco.accumulator[5] ),
    .X(_0588_));
 sky130_fd_sc_hd__nand2_1 _1288_ (.A(\gps_channel0.ca_nco.step[5] ),
    .B(\gps_channel0.ca_nco.accumulator[5] ),
    .Y(_0589_));
 sky130_fd_sc_hd__nand2_1 _1289_ (.A(_0588_),
    .B(_0589_),
    .Y(_0590_));
 sky130_fd_sc_hd__a2111o_1 _1290_ (.A1(_0578_),
    .A2(_0584_),
    .B1(_0586_),
    .C1(_0587_),
    .D1(_0590_),
    .X(_0591_));
 sky130_fd_sc_hd__nor2_1 _1291_ (.A(\gps_channel0.ca_nco.step[7] ),
    .B(\gps_channel0.ca_nco.accumulator[7] ),
    .Y(_0592_));
 sky130_fd_sc_hd__nand2_1 _1292_ (.A(\gps_channel0.ca_nco.step[6] ),
    .B(\gps_channel0.ca_nco.accumulator[6] ),
    .Y(_0593_));
 sky130_fd_sc_hd__a22o_1 _1293_ (.A1(\gps_channel0.ca_nco.step[4] ),
    .A2(\gps_channel0.ca_nco.accumulator[4] ),
    .B1(\gps_channel0.ca_nco.accumulator[5] ),
    .B2(\gps_channel0.ca_nco.step[5] ),
    .X(_0594_));
 sky130_fd_sc_hd__nand2_1 _1294_ (.A(_0588_),
    .B(_0594_),
    .Y(_0595_));
 sky130_fd_sc_hd__nand2_1 _1295_ (.A(\gps_channel0.ca_nco.step[7] ),
    .B(\gps_channel0.ca_nco.accumulator[7] ),
    .Y(_0596_));
 sky130_fd_sc_hd__o211a_1 _1296_ (.A1(_0592_),
    .A2(_0593_),
    .B1(_0595_),
    .C1(_0596_),
    .X(_0597_));
 sky130_fd_sc_hd__nor2_1 _1297_ (.A(\gps_channel0.ca_nco.step[6] ),
    .B(\gps_channel0.ca_nco.accumulator[6] ),
    .Y(_0598_));
 sky130_fd_sc_hd__a21o_1 _1298_ (.A1(_0596_),
    .A2(_0598_),
    .B1(_0592_),
    .X(_0599_));
 sky130_fd_sc_hd__or2b_1 _1299_ (.A(_0575_),
    .B_N(_0573_),
    .X(_0600_));
 sky130_fd_sc_hd__or2_1 _1300_ (.A(\gps_channel0.ca_nco.step[8] ),
    .B(\gps_channel0.ca_nco.accumulator[8] ),
    .X(_0601_));
 sky130_fd_sc_hd__nand2_1 _1301_ (.A(_0574_),
    .B(_0601_),
    .Y(_0602_));
 sky130_fd_sc_hd__or2_1 _1302_ (.A(_0600_),
    .B(_0602_),
    .X(_0603_));
 sky130_fd_sc_hd__a2111o_1 _1303_ (.A1(_0591_),
    .A2(_0597_),
    .B1(_0599_),
    .C1(_0572_),
    .D1(_0603_),
    .X(_0604_));
 sky130_fd_sc_hd__nand2_1 _1304_ (.A(\gps_channel0.ca_nco.step[12] ),
    .B(\gps_channel0.ca_nco.accumulator[12] ),
    .Y(_0605_));
 sky130_fd_sc_hd__or2_1 _1305_ (.A(\gps_channel0.ca_nco.step[12] ),
    .B(\gps_channel0.ca_nco.accumulator[12] ),
    .X(_0606_));
 sky130_fd_sc_hd__nand2_1 _1306_ (.A(_0605_),
    .B(_0606_),
    .Y(_0607_));
 sky130_fd_sc_hd__a21oi_2 _1307_ (.A1(_0577_),
    .A2(_0604_),
    .B1(_0607_),
    .Y(_0608_));
 sky130_fd_sc_hd__nand2_1 _1308_ (.A(\gps_channel0.ca_nco.step[15] ),
    .B(\gps_channel0.ca_nco.accumulator[15] ),
    .Y(_0609_));
 sky130_fd_sc_hd__or2_1 _1309_ (.A(\gps_channel0.ca_nco.step[15] ),
    .B(\gps_channel0.ca_nco.accumulator[15] ),
    .X(_0610_));
 sky130_fd_sc_hd__nand2_1 _1310_ (.A(_0609_),
    .B(_0610_),
    .Y(_0611_));
 sky130_fd_sc_hd__nand2_1 _1311_ (.A(\gps_channel0.ca_nco.step[14] ),
    .B(\gps_channel0.ca_nco.accumulator[14] ),
    .Y(_0612_));
 sky130_fd_sc_hd__or2_1 _1312_ (.A(\gps_channel0.ca_nco.step[14] ),
    .B(\gps_channel0.ca_nco.accumulator[14] ),
    .X(_0613_));
 sky130_fd_sc_hd__nand2_1 _1313_ (.A(_0612_),
    .B(_0613_),
    .Y(_0614_));
 sky130_fd_sc_hd__nor2_1 _1314_ (.A(_0611_),
    .B(_0614_),
    .Y(_0615_));
 sky130_fd_sc_hd__nor2_1 _1315_ (.A(\gps_channel0.ca_nco.step[13] ),
    .B(\gps_channel0.ca_nco.accumulator[13] ),
    .Y(_0616_));
 sky130_fd_sc_hd__nand2_1 _1316_ (.A(\gps_channel0.ca_nco.step[13] ),
    .B(\gps_channel0.ca_nco.accumulator[13] ),
    .Y(_0617_));
 sky130_fd_sc_hd__and2b_1 _1317_ (.A_N(_0616_),
    .B(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__a21oi_1 _1318_ (.A1(_0605_),
    .A2(_0617_),
    .B1(_0616_),
    .Y(_0619_));
 sky130_fd_sc_hd__and3_1 _1319_ (.A(\gps_channel0.ca_nco.step[14] ),
    .B(\gps_channel0.ca_nco.accumulator[14] ),
    .C(_0610_),
    .X(_0620_));
 sky130_fd_sc_hd__a221o_1 _1320_ (.A1(\gps_channel0.ca_nco.step[15] ),
    .A2(\gps_channel0.ca_nco.accumulator[15] ),
    .B1(_0615_),
    .B2(_0619_),
    .C1(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__a31o_2 _1321_ (.A1(_0608_),
    .A2(_0615_),
    .A3(_0618_),
    .B1(_0621_),
    .X(_0622_));
 sky130_fd_sc_hd__clkbuf_4 _1322_ (.A(\gps_channel0.ca_nco.step[16] ),
    .X(_0623_));
 sky130_fd_sc_hd__nor2_1 _1323_ (.A(_0623_),
    .B(\gps_channel0.ca_nco.accumulator[16] ),
    .Y(_0624_));
 sky130_fd_sc_hd__and2_1 _1324_ (.A(_0623_),
    .B(\gps_channel0.ca_nco.accumulator[16] ),
    .X(_0625_));
 sky130_fd_sc_hd__nor2_1 _1325_ (.A(_0624_),
    .B(_0625_),
    .Y(_0626_));
 sky130_fd_sc_hd__and2_1 _1326_ (.A(_0622_),
    .B(_0626_),
    .X(_0627_));
 sky130_fd_sc_hd__or2_1 _1327_ (.A(\gps_channel0.ca_nco.phase_sync ),
    .B(net3),
    .X(_0628_));
 sky130_fd_sc_hd__buf_4 _1328_ (.A(_0628_),
    .X(_0629_));
 sky130_fd_sc_hd__nor2_1 _1329_ (.A(net19),
    .B(_0628_),
    .Y(_0630_));
 sky130_fd_sc_hd__nor2_4 _1330_ (.A(_0629_),
    .B(_0630_),
    .Y(_0631_));
 sky130_fd_sc_hd__o21ai_1 _1331_ (.A1(_0622_),
    .A2(_0626_),
    .B1(_0631_),
    .Y(_0632_));
 sky130_fd_sc_hd__buf_4 _1332_ (.A(_0630_),
    .X(_0633_));
 sky130_fd_sc_hd__clkbuf_4 _1333_ (.A(_0633_),
    .X(_0634_));
 sky130_fd_sc_hd__a2bb2o_1 _1334_ (.A1_N(_0627_),
    .A2_N(_0632_),
    .B1(\gps_channel0.ca_nco.accumulator[16] ),
    .B2(_0634_),
    .X(_0046_));
 sky130_fd_sc_hd__clkbuf_4 _1335_ (.A(_0631_),
    .X(_0635_));
 sky130_fd_sc_hd__xor2_1 _1336_ (.A(_0623_),
    .B(\gps_channel0.ca_nco.accumulator[17] ),
    .X(_0636_));
 sky130_fd_sc_hd__o21ai_1 _1337_ (.A1(_0625_),
    .A2(_0627_),
    .B1(_0636_),
    .Y(_0637_));
 sky130_fd_sc_hd__or3_1 _1338_ (.A(_0625_),
    .B(_0627_),
    .C(_0636_),
    .X(_0638_));
 sky130_fd_sc_hd__a32o_1 _1339_ (.A1(_0635_),
    .A2(_0637_),
    .A3(_0638_),
    .B1(_0634_),
    .B2(\gps_channel0.ca_nco.accumulator[17] ),
    .X(_0047_));
 sky130_fd_sc_hd__nand2_1 _1340_ (.A(_0627_),
    .B(_0636_),
    .Y(_0639_));
 sky130_fd_sc_hd__buf_2 _1341_ (.A(_0623_),
    .X(_0640_));
 sky130_fd_sc_hd__o21ai_1 _1342_ (.A1(\gps_channel0.ca_nco.accumulator[16] ),
    .A2(\gps_channel0.ca_nco.accumulator[17] ),
    .B1(_0640_),
    .Y(_0641_));
 sky130_fd_sc_hd__nand2_1 _1343_ (.A(_0623_),
    .B(\gps_channel0.ca_nco.accumulator[18] ),
    .Y(_0642_));
 sky130_fd_sc_hd__or2_1 _1344_ (.A(_0623_),
    .B(\gps_channel0.ca_nco.accumulator[18] ),
    .X(_0643_));
 sky130_fd_sc_hd__nand2_1 _1345_ (.A(_0642_),
    .B(_0643_),
    .Y(_0644_));
 sky130_fd_sc_hd__a21o_1 _1346_ (.A1(_0639_),
    .A2(_0641_),
    .B1(_0644_),
    .X(_0645_));
 sky130_fd_sc_hd__nand3_1 _1347_ (.A(_0644_),
    .B(_0639_),
    .C(_0641_),
    .Y(_0646_));
 sky130_fd_sc_hd__clkbuf_4 _1348_ (.A(_0630_),
    .X(_0647_));
 sky130_fd_sc_hd__a32o_1 _1349_ (.A1(_0635_),
    .A2(_0645_),
    .A3(_0646_),
    .B1(_0647_),
    .B2(\gps_channel0.ca_nco.accumulator[18] ),
    .X(_0048_));
 sky130_fd_sc_hd__xnor2_1 _1350_ (.A(_0623_),
    .B(\gps_channel0.ca_nco.accumulator[19] ),
    .Y(_0648_));
 sky130_fd_sc_hd__a21oi_1 _1351_ (.A1(_0642_),
    .A2(_0645_),
    .B1(_0648_),
    .Y(_0649_));
 sky130_fd_sc_hd__clkinv_2 _1352_ (.A(_0631_),
    .Y(_0650_));
 sky130_fd_sc_hd__a31o_1 _1353_ (.A1(_0642_),
    .A2(_0645_),
    .A3(_0648_),
    .B1(_0650_),
    .X(_0651_));
 sky130_fd_sc_hd__a2bb2o_1 _1354_ (.A1_N(_0649_),
    .A2_N(_0651_),
    .B1(\gps_channel0.ca_nco.accumulator[19] ),
    .B2(_0634_),
    .X(_0049_));
 sky130_fd_sc_hd__or2_1 _1355_ (.A(\gps_channel0.ca_nco.step[16] ),
    .B(\gps_channel0.ca_nco.accumulator[20] ),
    .X(_0652_));
 sky130_fd_sc_hd__nand2_1 _1356_ (.A(\gps_channel0.ca_nco.step[16] ),
    .B(\gps_channel0.ca_nco.accumulator[20] ),
    .Y(_0653_));
 sky130_fd_sc_hd__nand2_1 _1357_ (.A(_0652_),
    .B(_0653_),
    .Y(_0654_));
 sky130_fd_sc_hd__nor2_1 _1358_ (.A(_0644_),
    .B(_0648_),
    .Y(_0655_));
 sky130_fd_sc_hd__and3_1 _1359_ (.A(_0626_),
    .B(_0636_),
    .C(_0655_),
    .X(_0656_));
 sky130_fd_sc_hd__o41a_1 _1360_ (.A1(\gps_channel0.ca_nco.accumulator[16] ),
    .A2(\gps_channel0.ca_nco.accumulator[17] ),
    .A3(\gps_channel0.ca_nco.accumulator[18] ),
    .A4(\gps_channel0.ca_nco.accumulator[19] ),
    .B1(_0623_),
    .X(_0657_));
 sky130_fd_sc_hd__a21oi_2 _1361_ (.A1(_0622_),
    .A2(_0656_),
    .B1(_0657_),
    .Y(_0658_));
 sky130_fd_sc_hd__or2_1 _1362_ (.A(_0654_),
    .B(_0658_),
    .X(_0659_));
 sky130_fd_sc_hd__nand2_1 _1363_ (.A(_0654_),
    .B(_0658_),
    .Y(_0660_));
 sky130_fd_sc_hd__a32o_1 _1364_ (.A1(_0635_),
    .A2(_0659_),
    .A3(_0660_),
    .B1(_0647_),
    .B2(\gps_channel0.ca_nco.accumulator[20] ),
    .X(_0050_));
 sky130_fd_sc_hd__xnor2_1 _1365_ (.A(\gps_channel0.ca_nco.step[16] ),
    .B(\gps_channel0.ca_nco.accumulator[21] ),
    .Y(_0661_));
 sky130_fd_sc_hd__o21a_1 _1366_ (.A1(_0654_),
    .A2(_0658_),
    .B1(_0653_),
    .X(_0662_));
 sky130_fd_sc_hd__xor2_1 _1367_ (.A(_0661_),
    .B(_0662_),
    .X(_0663_));
 sky130_fd_sc_hd__a22o_1 _1368_ (.A1(\gps_channel0.ca_nco.accumulator[21] ),
    .A2(_0634_),
    .B1(_0635_),
    .B2(_0663_),
    .X(_0051_));
 sky130_fd_sc_hd__nand2_1 _1369_ (.A(\gps_channel0.ca_nco.step[16] ),
    .B(\gps_channel0.ca_nco.accumulator[22] ),
    .Y(_0664_));
 sky130_fd_sc_hd__or2_1 _1370_ (.A(\gps_channel0.ca_nco.step[16] ),
    .B(\gps_channel0.ca_nco.accumulator[22] ),
    .X(_0665_));
 sky130_fd_sc_hd__nand2_1 _1371_ (.A(_0664_),
    .B(_0665_),
    .Y(_0666_));
 sky130_fd_sc_hd__or3_1 _1372_ (.A(_0654_),
    .B(_0658_),
    .C(_0661_),
    .X(_0667_));
 sky130_fd_sc_hd__o21ai_1 _1373_ (.A1(\gps_channel0.ca_nco.accumulator[20] ),
    .A2(\gps_channel0.ca_nco.accumulator[21] ),
    .B1(_0640_),
    .Y(_0668_));
 sky130_fd_sc_hd__and3_1 _1374_ (.A(_0666_),
    .B(_0667_),
    .C(_0668_),
    .X(_0669_));
 sky130_fd_sc_hd__a21o_1 _1375_ (.A1(_0667_),
    .A2(_0668_),
    .B1(_0666_),
    .X(_0670_));
 sky130_fd_sc_hd__nand2_1 _1376_ (.A(_0631_),
    .B(_0670_),
    .Y(_0671_));
 sky130_fd_sc_hd__a2bb2o_1 _1377_ (.A1_N(_0669_),
    .A2_N(_0671_),
    .B1(\gps_channel0.ca_nco.accumulator[22] ),
    .B2(_0634_),
    .X(_0052_));
 sky130_fd_sc_hd__xor2_1 _1378_ (.A(\gps_channel0.ca_nco.step[16] ),
    .B(\gps_channel0.ca_nco.accumulator[23] ),
    .X(_0672_));
 sky130_fd_sc_hd__inv_2 _1379_ (.A(_0672_),
    .Y(_0673_));
 sky130_fd_sc_hd__nand3_1 _1380_ (.A(_0664_),
    .B(_0670_),
    .C(_0673_),
    .Y(_0674_));
 sky130_fd_sc_hd__a21o_1 _1381_ (.A1(_0664_),
    .A2(_0670_),
    .B1(_0673_),
    .X(_0675_));
 sky130_fd_sc_hd__a32o_1 _1382_ (.A1(_0631_),
    .A2(_0674_),
    .A3(_0675_),
    .B1(_0647_),
    .B2(\gps_channel0.ca_nco.accumulator[23] ),
    .X(_0053_));
 sky130_fd_sc_hd__inv_2 _1383_ (.A(_0657_),
    .Y(_0676_));
 sky130_fd_sc_hd__or4_1 _1384_ (.A(_0654_),
    .B(_0661_),
    .C(_0666_),
    .D(_0673_),
    .X(_0677_));
 sky130_fd_sc_hd__inv_2 _1385_ (.A(_0677_),
    .Y(_0678_));
 sky130_fd_sc_hd__o41a_1 _1386_ (.A1(\gps_channel0.ca_nco.accumulator[20] ),
    .A2(\gps_channel0.ca_nco.accumulator[21] ),
    .A3(\gps_channel0.ca_nco.accumulator[22] ),
    .A4(\gps_channel0.ca_nco.accumulator[23] ),
    .B1(_0640_),
    .X(_0679_));
 sky130_fd_sc_hd__a31oi_1 _1387_ (.A1(_0622_),
    .A2(_0656_),
    .A3(_0678_),
    .B1(_0679_),
    .Y(_0680_));
 sky130_fd_sc_hd__and2_1 _1388_ (.A(_0676_),
    .B(_0680_),
    .X(_0681_));
 sky130_fd_sc_hd__xnor2_1 _1389_ (.A(_0623_),
    .B(\gps_channel0.ca_nco.accumulator[24] ),
    .Y(_0682_));
 sky130_fd_sc_hd__xor2_1 _1390_ (.A(_0681_),
    .B(_0682_),
    .X(_0683_));
 sky130_fd_sc_hd__a22o_1 _1391_ (.A1(\gps_channel0.ca_nco.accumulator[24] ),
    .A2(_0634_),
    .B1(_0635_),
    .B2(_0683_),
    .X(_0054_));
 sky130_fd_sc_hd__xor2_1 _1392_ (.A(_0623_),
    .B(\gps_channel0.ca_nco.accumulator[25] ),
    .X(_0684_));
 sky130_fd_sc_hd__a2bb2o_1 _1393_ (.A1_N(_0681_),
    .A2_N(_0682_),
    .B1(_0640_),
    .B2(\gps_channel0.ca_nco.accumulator[24] ),
    .X(_0685_));
 sky130_fd_sc_hd__nand2_1 _1394_ (.A(_0684_),
    .B(_0685_),
    .Y(_0686_));
 sky130_fd_sc_hd__o21a_1 _1395_ (.A1(_0684_),
    .A2(_0685_),
    .B1(_0631_),
    .X(_0687_));
 sky130_fd_sc_hd__a22o_1 _1396_ (.A1(\gps_channel0.ca_nco.accumulator[25] ),
    .A2(_0634_),
    .B1(_0686_),
    .B2(_0687_),
    .X(_0055_));
 sky130_fd_sc_hd__or2b_1 _1397_ (.A(_0682_),
    .B_N(_0684_),
    .X(_0688_));
 sky130_fd_sc_hd__a21o_1 _1398_ (.A1(_0676_),
    .A2(_0680_),
    .B1(_0688_),
    .X(_0689_));
 sky130_fd_sc_hd__o21ai_2 _1399_ (.A1(\gps_channel0.ca_nco.accumulator[24] ),
    .A2(\gps_channel0.ca_nco.accumulator[25] ),
    .B1(_0640_),
    .Y(_0690_));
 sky130_fd_sc_hd__or2_1 _1400_ (.A(_0640_),
    .B(\gps_channel0.ca_nco.accumulator[26] ),
    .X(_0691_));
 sky130_fd_sc_hd__nand2_1 _1401_ (.A(_0640_),
    .B(\gps_channel0.ca_nco.accumulator[26] ),
    .Y(_0692_));
 sky130_fd_sc_hd__nand2_1 _1402_ (.A(_0691_),
    .B(_0692_),
    .Y(_0693_));
 sky130_fd_sc_hd__a21o_1 _1403_ (.A1(_0689_),
    .A2(_0690_),
    .B1(_0693_),
    .X(_0694_));
 sky130_fd_sc_hd__a31oi_1 _1404_ (.A1(_0693_),
    .A2(_0689_),
    .A3(_0690_),
    .B1(_0650_),
    .Y(_0695_));
 sky130_fd_sc_hd__a22o_1 _1405_ (.A1(\gps_channel0.ca_nco.accumulator[26] ),
    .A2(_0634_),
    .B1(_0694_),
    .B2(_0695_),
    .X(_0056_));
 sky130_fd_sc_hd__xnor2_1 _1406_ (.A(_0640_),
    .B(\gps_channel0.ca_nco.accumulator[27] ),
    .Y(_0696_));
 sky130_fd_sc_hd__a21oi_1 _1407_ (.A1(_0692_),
    .A2(_0694_),
    .B1(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__a31o_1 _1408_ (.A1(_0692_),
    .A2(_0694_),
    .A3(_0696_),
    .B1(_0650_),
    .X(_0698_));
 sky130_fd_sc_hd__a2bb2o_1 _1409_ (.A1_N(_0697_),
    .A2_N(_0698_),
    .B1(\gps_channel0.ca_nco.accumulator[27] ),
    .B2(_0634_),
    .X(_0057_));
 sky130_fd_sc_hd__or2_1 _1410_ (.A(_0693_),
    .B(_0696_),
    .X(_0699_));
 sky130_fd_sc_hd__o21ai_1 _1411_ (.A1(\gps_channel0.ca_nco.accumulator[26] ),
    .A2(\gps_channel0.ca_nco.accumulator[27] ),
    .B1(_0640_),
    .Y(_0700_));
 sky130_fd_sc_hd__o211ai_4 _1412_ (.A1(_0689_),
    .A2(_0699_),
    .B1(_0700_),
    .C1(_0690_),
    .Y(_0701_));
 sky130_fd_sc_hd__a31oi_1 _1413_ (.A1(net19),
    .A2(\gps_channel0.ca_nco.accumulator[28] ),
    .A3(_0701_),
    .B1(_0629_),
    .Y(_0702_));
 sky130_fd_sc_hd__a21o_1 _1414_ (.A1(_0631_),
    .A2(_0701_),
    .B1(\gps_channel0.ca_nco.accumulator[28] ),
    .X(_0703_));
 sky130_fd_sc_hd__and2_1 _1415_ (.A(_0702_),
    .B(_0703_),
    .X(_0704_));
 sky130_fd_sc_hd__clkbuf_1 _1416_ (.A(_0704_),
    .X(_0058_));
 sky130_fd_sc_hd__and3_1 _1417_ (.A(\gps_channel0.ca_nco.accumulator[28] ),
    .B(_0631_),
    .C(_0701_),
    .X(_0705_));
 sky130_fd_sc_hd__mux2_1 _1418_ (.A0(_0705_),
    .A1(_0702_),
    .S(\gps_channel0.ca_nco.accumulator[29] ),
    .X(_0706_));
 sky130_fd_sc_hd__clkbuf_1 _1419_ (.A(_0706_),
    .X(_0059_));
 sky130_fd_sc_hd__and2_1 _1420_ (.A(\gps_channel0.ca_nco.accumulator[28] ),
    .B(\gps_channel0.ca_nco.accumulator[29] ),
    .X(_0707_));
 sky130_fd_sc_hd__a21oi_1 _1421_ (.A1(_0701_),
    .A2(_0707_),
    .B1(\gps_channel0.ca_nco.accumulator[30] ),
    .Y(_0708_));
 sky130_fd_sc_hd__a31o_1 _1422_ (.A1(\gps_channel0.ca_nco.accumulator[30] ),
    .A2(_0701_),
    .A3(_0707_),
    .B1(_0650_),
    .X(_0709_));
 sky130_fd_sc_hd__a2bb2o_1 _1423_ (.A1_N(_0708_),
    .A2_N(_0709_),
    .B1(\gps_channel0.ca_nco.accumulator[30] ),
    .B2(_0634_),
    .X(_0060_));
 sky130_fd_sc_hd__inv_2 _1424_ (.A(\gps_channel0.ca_nco.accumulator[31] ),
    .Y(_0010_));
 sky130_fd_sc_hd__nor2_1 _1425_ (.A(_0010_),
    .B(_0647_),
    .Y(_0710_));
 sky130_fd_sc_hd__and4_1 _1426_ (.A(\gps_channel0.ca_nco.accumulator[30] ),
    .B(_0631_),
    .C(_0701_),
    .D(_0707_),
    .X(_0711_));
 sky130_fd_sc_hd__buf_4 _1427_ (.A(\gps_channel0.ca_nco.accumulator[31] ),
    .X(_0712_));
 sky130_fd_sc_hd__o2bb2a_1 _1428_ (.A1_N(_0709_),
    .A2_N(_0710_),
    .B1(_0711_),
    .B2(_0712_),
    .X(_0061_));
 sky130_fd_sc_hd__nand2_1 _1429_ (.A(\gps_channel0.ca_nco.step[0] ),
    .B(net19),
    .Y(_0713_));
 sky130_fd_sc_hd__xnor2_1 _1430_ (.A(\gps_channel0.ca_nco.accumulator[0] ),
    .B(_0713_),
    .Y(_0714_));
 sky130_fd_sc_hd__nor2_8 _1431_ (.A(\gps_channel0.ca_nco.phase_sync ),
    .B(net3),
    .Y(_0715_));
 sky130_fd_sc_hd__mux2_1 _1432_ (.A0(\gps_channel0.ca_nco.phase_in[0] ),
    .A1(_0714_),
    .S(_0715_),
    .X(_0716_));
 sky130_fd_sc_hd__clkbuf_1 _1433_ (.A(_0716_),
    .X(_0062_));
 sky130_fd_sc_hd__a21oi_1 _1434_ (.A1(\gps_channel0.ca_nco.step[0] ),
    .A2(\gps_channel0.ca_nco.accumulator[0] ),
    .B1(_0580_),
    .Y(_0717_));
 sky130_fd_sc_hd__a311oi_1 _1435_ (.A1(\gps_channel0.ca_nco.step[0] ),
    .A2(\gps_channel0.ca_nco.accumulator[0] ),
    .A3(_0580_),
    .B1(_0650_),
    .C1(_0717_),
    .Y(_0718_));
 sky130_fd_sc_hd__a221o_1 _1436_ (.A1(\gps_channel0.ca_nco.phase_in[1] ),
    .A2(_0629_),
    .B1(_0647_),
    .B2(\gps_channel0.ca_nco.accumulator[1] ),
    .C1(_0718_),
    .X(_0063_));
 sky130_fd_sc_hd__nand2_1 _1437_ (.A(_0583_),
    .B(_0579_),
    .Y(_0719_));
 sky130_fd_sc_hd__xnor2_1 _1438_ (.A(_0719_),
    .B(_0582_),
    .Y(_0720_));
 sky130_fd_sc_hd__mux2_1 _1439_ (.A0(\gps_channel0.ca_nco.phase_in[2] ),
    .A1(_0720_),
    .S(_0715_),
    .X(_0721_));
 sky130_fd_sc_hd__mux2_1 _1440_ (.A0(_0721_),
    .A1(\gps_channel0.ca_nco.accumulator[2] ),
    .S(_0633_),
    .X(_0722_));
 sky130_fd_sc_hd__clkbuf_1 _1441_ (.A(_0722_),
    .X(_0064_));
 sky130_fd_sc_hd__and2b_1 _1442_ (.A_N(_0587_),
    .B(_0578_),
    .X(_0723_));
 sky130_fd_sc_hd__xnor2_1 _1443_ (.A(_0584_),
    .B(_0723_),
    .Y(_0724_));
 sky130_fd_sc_hd__mux2_1 _1444_ (.A0(\gps_channel0.ca_nco.phase_in[3] ),
    .A1(_0724_),
    .S(_0715_),
    .X(_0725_));
 sky130_fd_sc_hd__mux2_1 _1445_ (.A0(_0725_),
    .A1(\gps_channel0.ca_nco.accumulator[3] ),
    .S(_0633_),
    .X(_0726_));
 sky130_fd_sc_hd__clkbuf_1 _1446_ (.A(_0726_),
    .X(_0065_));
 sky130_fd_sc_hd__a21oi_1 _1447_ (.A1(_0578_),
    .A2(_0584_),
    .B1(_0587_),
    .Y(_0727_));
 sky130_fd_sc_hd__nand2_1 _1448_ (.A(_0727_),
    .B(_0585_),
    .Y(_0728_));
 sky130_fd_sc_hd__or2_1 _1449_ (.A(_0727_),
    .B(_0585_),
    .X(_0729_));
 sky130_fd_sc_hd__a22o_1 _1450_ (.A1(\gps_channel0.ca_nco.phase_in[4] ),
    .A2(_0629_),
    .B1(_0647_),
    .B2(\gps_channel0.ca_nco.accumulator[4] ),
    .X(_0730_));
 sky130_fd_sc_hd__a31o_1 _1451_ (.A1(_0728_),
    .A2(_0635_),
    .A3(_0729_),
    .B1(_0730_),
    .X(_0066_));
 sky130_fd_sc_hd__a21bo_1 _1452_ (.A1(\gps_channel0.ca_nco.step[4] ),
    .A2(\gps_channel0.ca_nco.accumulator[4] ),
    .B1_N(_0728_),
    .X(_0731_));
 sky130_fd_sc_hd__xnor2_1 _1453_ (.A(_0590_),
    .B(_0731_),
    .Y(_0732_));
 sky130_fd_sc_hd__mux2_1 _1454_ (.A0(\gps_channel0.ca_nco.phase_in[5] ),
    .A1(_0732_),
    .S(_0715_),
    .X(_0733_));
 sky130_fd_sc_hd__mux2_1 _1455_ (.A0(_0733_),
    .A1(\gps_channel0.ca_nco.accumulator[5] ),
    .S(_0633_),
    .X(_0734_));
 sky130_fd_sc_hd__clkbuf_1 _1456_ (.A(_0734_),
    .X(_0067_));
 sky130_fd_sc_hd__and2_1 _1457_ (.A(\gps_channel0.ca_nco.step[6] ),
    .B(\gps_channel0.ca_nco.accumulator[6] ),
    .X(_0735_));
 sky130_fd_sc_hd__o211ai_1 _1458_ (.A1(_0735_),
    .A2(_0598_),
    .B1(_0591_),
    .C1(_0595_),
    .Y(_0736_));
 sky130_fd_sc_hd__a211o_1 _1459_ (.A1(_0591_),
    .A2(_0595_),
    .B1(_0735_),
    .C1(_0598_),
    .X(_0737_));
 sky130_fd_sc_hd__a22o_1 _1460_ (.A1(\gps_channel0.ca_nco.phase_in[6] ),
    .A2(_0629_),
    .B1(_0633_),
    .B2(\gps_channel0.ca_nco.accumulator[6] ),
    .X(_0738_));
 sky130_fd_sc_hd__a31o_1 _1461_ (.A1(_0635_),
    .A2(_0736_),
    .A3(_0737_),
    .B1(_0738_),
    .X(_0068_));
 sky130_fd_sc_hd__and2_1 _1462_ (.A(\gps_channel0.ca_nco.step[7] ),
    .B(\gps_channel0.ca_nco.accumulator[7] ),
    .X(_0739_));
 sky130_fd_sc_hd__nor2_1 _1463_ (.A(_0739_),
    .B(_0592_),
    .Y(_0740_));
 sky130_fd_sc_hd__a21oi_1 _1464_ (.A1(_0593_),
    .A2(_0737_),
    .B1(_0740_),
    .Y(_0741_));
 sky130_fd_sc_hd__a31o_1 _1465_ (.A1(_0593_),
    .A2(_0740_),
    .A3(_0737_),
    .B1(_0629_),
    .X(_0742_));
 sky130_fd_sc_hd__o22a_1 _1466_ (.A1(\gps_channel0.ca_nco.phase_in[7] ),
    .A2(_0715_),
    .B1(_0741_),
    .B2(_0742_),
    .X(_0743_));
 sky130_fd_sc_hd__mux2_1 _1467_ (.A0(_0743_),
    .A1(\gps_channel0.ca_nco.accumulator[7] ),
    .S(_0633_),
    .X(_0744_));
 sky130_fd_sc_hd__clkbuf_1 _1468_ (.A(_0744_),
    .X(_0069_));
 sky130_fd_sc_hd__a21o_1 _1469_ (.A1(_0591_),
    .A2(_0597_),
    .B1(_0599_),
    .X(_0745_));
 sky130_fd_sc_hd__or2_1 _1470_ (.A(_0745_),
    .B(_0602_),
    .X(_0746_));
 sky130_fd_sc_hd__nand2_1 _1471_ (.A(_0745_),
    .B(_0602_),
    .Y(_0747_));
 sky130_fd_sc_hd__and2_1 _1472_ (.A(_0746_),
    .B(_0747_),
    .X(_0748_));
 sky130_fd_sc_hd__a22o_1 _1473_ (.A1(\gps_channel0.ca_nco.phase_in[8] ),
    .A2(_0629_),
    .B1(_0647_),
    .B2(\gps_channel0.ca_nco.accumulator[8] ),
    .X(_0749_));
 sky130_fd_sc_hd__a21o_1 _1474_ (.A1(_0635_),
    .A2(_0748_),
    .B1(_0749_),
    .X(_0070_));
 sky130_fd_sc_hd__nand2_1 _1475_ (.A(_0574_),
    .B(_0746_),
    .Y(_0750_));
 sky130_fd_sc_hd__xnor2_1 _1476_ (.A(_0600_),
    .B(_0750_),
    .Y(_0182_));
 sky130_fd_sc_hd__mux2_1 _1477_ (.A0(\gps_channel0.ca_nco.phase_in[9] ),
    .A1(_0182_),
    .S(_0715_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _1478_ (.A0(_0183_),
    .A1(\gps_channel0.ca_nco.accumulator[9] ),
    .S(_0633_),
    .X(_0184_));
 sky130_fd_sc_hd__clkbuf_1 _1479_ (.A(_0184_),
    .X(_0071_));
 sky130_fd_sc_hd__o21a_1 _1480_ (.A1(_0600_),
    .A2(_0746_),
    .B1(_0576_),
    .X(_0185_));
 sky130_fd_sc_hd__xor2_1 _1481_ (.A(_0571_),
    .B(_0185_),
    .X(_0186_));
 sky130_fd_sc_hd__and3_1 _1482_ (.A(net19),
    .B(_0715_),
    .C(_0186_),
    .X(_0187_));
 sky130_fd_sc_hd__a221o_1 _1483_ (.A1(\gps_channel0.ca_nco.phase_in[10] ),
    .A2(_0629_),
    .B1(_0647_),
    .B2(\gps_channel0.ca_nco.accumulator[10] ),
    .C1(_0187_),
    .X(_0072_));
 sky130_fd_sc_hd__o21ai_1 _1484_ (.A1(_0571_),
    .A2(_0185_),
    .B1(_0567_),
    .Y(_0188_));
 sky130_fd_sc_hd__xnor2_1 _1485_ (.A(_0569_),
    .B(_0188_),
    .Y(_0189_));
 sky130_fd_sc_hd__a22o_1 _1486_ (.A1(\gps_channel0.ca_nco.phase_in[11] ),
    .A2(_0629_),
    .B1(_0647_),
    .B2(\gps_channel0.ca_nco.accumulator[11] ),
    .X(_0190_));
 sky130_fd_sc_hd__a21o_1 _1487_ (.A1(_0635_),
    .A2(_0189_),
    .B1(_0190_),
    .X(_0073_));
 sky130_fd_sc_hd__and3_1 _1488_ (.A(_0577_),
    .B(_0604_),
    .C(_0607_),
    .X(_0191_));
 sky130_fd_sc_hd__nor2_1 _1489_ (.A(_0608_),
    .B(_0191_),
    .Y(_0192_));
 sky130_fd_sc_hd__a22o_1 _1490_ (.A1(\gps_channel0.ca_nco.phase_in[12] ),
    .A2(_0629_),
    .B1(_0647_),
    .B2(\gps_channel0.ca_nco.accumulator[12] ),
    .X(_0193_));
 sky130_fd_sc_hd__a21o_1 _1491_ (.A1(_0635_),
    .A2(_0192_),
    .B1(_0193_),
    .X(_0074_));
 sky130_fd_sc_hd__a21oi_1 _1492_ (.A1(\gps_channel0.ca_nco.step[12] ),
    .A2(\gps_channel0.ca_nco.accumulator[12] ),
    .B1(_0608_),
    .Y(_0194_));
 sky130_fd_sc_hd__xnor2_1 _1493_ (.A(_0618_),
    .B(_0194_),
    .Y(_0195_));
 sky130_fd_sc_hd__mux2_1 _1494_ (.A0(\gps_channel0.ca_nco.phase_in[13] ),
    .A1(_0195_),
    .S(_0715_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _1495_ (.A0(_0196_),
    .A1(\gps_channel0.ca_nco.accumulator[13] ),
    .S(_0633_),
    .X(_0197_));
 sky130_fd_sc_hd__clkbuf_1 _1496_ (.A(_0197_),
    .X(_0075_));
 sky130_fd_sc_hd__a21oi_1 _1497_ (.A1(_0608_),
    .A2(_0618_),
    .B1(_0619_),
    .Y(_0198_));
 sky130_fd_sc_hd__xor2_1 _1498_ (.A(_0614_),
    .B(_0198_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _1499_ (.A0(\gps_channel0.ca_nco.phase_in[14] ),
    .A1(_0199_),
    .S(_0715_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _1500_ (.A0(_0200_),
    .A1(\gps_channel0.ca_nco.accumulator[14] ),
    .S(_0633_),
    .X(_0201_));
 sky130_fd_sc_hd__clkbuf_1 _1501_ (.A(_0201_),
    .X(_0076_));
 sky130_fd_sc_hd__o21ai_1 _1502_ (.A1(_0614_),
    .A2(_0198_),
    .B1(_0612_),
    .Y(_0202_));
 sky130_fd_sc_hd__xnor2_1 _1503_ (.A(_0611_),
    .B(_0202_),
    .Y(_0203_));
 sky130_fd_sc_hd__mux2_1 _1504_ (.A0(\gps_channel0.ca_nco.phase_in[15] ),
    .A1(_0203_),
    .S(_0715_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _1505_ (.A0(_0204_),
    .A1(\gps_channel0.ca_nco.accumulator[15] ),
    .S(_0633_),
    .X(_0205_));
 sky130_fd_sc_hd__clkbuf_1 _1506_ (.A(_0205_),
    .X(_0077_));
 sky130_fd_sc_hd__clkinv_2 _1507_ (.A(net24),
    .Y(_0206_));
 sky130_fd_sc_hd__or2_1 _1508_ (.A(net25),
    .B(net23),
    .X(_0207_));
 sky130_fd_sc_hd__or2_1 _1509_ (.A(_0206_),
    .B(_0207_),
    .X(_0208_));
 sky130_fd_sc_hd__clkbuf_2 _1510_ (.A(_0208_),
    .X(_0209_));
 sky130_fd_sc_hd__buf_2 _1511_ (.A(_0209_),
    .X(_0210_));
 sky130_fd_sc_hd__nor2_2 _1512_ (.A(_0206_),
    .B(_0207_),
    .Y(_0211_));
 sky130_fd_sc_hd__buf_2 _1513_ (.A(_0211_),
    .X(_0212_));
 sky130_fd_sc_hd__buf_2 _1514_ (.A(net3),
    .X(_0213_));
 sky130_fd_sc_hd__o21ba_1 _1515_ (.A1(\gps_channel0.lo_nco.phase_in[0] ),
    .A2(_0212_),
    .B1_N(_0213_),
    .X(_0214_));
 sky130_fd_sc_hd__o21a_1 _1516_ (.A1(net4),
    .A2(_0210_),
    .B1(_0214_),
    .X(_0078_));
 sky130_fd_sc_hd__o21ba_1 _1517_ (.A1(\gps_channel0.lo_nco.phase_in[1] ),
    .A2(_0212_),
    .B1_N(_0213_),
    .X(_0215_));
 sky130_fd_sc_hd__o21a_1 _1518_ (.A1(net5),
    .A2(_0210_),
    .B1(_0215_),
    .X(_0079_));
 sky130_fd_sc_hd__o21ba_1 _1519_ (.A1(\gps_channel0.lo_nco.phase_in[2] ),
    .A2(_0212_),
    .B1_N(_0213_),
    .X(_0216_));
 sky130_fd_sc_hd__o21a_1 _1520_ (.A1(net6),
    .A2(_0210_),
    .B1(_0216_),
    .X(_0080_));
 sky130_fd_sc_hd__o21ba_1 _1521_ (.A1(\gps_channel0.lo_nco.phase_in[3] ),
    .A2(_0212_),
    .B1_N(_0213_),
    .X(_0217_));
 sky130_fd_sc_hd__o21a_1 _1522_ (.A1(net7),
    .A2(_0210_),
    .B1(_0217_),
    .X(_0081_));
 sky130_fd_sc_hd__o21ba_1 _1523_ (.A1(\gps_channel0.lo_nco.phase_in[4] ),
    .A2(_0212_),
    .B1_N(_0213_),
    .X(_0218_));
 sky130_fd_sc_hd__o21a_1 _1524_ (.A1(net9),
    .A2(_0210_),
    .B1(_0218_),
    .X(_0082_));
 sky130_fd_sc_hd__o21ba_1 _1525_ (.A1(\gps_channel0.lo_nco.phase_in[5] ),
    .A2(_0212_),
    .B1_N(_0213_),
    .X(_0219_));
 sky130_fd_sc_hd__o21a_1 _1526_ (.A1(net10),
    .A2(_0210_),
    .B1(_0219_),
    .X(_0083_));
 sky130_fd_sc_hd__buf_2 _1527_ (.A(net3),
    .X(_0220_));
 sky130_fd_sc_hd__clkbuf_2 _1528_ (.A(_0220_),
    .X(_0221_));
 sky130_fd_sc_hd__o21ba_1 _1529_ (.A1(\gps_channel0.lo_nco.phase_in[6] ),
    .A2(_0212_),
    .B1_N(_0221_),
    .X(_0222_));
 sky130_fd_sc_hd__o21a_1 _1530_ (.A1(net11),
    .A2(_0210_),
    .B1(_0222_),
    .X(_0084_));
 sky130_fd_sc_hd__o21ba_1 _1531_ (.A1(\gps_channel0.lo_nco.phase_in[7] ),
    .A2(_0212_),
    .B1_N(_0221_),
    .X(_0223_));
 sky130_fd_sc_hd__o21a_1 _1532_ (.A1(net12),
    .A2(_0210_),
    .B1(_0223_),
    .X(_0085_));
 sky130_fd_sc_hd__o21ba_1 _1533_ (.A1(\gps_channel0.lo_nco.phase_in[8] ),
    .A2(_0212_),
    .B1_N(_0221_),
    .X(_0224_));
 sky130_fd_sc_hd__o21a_1 _1534_ (.A1(net13),
    .A2(_0210_),
    .B1(_0224_),
    .X(_0086_));
 sky130_fd_sc_hd__o21ba_1 _1535_ (.A1(\gps_channel0.lo_nco.phase_in[9] ),
    .A2(_0211_),
    .B1_N(_0221_),
    .X(_0225_));
 sky130_fd_sc_hd__o21a_1 _1536_ (.A1(net14),
    .A2(_0210_),
    .B1(_0225_),
    .X(_0087_));
 sky130_fd_sc_hd__o21ba_1 _1537_ (.A1(\gps_channel0.lo_nco.phase_in[10] ),
    .A2(_0211_),
    .B1_N(_0221_),
    .X(_0226_));
 sky130_fd_sc_hd__o21a_1 _1538_ (.A1(net15),
    .A2(_0209_),
    .B1(_0226_),
    .X(_0088_));
 sky130_fd_sc_hd__o21ba_1 _1539_ (.A1(\gps_channel0.lo_nco.phase_in[11] ),
    .A2(_0211_),
    .B1_N(_0221_),
    .X(_0227_));
 sky130_fd_sc_hd__o21a_1 _1540_ (.A1(net16),
    .A2(_0209_),
    .B1(_0227_),
    .X(_0089_));
 sky130_fd_sc_hd__o21ba_1 _1541_ (.A1(\gps_channel0.lo_nco.phase_in[12] ),
    .A2(_0211_),
    .B1_N(_0221_),
    .X(_0228_));
 sky130_fd_sc_hd__o21a_1 _1542_ (.A1(net17),
    .A2(_0209_),
    .B1(_0228_),
    .X(_0090_));
 sky130_fd_sc_hd__o21ba_1 _1543_ (.A1(\gps_channel0.lo_nco.phase_in[13] ),
    .A2(_0211_),
    .B1_N(_0221_),
    .X(_0229_));
 sky130_fd_sc_hd__o21a_1 _1544_ (.A1(net18),
    .A2(_0209_),
    .B1(_0229_),
    .X(_0091_));
 sky130_fd_sc_hd__o21ba_1 _1545_ (.A1(\gps_channel0.lo_nco.phase_in[14] ),
    .A2(_0211_),
    .B1_N(_0221_),
    .X(_0230_));
 sky130_fd_sc_hd__o21a_1 _1546_ (.A1(net20),
    .A2(_0209_),
    .B1(_0230_),
    .X(_0092_));
 sky130_fd_sc_hd__o21ba_1 _1547_ (.A1(\gps_channel0.lo_nco.phase_in[15] ),
    .A2(_0211_),
    .B1_N(_0221_),
    .X(_0231_));
 sky130_fd_sc_hd__o21a_1 _1548_ (.A1(net21),
    .A2(_0209_),
    .B1(_0231_),
    .X(_0093_));
 sky130_fd_sc_hd__clkbuf_8 _1549_ (.A(\gps_channel0.ca_nco.accumulator[31] ),
    .X(_0232_));
 sky130_fd_sc_hd__clkinv_2 _1550_ (.A(_0232_),
    .Y(_0011_));
 sky130_fd_sc_hd__clkinv_2 _1551_ (.A(_0232_),
    .Y(_0012_));
 sky130_fd_sc_hd__clkinv_2 _1552_ (.A(_0232_),
    .Y(_0013_));
 sky130_fd_sc_hd__clkinv_2 _1553_ (.A(_0232_),
    .Y(_0014_));
 sky130_fd_sc_hd__clkinv_2 _1554_ (.A(_0232_),
    .Y(_0015_));
 sky130_fd_sc_hd__clkinv_2 _1555_ (.A(_0232_),
    .Y(_0016_));
 sky130_fd_sc_hd__clkinv_2 _1556_ (.A(_0232_),
    .Y(_0017_));
 sky130_fd_sc_hd__clkinv_2 _1557_ (.A(_0232_),
    .Y(_0018_));
 sky130_fd_sc_hd__clkinv_2 _1558_ (.A(_0232_),
    .Y(_0019_));
 sky130_fd_sc_hd__clkinv_2 _1559_ (.A(_0232_),
    .Y(_0020_));
 sky130_fd_sc_hd__clkinv_2 _1560_ (.A(_0712_),
    .Y(_0021_));
 sky130_fd_sc_hd__clkinv_2 _1561_ (.A(_0712_),
    .Y(_0022_));
 sky130_fd_sc_hd__clkinv_2 _1562_ (.A(_0712_),
    .Y(_0023_));
 sky130_fd_sc_hd__clkinv_2 _1563_ (.A(_0712_),
    .Y(_0024_));
 sky130_fd_sc_hd__clkinv_2 _1564_ (.A(_0712_),
    .Y(_0025_));
 sky130_fd_sc_hd__clkinv_2 _1565_ (.A(_0712_),
    .Y(_0026_));
 sky130_fd_sc_hd__clkinv_2 _1566_ (.A(_0712_),
    .Y(_0027_));
 sky130_fd_sc_hd__clkinv_2 _1567_ (.A(_0712_),
    .Y(_0028_));
 sky130_fd_sc_hd__clkinv_2 _1568_ (.A(_0712_),
    .Y(_0029_));
 sky130_fd_sc_hd__or3_1 _1569_ (.A(_0555_),
    .B(_0559_),
    .C(_0560_),
    .X(_0233_));
 sky130_fd_sc_hd__or3_1 _1570_ (.A(_0543_),
    .B(_0549_),
    .C(_0233_),
    .X(_0234_));
 sky130_fd_sc_hd__a21oi_1 _1571_ (.A1(_0535_),
    .A2(_0539_),
    .B1(_0234_),
    .Y(_0235_));
 sky130_fd_sc_hd__a211oi_1 _1572_ (.A1(_0541_),
    .A2(_0548_),
    .B1(_0233_),
    .C1(_0547_),
    .Y(_0236_));
 sky130_fd_sc_hd__nor2_1 _1573_ (.A(_0554_),
    .B(_0559_),
    .Y(_0237_));
 sky130_fd_sc_hd__or3_1 _1574_ (.A(_0560_),
    .B(_0236_),
    .C(_0237_),
    .X(_0238_));
 sky130_fd_sc_hd__or2_1 _1575_ (.A(_0235_),
    .B(_0238_),
    .X(_0239_));
 sky130_fd_sc_hd__clkbuf_4 _1576_ (.A(\gps_channel0.lo_nco.step[16] ),
    .X(_0240_));
 sky130_fd_sc_hd__xor2_1 _1577_ (.A(_0240_),
    .B(\gps_channel0.lo_nco.accumulator[16] ),
    .X(_0241_));
 sky130_fd_sc_hd__and2_1 _1578_ (.A(_0239_),
    .B(_0241_),
    .X(_0242_));
 sky130_fd_sc_hd__o21ai_1 _1579_ (.A1(_0239_),
    .A2(_0241_),
    .B1(_0501_),
    .Y(_0243_));
 sky130_fd_sc_hd__a2bb2o_1 _1580_ (.A1_N(_0242_),
    .A2_N(_0243_),
    .B1(\gps_channel0.lo_nco.accumulator[16] ),
    .B2(_0525_),
    .X(_0104_));
 sky130_fd_sc_hd__xor2_1 _1581_ (.A(_0240_),
    .B(\gps_channel0.lo_nco.accumulator[17] ),
    .X(_0244_));
 sky130_fd_sc_hd__buf_2 _1582_ (.A(_0240_),
    .X(_0245_));
 sky130_fd_sc_hd__a21oi_1 _1583_ (.A1(_0245_),
    .A2(\gps_channel0.lo_nco.accumulator[16] ),
    .B1(_0242_),
    .Y(_0246_));
 sky130_fd_sc_hd__xnor2_1 _1584_ (.A(_0244_),
    .B(_0246_),
    .Y(_0247_));
 sky130_fd_sc_hd__a22o_1 _1585_ (.A1(\gps_channel0.lo_nco.accumulator[17] ),
    .A2(_0525_),
    .B1(_0247_),
    .B2(_0501_),
    .X(_0105_));
 sky130_fd_sc_hd__o21ai_1 _1586_ (.A1(\gps_channel0.lo_nco.accumulator[16] ),
    .A2(\gps_channel0.lo_nco.accumulator[17] ),
    .B1(_0245_),
    .Y(_0248_));
 sky130_fd_sc_hd__nand2_1 _1587_ (.A(_0242_),
    .B(_0244_),
    .Y(_0249_));
 sky130_fd_sc_hd__nand2_1 _1588_ (.A(_0240_),
    .B(\gps_channel0.lo_nco.accumulator[18] ),
    .Y(_0250_));
 sky130_fd_sc_hd__or2_1 _1589_ (.A(_0240_),
    .B(\gps_channel0.lo_nco.accumulator[18] ),
    .X(_0251_));
 sky130_fd_sc_hd__nand2_1 _1590_ (.A(_0250_),
    .B(_0251_),
    .Y(_0252_));
 sky130_fd_sc_hd__a21o_1 _1591_ (.A1(_0248_),
    .A2(_0249_),
    .B1(_0252_),
    .X(_0253_));
 sky130_fd_sc_hd__nand3_1 _1592_ (.A(_0252_),
    .B(_0248_),
    .C(_0249_),
    .Y(_0254_));
 sky130_fd_sc_hd__a32o_1 _1593_ (.A1(_0501_),
    .A2(_0253_),
    .A3(_0254_),
    .B1(_0525_),
    .B2(\gps_channel0.lo_nco.accumulator[18] ),
    .X(_0106_));
 sky130_fd_sc_hd__xnor2_1 _1594_ (.A(_0240_),
    .B(\gps_channel0.lo_nco.accumulator[19] ),
    .Y(_0255_));
 sky130_fd_sc_hd__a21oi_1 _1595_ (.A1(_0250_),
    .A2(_0253_),
    .B1(_0255_),
    .Y(_0256_));
 sky130_fd_sc_hd__a31o_1 _1596_ (.A1(_0250_),
    .A2(_0253_),
    .A3(_0255_),
    .B1(_0454_),
    .X(_0257_));
 sky130_fd_sc_hd__a2bb2o_1 _1597_ (.A1_N(_0256_),
    .A2_N(_0257_),
    .B1(\gps_channel0.lo_nco.accumulator[19] ),
    .B2(_0525_),
    .X(_0107_));
 sky130_fd_sc_hd__o41a_1 _1598_ (.A1(\gps_channel0.lo_nco.accumulator[16] ),
    .A2(\gps_channel0.lo_nco.accumulator[17] ),
    .A3(\gps_channel0.lo_nco.accumulator[18] ),
    .A4(\gps_channel0.lo_nco.accumulator[19] ),
    .B1(_0245_),
    .X(_0258_));
 sky130_fd_sc_hd__nor2_1 _1599_ (.A(_0252_),
    .B(_0255_),
    .Y(_0259_));
 sky130_fd_sc_hd__and3_1 _1600_ (.A(_0241_),
    .B(_0244_),
    .C(_0259_),
    .X(_0260_));
 sky130_fd_sc_hd__o21a_1 _1601_ (.A1(_0235_),
    .A2(_0238_),
    .B1(_0260_),
    .X(_0261_));
 sky130_fd_sc_hd__xor2_1 _1602_ (.A(_0245_),
    .B(\gps_channel0.lo_nco.accumulator[20] ),
    .X(_0262_));
 sky130_fd_sc_hd__o21a_1 _1603_ (.A1(_0258_),
    .A2(_0261_),
    .B1(_0262_),
    .X(_0263_));
 sky130_fd_sc_hd__o31ai_1 _1604_ (.A1(_0262_),
    .A2(_0258_),
    .A3(_0261_),
    .B1(_0501_),
    .Y(_0264_));
 sky130_fd_sc_hd__a2bb2o_1 _1605_ (.A1_N(_0263_),
    .A2_N(_0264_),
    .B1(\gps_channel0.lo_nco.accumulator[20] ),
    .B2(_0525_),
    .X(_0108_));
 sky130_fd_sc_hd__xor2_1 _1606_ (.A(_0240_),
    .B(\gps_channel0.lo_nco.accumulator[21] ),
    .X(_0265_));
 sky130_fd_sc_hd__a21oi_1 _1607_ (.A1(_0245_),
    .A2(\gps_channel0.lo_nco.accumulator[20] ),
    .B1(_0263_),
    .Y(_0266_));
 sky130_fd_sc_hd__xnor2_1 _1608_ (.A(_0265_),
    .B(_0266_),
    .Y(_0267_));
 sky130_fd_sc_hd__a22o_1 _1609_ (.A1(\gps_channel0.lo_nco.accumulator[21] ),
    .A2(_0525_),
    .B1(_0267_),
    .B2(_0501_),
    .X(_0109_));
 sky130_fd_sc_hd__or2_1 _1610_ (.A(_0240_),
    .B(\gps_channel0.lo_nco.accumulator[22] ),
    .X(_0268_));
 sky130_fd_sc_hd__nand2_1 _1611_ (.A(_0240_),
    .B(\gps_channel0.lo_nco.accumulator[22] ),
    .Y(_0269_));
 sky130_fd_sc_hd__and2_1 _1612_ (.A(_0268_),
    .B(_0269_),
    .X(_0270_));
 sky130_fd_sc_hd__o21a_1 _1613_ (.A1(\gps_channel0.lo_nco.accumulator[20] ),
    .A2(\gps_channel0.lo_nco.accumulator[21] ),
    .B1(_0245_),
    .X(_0271_));
 sky130_fd_sc_hd__a21o_1 _1614_ (.A1(_0263_),
    .A2(_0265_),
    .B1(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__or2_1 _1615_ (.A(_0270_),
    .B(_0272_),
    .X(_0273_));
 sky130_fd_sc_hd__nand2_1 _1616_ (.A(_0270_),
    .B(_0272_),
    .Y(_0274_));
 sky130_fd_sc_hd__a32o_1 _1617_ (.A1(_0501_),
    .A2(_0273_),
    .A3(_0274_),
    .B1(_0525_),
    .B2(\gps_channel0.lo_nco.accumulator[22] ),
    .X(_0110_));
 sky130_fd_sc_hd__xnor2_2 _1618_ (.A(_0240_),
    .B(\gps_channel0.lo_nco.accumulator[23] ),
    .Y(_0275_));
 sky130_fd_sc_hd__a21oi_1 _1619_ (.A1(_0269_),
    .A2(_0274_),
    .B1(_0275_),
    .Y(_0276_));
 sky130_fd_sc_hd__a31o_1 _1620_ (.A1(_0269_),
    .A2(_0274_),
    .A3(_0275_),
    .B1(_0454_),
    .X(_0277_));
 sky130_fd_sc_hd__a2bb2o_1 _1621_ (.A1_N(_0276_),
    .A2_N(_0277_),
    .B1(\gps_channel0.lo_nco.accumulator[23] ),
    .B2(_0525_),
    .X(_0111_));
 sky130_fd_sc_hd__o21a_1 _1622_ (.A1(\gps_channel0.lo_nco.accumulator[22] ),
    .A2(\gps_channel0.lo_nco.accumulator[23] ),
    .B1(_0245_),
    .X(_0278_));
 sky130_fd_sc_hd__or3_1 _1623_ (.A(_0258_),
    .B(_0271_),
    .C(_0278_),
    .X(_0279_));
 sky130_fd_sc_hd__clkinv_2 _1624_ (.A(_0275_),
    .Y(_0280_));
 sky130_fd_sc_hd__and4_1 _1625_ (.A(_0262_),
    .B(_0265_),
    .C(_0270_),
    .D(_0280_),
    .X(_0281_));
 sky130_fd_sc_hd__o211a_1 _1626_ (.A1(_0235_),
    .A2(_0238_),
    .B1(_0260_),
    .C1(_0281_),
    .X(_0282_));
 sky130_fd_sc_hd__and2_1 _1627_ (.A(_0245_),
    .B(\gps_channel0.lo_nco.accumulator[24] ),
    .X(_0283_));
 sky130_fd_sc_hd__or2_1 _1628_ (.A(_0245_),
    .B(\gps_channel0.lo_nco.accumulator[24] ),
    .X(_0284_));
 sky130_fd_sc_hd__and2b_1 _1629_ (.A_N(_0283_),
    .B(_0284_),
    .X(_0285_));
 sky130_fd_sc_hd__o21ai_1 _1630_ (.A1(_0279_),
    .A2(_0282_),
    .B1(_0285_),
    .Y(_0286_));
 sky130_fd_sc_hd__or3_1 _1631_ (.A(_0279_),
    .B(_0282_),
    .C(_0285_),
    .X(_0287_));
 sky130_fd_sc_hd__a32o_1 _1632_ (.A1(_0501_),
    .A2(_0286_),
    .A3(_0287_),
    .B1(_0451_),
    .B2(\gps_channel0.lo_nco.accumulator[24] ),
    .X(_0112_));
 sky130_fd_sc_hd__o31a_1 _1633_ (.A1(_0279_),
    .A2(_0282_),
    .A3(_0283_),
    .B1(_0284_),
    .X(_0288_));
 sky130_fd_sc_hd__and2_1 _1634_ (.A(\gps_channel0.lo_nco.accumulator[25] ),
    .B(_0288_),
    .X(_0289_));
 sky130_fd_sc_hd__a21oi_1 _1635_ (.A1(net8),
    .A2(_0288_),
    .B1(\gps_channel0.lo_nco.accumulator[25] ),
    .Y(_0290_));
 sky130_fd_sc_hd__a211oi_1 _1636_ (.A1(net8),
    .A2(_0289_),
    .B1(_0290_),
    .C1(_0450_),
    .Y(_0113_));
 sky130_fd_sc_hd__a31oi_1 _1637_ (.A1(net8),
    .A2(\gps_channel0.lo_nco.accumulator[26] ),
    .A3(_0289_),
    .B1(_0450_),
    .Y(_0291_));
 sky130_fd_sc_hd__a31o_1 _1638_ (.A1(\gps_channel0.lo_nco.accumulator[25] ),
    .A2(_0486_),
    .A3(_0288_),
    .B1(\gps_channel0.lo_nco.accumulator[26] ),
    .X(_0292_));
 sky130_fd_sc_hd__and2_1 _1639_ (.A(_0291_),
    .B(_0292_),
    .X(_0293_));
 sky130_fd_sc_hd__clkbuf_1 _1640_ (.A(_0293_),
    .X(_0114_));
 sky130_fd_sc_hd__and3_1 _1641_ (.A(\gps_channel0.lo_nco.accumulator[26] ),
    .B(_0486_),
    .C(_0289_),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _1642_ (.A0(_0294_),
    .A1(_0291_),
    .S(\gps_channel0.lo_nco.accumulator[27] ),
    .X(_0295_));
 sky130_fd_sc_hd__clkbuf_1 _1643_ (.A(_0295_),
    .X(_0115_));
 sky130_fd_sc_hd__and3_1 _1644_ (.A(\gps_channel0.lo_nco.accumulator[26] ),
    .B(\gps_channel0.lo_nco.accumulator[27] ),
    .C(_0289_),
    .X(_0296_));
 sky130_fd_sc_hd__a31oi_1 _1645_ (.A1(net8),
    .A2(\gps_channel0.lo_nco.accumulator[28] ),
    .A3(_0296_),
    .B1(_0450_),
    .Y(_0297_));
 sky130_fd_sc_hd__a21o_1 _1646_ (.A1(_0486_),
    .A2(_0296_),
    .B1(\gps_channel0.lo_nco.accumulator[28] ),
    .X(_0298_));
 sky130_fd_sc_hd__and2_1 _1647_ (.A(_0297_),
    .B(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__clkbuf_1 _1648_ (.A(_0299_),
    .X(_0116_));
 sky130_fd_sc_hd__and3_1 _1649_ (.A(\gps_channel0.lo_nco.accumulator[28] ),
    .B(_0486_),
    .C(_0296_),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _1650_ (.A0(_0300_),
    .A1(_0297_),
    .S(\gps_channel0.lo_nco.accumulator[29] ),
    .X(_0301_));
 sky130_fd_sc_hd__clkbuf_1 _1651_ (.A(_0301_),
    .X(_0117_));
 sky130_fd_sc_hd__and2_1 _1652_ (.A(\gps_channel0.lo_nco.accumulator[28] ),
    .B(\gps_channel0.lo_nco.accumulator[29] ),
    .X(_0302_));
 sky130_fd_sc_hd__a21o_1 _1653_ (.A1(_0296_),
    .A2(_0302_),
    .B1(\gps_channel0.lo_nco.accumulator[30] ),
    .X(_0303_));
 sky130_fd_sc_hd__a31oi_1 _1654_ (.A1(\gps_channel0.lo_nco.accumulator[30] ),
    .A2(_0296_),
    .A3(_0302_),
    .B1(_0454_),
    .Y(_0304_));
 sky130_fd_sc_hd__a22o_1 _1655_ (.A1(\gps_channel0.lo_nco.accumulator[30] ),
    .A2(_0525_),
    .B1(_0303_),
    .B2(_0304_),
    .X(_0118_));
 sky130_fd_sc_hd__inv_2 _1656_ (.A(\gps_channel0.lo_i ),
    .Y(_0305_));
 sky130_fd_sc_hd__a41o_1 _1657_ (.A1(\gps_channel0.lo_nco.accumulator[30] ),
    .A2(_0486_),
    .A3(_0296_),
    .A4(_0302_),
    .B1(\gps_channel0.lo_i ),
    .X(_0306_));
 sky130_fd_sc_hd__o31a_1 _1658_ (.A1(_0305_),
    .A2(_0451_),
    .A3(_0304_),
    .B1(_0306_),
    .X(_0119_));
 sky130_fd_sc_hd__and3_1 _1659_ (.A(net25),
    .B(net23),
    .C(_0206_),
    .X(_0307_));
 sky130_fd_sc_hd__buf_4 _1660_ (.A(_0307_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _1661_ (.A0(\gps_channel0.ca_gen.g2_init[1] ),
    .A1(net4),
    .S(_0308_),
    .X(_0309_));
 sky130_fd_sc_hd__or2_1 _1662_ (.A(_0213_),
    .B(_0309_),
    .X(_0310_));
 sky130_fd_sc_hd__clkbuf_1 _1663_ (.A(_0310_),
    .X(_0120_));
 sky130_fd_sc_hd__clkbuf_4 _1664_ (.A(_0220_),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _1665_ (.A0(\gps_channel0.ca_gen.g2_init[2] ),
    .A1(net5),
    .S(_0308_),
    .X(_0312_));
 sky130_fd_sc_hd__and2b_1 _1666_ (.A_N(_0311_),
    .B(_0312_),
    .X(_0313_));
 sky130_fd_sc_hd__clkbuf_1 _1667_ (.A(_0313_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _1668_ (.A0(\gps_channel0.ca_gen.g2_init[3] ),
    .A1(net6),
    .S(_0308_),
    .X(_0314_));
 sky130_fd_sc_hd__and2b_1 _1669_ (.A_N(_0311_),
    .B(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__clkbuf_1 _1670_ (.A(_0315_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _1671_ (.A0(\gps_channel0.ca_gen.g2_init[4] ),
    .A1(net7),
    .S(_0308_),
    .X(_0316_));
 sky130_fd_sc_hd__and2b_1 _1672_ (.A_N(_0311_),
    .B(_0316_),
    .X(_0317_));
 sky130_fd_sc_hd__clkbuf_1 _1673_ (.A(_0317_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _1674_ (.A0(\gps_channel0.ca_gen.g2_init[5] ),
    .A1(net9),
    .S(_0308_),
    .X(_0318_));
 sky130_fd_sc_hd__and2b_1 _1675_ (.A_N(_0311_),
    .B(_0318_),
    .X(_0319_));
 sky130_fd_sc_hd__clkbuf_1 _1676_ (.A(_0319_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _1677_ (.A0(\gps_channel0.ca_gen.g2_init[6] ),
    .A1(net10),
    .S(_0308_),
    .X(_0320_));
 sky130_fd_sc_hd__or2_1 _1678_ (.A(_0213_),
    .B(_0320_),
    .X(_0321_));
 sky130_fd_sc_hd__clkbuf_1 _1679_ (.A(_0321_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _1680_ (.A0(\gps_channel0.ca_gen.g2_init[7] ),
    .A1(net11),
    .S(_0308_),
    .X(_0322_));
 sky130_fd_sc_hd__or2_1 _1681_ (.A(_0213_),
    .B(_0322_),
    .X(_0323_));
 sky130_fd_sc_hd__clkbuf_1 _1682_ (.A(_0323_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _1683_ (.A0(\gps_channel0.ca_gen.g2_init[8] ),
    .A1(net12),
    .S(_0308_),
    .X(_0324_));
 sky130_fd_sc_hd__and2b_1 _1684_ (.A_N(_0311_),
    .B(_0324_),
    .X(_0325_));
 sky130_fd_sc_hd__clkbuf_1 _1685_ (.A(_0325_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _1686_ (.A0(\gps_channel0.ca_gen.g2_init[9] ),
    .A1(net13),
    .S(_0308_),
    .X(_0326_));
 sky130_fd_sc_hd__or2_1 _1687_ (.A(_0213_),
    .B(_0326_),
    .X(_0327_));
 sky130_fd_sc_hd__clkbuf_1 _1688_ (.A(_0327_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _1689_ (.A0(\gps_channel0.ca_gen.g2_init[10] ),
    .A1(net14),
    .S(_0308_),
    .X(_0328_));
 sky130_fd_sc_hd__and2b_1 _1690_ (.A_N(_0311_),
    .B(_0328_),
    .X(_0329_));
 sky130_fd_sc_hd__clkbuf_1 _1691_ (.A(_0329_),
    .X(_0129_));
 sky130_fd_sc_hd__inv_2 _1692_ (.A(net25),
    .Y(_0330_));
 sky130_fd_sc_hd__mux2_1 _1693_ (.A0(_0330_),
    .A1(net23),
    .S(_0206_),
    .X(_0331_));
 sky130_fd_sc_hd__and3b_1 _1694_ (.A_N(net23),
    .B(_0206_),
    .C(net25),
    .X(_0332_));
 sky130_fd_sc_hd__buf_2 _1695_ (.A(_0332_),
    .X(_0333_));
 sky130_fd_sc_hd__clkbuf_4 _1696_ (.A(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__a21oi_1 _1697_ (.A1(\gps_channel0.ca_nco.phase_sync ),
    .A2(_0331_),
    .B1(_0334_),
    .Y(_0335_));
 sky130_fd_sc_hd__nor2_1 _1698_ (.A(_0311_),
    .B(_0335_),
    .Y(_0130_));
 sky130_fd_sc_hd__o211a_1 _1699_ (.A1(_0330_),
    .A2(_0206_),
    .B1(_0207_),
    .C1(\gps_channel0.lo_nco.phase_sync ),
    .X(_0336_));
 sky130_fd_sc_hd__o21ba_1 _1700_ (.A1(_0212_),
    .A2(_0336_),
    .B1_N(_0311_),
    .X(_0131_));
 sky130_fd_sc_hd__and3_1 _1701_ (.A(_0330_),
    .B(net23),
    .C(_0206_),
    .X(_0337_));
 sky130_fd_sc_hd__clkbuf_2 _1702_ (.A(_0337_),
    .X(_0338_));
 sky130_fd_sc_hd__clkbuf_4 _1703_ (.A(_0338_),
    .X(_0339_));
 sky130_fd_sc_hd__or3b_1 _1704_ (.A(net25),
    .B(net24),
    .C_N(net23),
    .X(_0340_));
 sky130_fd_sc_hd__buf_2 _1705_ (.A(_0340_),
    .X(_0341_));
 sky130_fd_sc_hd__clkbuf_4 _1706_ (.A(_0341_),
    .X(_0342_));
 sky130_fd_sc_hd__buf_2 _1707_ (.A(net3),
    .X(_0343_));
 sky130_fd_sc_hd__o21ba_1 _1708_ (.A1(net4),
    .A2(_0342_),
    .B1_N(_0343_),
    .X(_0344_));
 sky130_fd_sc_hd__o21a_1 _1709_ (.A1(\gps_channel0.lo_nco.step[0] ),
    .A2(_0339_),
    .B1(_0344_),
    .X(_0132_));
 sky130_fd_sc_hd__o21ba_1 _1710_ (.A1(net5),
    .A2(_0342_),
    .B1_N(_0343_),
    .X(_0345_));
 sky130_fd_sc_hd__o21a_1 _1711_ (.A1(\gps_channel0.lo_nco.step[1] ),
    .A2(_0339_),
    .B1(_0345_),
    .X(_0133_));
 sky130_fd_sc_hd__o21ba_1 _1712_ (.A1(net6),
    .A2(_0342_),
    .B1_N(_0343_),
    .X(_0346_));
 sky130_fd_sc_hd__o21a_1 _1713_ (.A1(\gps_channel0.lo_nco.step[2] ),
    .A2(_0339_),
    .B1(_0346_),
    .X(_0134_));
 sky130_fd_sc_hd__o21ba_1 _1714_ (.A1(net7),
    .A2(_0342_),
    .B1_N(_0343_),
    .X(_0347_));
 sky130_fd_sc_hd__o21a_1 _1715_ (.A1(\gps_channel0.lo_nco.step[3] ),
    .A2(_0339_),
    .B1(_0347_),
    .X(_0135_));
 sky130_fd_sc_hd__o21ba_1 _1716_ (.A1(net9),
    .A2(_0342_),
    .B1_N(_0343_),
    .X(_0348_));
 sky130_fd_sc_hd__o21a_1 _1717_ (.A1(\gps_channel0.lo_nco.step[4] ),
    .A2(_0339_),
    .B1(_0348_),
    .X(_0136_));
 sky130_fd_sc_hd__o21ba_1 _1718_ (.A1(net10),
    .A2(_0342_),
    .B1_N(_0343_),
    .X(_0349_));
 sky130_fd_sc_hd__o21a_1 _1719_ (.A1(\gps_channel0.lo_nco.step[5] ),
    .A2(_0339_),
    .B1(_0349_),
    .X(_0137_));
 sky130_fd_sc_hd__o21ba_1 _1720_ (.A1(net11),
    .A2(_0342_),
    .B1_N(_0343_),
    .X(_0350_));
 sky130_fd_sc_hd__o21a_1 _1721_ (.A1(\gps_channel0.lo_nco.step[6] ),
    .A2(_0339_),
    .B1(_0350_),
    .X(_0138_));
 sky130_fd_sc_hd__o21ba_1 _1722_ (.A1(net12),
    .A2(_0342_),
    .B1_N(_0343_),
    .X(_0351_));
 sky130_fd_sc_hd__o21a_1 _1723_ (.A1(\gps_channel0.lo_nco.step[7] ),
    .A2(_0339_),
    .B1(_0351_),
    .X(_0139_));
 sky130_fd_sc_hd__o21ba_1 _1724_ (.A1(net13),
    .A2(_0342_),
    .B1_N(_0343_),
    .X(_0352_));
 sky130_fd_sc_hd__o21a_1 _1725_ (.A1(\gps_channel0.lo_nco.step[8] ),
    .A2(_0339_),
    .B1(_0352_),
    .X(_0140_));
 sky130_fd_sc_hd__o21ba_1 _1726_ (.A1(net14),
    .A2(_0341_),
    .B1_N(_0343_),
    .X(_0353_));
 sky130_fd_sc_hd__o21a_1 _1727_ (.A1(\gps_channel0.lo_nco.step[9] ),
    .A2(_0339_),
    .B1(_0353_),
    .X(_0141_));
 sky130_fd_sc_hd__buf_2 _1728_ (.A(net3),
    .X(_0354_));
 sky130_fd_sc_hd__o21ba_1 _1729_ (.A1(net15),
    .A2(_0341_),
    .B1_N(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__o21a_1 _1730_ (.A1(\gps_channel0.lo_nco.step[10] ),
    .A2(_0338_),
    .B1(_0355_),
    .X(_0142_));
 sky130_fd_sc_hd__o21ba_1 _1731_ (.A1(net16),
    .A2(_0341_),
    .B1_N(_0354_),
    .X(_0356_));
 sky130_fd_sc_hd__o21a_1 _1732_ (.A1(\gps_channel0.lo_nco.step[11] ),
    .A2(_0338_),
    .B1(_0356_),
    .X(_0143_));
 sky130_fd_sc_hd__o21ba_1 _1733_ (.A1(net17),
    .A2(_0341_),
    .B1_N(_0354_),
    .X(_0357_));
 sky130_fd_sc_hd__o21a_1 _1734_ (.A1(\gps_channel0.lo_nco.step[12] ),
    .A2(_0338_),
    .B1(_0357_),
    .X(_0144_));
 sky130_fd_sc_hd__o21ba_1 _1735_ (.A1(net18),
    .A2(_0341_),
    .B1_N(_0354_),
    .X(_0358_));
 sky130_fd_sc_hd__o21a_1 _1736_ (.A1(\gps_channel0.lo_nco.step[13] ),
    .A2(_0338_),
    .B1(_0358_),
    .X(_0145_));
 sky130_fd_sc_hd__o21ba_1 _1737_ (.A1(net20),
    .A2(_0341_),
    .B1_N(_0354_),
    .X(_0359_));
 sky130_fd_sc_hd__o21a_1 _1738_ (.A1(\gps_channel0.lo_nco.step[14] ),
    .A2(_0338_),
    .B1(_0359_),
    .X(_0146_));
 sky130_fd_sc_hd__o21ba_1 _1739_ (.A1(net21),
    .A2(_0341_),
    .B1_N(_0354_),
    .X(_0360_));
 sky130_fd_sc_hd__o21a_1 _1740_ (.A1(\gps_channel0.lo_nco.step[15] ),
    .A2(_0338_),
    .B1(_0360_),
    .X(_0147_));
 sky130_fd_sc_hd__a21o_1 _1741_ (.A1(_0245_),
    .A2(_0342_),
    .B1(_0311_),
    .X(_0148_));
 sky130_fd_sc_hd__or3b_1 _1742_ (.A(_0206_),
    .B(net25),
    .C_N(net23),
    .X(_0361_));
 sky130_fd_sc_hd__clkbuf_4 _1743_ (.A(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__clkbuf_4 _1744_ (.A(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__and3_2 _1745_ (.A(_0330_),
    .B(net23),
    .C(net24),
    .X(_0364_));
 sky130_fd_sc_hd__clkbuf_4 _1746_ (.A(_0364_),
    .X(_0365_));
 sky130_fd_sc_hd__o21ba_1 _1747_ (.A1(\gps_channel0.ca_nco.step[0] ),
    .A2(_0365_),
    .B1_N(_0354_),
    .X(_0366_));
 sky130_fd_sc_hd__o21a_1 _1748_ (.A1(net4),
    .A2(_0363_),
    .B1(_0366_),
    .X(_0149_));
 sky130_fd_sc_hd__o21ba_1 _1749_ (.A1(\gps_channel0.ca_nco.step[1] ),
    .A2(_0365_),
    .B1_N(_0354_),
    .X(_0367_));
 sky130_fd_sc_hd__o21a_1 _1750_ (.A1(net5),
    .A2(_0363_),
    .B1(_0367_),
    .X(_0150_));
 sky130_fd_sc_hd__o21ba_1 _1751_ (.A1(\gps_channel0.ca_nco.step[2] ),
    .A2(_0365_),
    .B1_N(_0354_),
    .X(_0368_));
 sky130_fd_sc_hd__o21a_1 _1752_ (.A1(net6),
    .A2(_0363_),
    .B1(_0368_),
    .X(_0151_));
 sky130_fd_sc_hd__o21ba_1 _1753_ (.A1(\gps_channel0.ca_nco.step[3] ),
    .A2(_0365_),
    .B1_N(_0354_),
    .X(_0369_));
 sky130_fd_sc_hd__o21a_1 _1754_ (.A1(net7),
    .A2(_0363_),
    .B1(_0369_),
    .X(_0152_));
 sky130_fd_sc_hd__buf_2 _1755_ (.A(net3),
    .X(_0370_));
 sky130_fd_sc_hd__o21ba_1 _1756_ (.A1(\gps_channel0.ca_nco.step[4] ),
    .A2(_0365_),
    .B1_N(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__o21a_1 _1757_ (.A1(net9),
    .A2(_0363_),
    .B1(_0371_),
    .X(_0153_));
 sky130_fd_sc_hd__o21ba_1 _1758_ (.A1(\gps_channel0.ca_nco.step[5] ),
    .A2(_0365_),
    .B1_N(_0370_),
    .X(_0372_));
 sky130_fd_sc_hd__o21a_1 _1759_ (.A1(net10),
    .A2(_0363_),
    .B1(_0372_),
    .X(_0154_));
 sky130_fd_sc_hd__o21ba_1 _1760_ (.A1(\gps_channel0.ca_nco.step[6] ),
    .A2(_0365_),
    .B1_N(_0370_),
    .X(_0373_));
 sky130_fd_sc_hd__o21a_1 _1761_ (.A1(net11),
    .A2(_0363_),
    .B1(_0373_),
    .X(_0155_));
 sky130_fd_sc_hd__o21ba_1 _1762_ (.A1(\gps_channel0.ca_nco.step[7] ),
    .A2(_0365_),
    .B1_N(_0370_),
    .X(_0374_));
 sky130_fd_sc_hd__o21a_1 _1763_ (.A1(net12),
    .A2(_0363_),
    .B1(_0374_),
    .X(_0156_));
 sky130_fd_sc_hd__o21ba_1 _1764_ (.A1(\gps_channel0.ca_nco.step[8] ),
    .A2(_0365_),
    .B1_N(_0370_),
    .X(_0375_));
 sky130_fd_sc_hd__o21a_1 _1765_ (.A1(net13),
    .A2(_0363_),
    .B1(_0375_),
    .X(_0157_));
 sky130_fd_sc_hd__o21ba_1 _1766_ (.A1(\gps_channel0.ca_nco.step[9] ),
    .A2(_0365_),
    .B1_N(_0370_),
    .X(_0376_));
 sky130_fd_sc_hd__o21a_1 _1767_ (.A1(net14),
    .A2(_0363_),
    .B1(_0376_),
    .X(_0158_));
 sky130_fd_sc_hd__o21ba_1 _1768_ (.A1(\gps_channel0.ca_nco.step[10] ),
    .A2(_0364_),
    .B1_N(_0370_),
    .X(_0377_));
 sky130_fd_sc_hd__o21a_1 _1769_ (.A1(net15),
    .A2(_0362_),
    .B1(_0377_),
    .X(_0159_));
 sky130_fd_sc_hd__o21ba_1 _1770_ (.A1(\gps_channel0.ca_nco.step[11] ),
    .A2(_0364_),
    .B1_N(_0370_),
    .X(_0378_));
 sky130_fd_sc_hd__o21a_1 _1771_ (.A1(net16),
    .A2(_0362_),
    .B1(_0378_),
    .X(_0160_));
 sky130_fd_sc_hd__o21ba_1 _1772_ (.A1(\gps_channel0.ca_nco.step[12] ),
    .A2(_0364_),
    .B1_N(_0370_),
    .X(_0379_));
 sky130_fd_sc_hd__o21a_1 _1773_ (.A1(net17),
    .A2(_0362_),
    .B1(_0379_),
    .X(_0161_));
 sky130_fd_sc_hd__o21ba_1 _1774_ (.A1(\gps_channel0.ca_nco.step[13] ),
    .A2(_0364_),
    .B1_N(_0370_),
    .X(_0380_));
 sky130_fd_sc_hd__o21a_1 _1775_ (.A1(net18),
    .A2(_0362_),
    .B1(_0380_),
    .X(_0162_));
 sky130_fd_sc_hd__buf_2 _1776_ (.A(net3),
    .X(_0381_));
 sky130_fd_sc_hd__o21ba_1 _1777_ (.A1(\gps_channel0.ca_nco.step[14] ),
    .A2(_0364_),
    .B1_N(_0381_),
    .X(_0382_));
 sky130_fd_sc_hd__o21a_1 _1778_ (.A1(net20),
    .A2(_0362_),
    .B1(_0382_),
    .X(_0163_));
 sky130_fd_sc_hd__o21ba_1 _1779_ (.A1(\gps_channel0.ca_nco.step[15] ),
    .A2(_0364_),
    .B1_N(_0381_),
    .X(_0383_));
 sky130_fd_sc_hd__o21a_1 _1780_ (.A1(net21),
    .A2(_0362_),
    .B1(_0383_),
    .X(_0164_));
 sky130_fd_sc_hd__a21o_1 _1781_ (.A1(_0640_),
    .A2(_0362_),
    .B1(_0311_),
    .X(_0165_));
 sky130_fd_sc_hd__or3_1 _1782_ (.A(_0330_),
    .B(net23),
    .C(net24),
    .X(_0384_));
 sky130_fd_sc_hd__buf_2 _1783_ (.A(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__buf_2 _1784_ (.A(_0385_),
    .X(_0386_));
 sky130_fd_sc_hd__o21ba_1 _1785_ (.A1(\gps_channel0.ca_nco.phase_in[0] ),
    .A2(_0334_),
    .B1_N(_0381_),
    .X(_0387_));
 sky130_fd_sc_hd__o21a_1 _1786_ (.A1(net4),
    .A2(_0386_),
    .B1(_0387_),
    .X(_0166_));
 sky130_fd_sc_hd__o21ba_1 _1787_ (.A1(\gps_channel0.ca_nco.phase_in[1] ),
    .A2(_0334_),
    .B1_N(_0381_),
    .X(_0388_));
 sky130_fd_sc_hd__o21a_1 _1788_ (.A1(net5),
    .A2(_0386_),
    .B1(_0388_),
    .X(_0167_));
 sky130_fd_sc_hd__o21ba_1 _1789_ (.A1(\gps_channel0.ca_nco.phase_in[2] ),
    .A2(_0334_),
    .B1_N(_0381_),
    .X(_0389_));
 sky130_fd_sc_hd__o21a_1 _1790_ (.A1(net6),
    .A2(_0386_),
    .B1(_0389_),
    .X(_0168_));
 sky130_fd_sc_hd__o21ba_1 _1791_ (.A1(\gps_channel0.ca_nco.phase_in[3] ),
    .A2(_0334_),
    .B1_N(_0381_),
    .X(_0390_));
 sky130_fd_sc_hd__o21a_1 _1792_ (.A1(net7),
    .A2(_0386_),
    .B1(_0390_),
    .X(_0169_));
 sky130_fd_sc_hd__o21ba_1 _1793_ (.A1(\gps_channel0.ca_nco.phase_in[4] ),
    .A2(_0334_),
    .B1_N(_0381_),
    .X(_0391_));
 sky130_fd_sc_hd__o21a_1 _1794_ (.A1(net9),
    .A2(_0386_),
    .B1(_0391_),
    .X(_0170_));
 sky130_fd_sc_hd__o21ba_1 _1795_ (.A1(\gps_channel0.ca_nco.phase_in[5] ),
    .A2(_0334_),
    .B1_N(_0381_),
    .X(_0392_));
 sky130_fd_sc_hd__o21a_1 _1796_ (.A1(net10),
    .A2(_0386_),
    .B1(_0392_),
    .X(_0171_));
 sky130_fd_sc_hd__o21ba_1 _1797_ (.A1(\gps_channel0.ca_nco.phase_in[6] ),
    .A2(_0334_),
    .B1_N(_0381_),
    .X(_0393_));
 sky130_fd_sc_hd__o21a_1 _1798_ (.A1(net11),
    .A2(_0386_),
    .B1(_0393_),
    .X(_0172_));
 sky130_fd_sc_hd__o21ba_1 _1799_ (.A1(\gps_channel0.ca_nco.phase_in[7] ),
    .A2(_0334_),
    .B1_N(_0381_),
    .X(_0394_));
 sky130_fd_sc_hd__o21a_1 _1800_ (.A1(net12),
    .A2(_0386_),
    .B1(_0394_),
    .X(_0173_));
 sky130_fd_sc_hd__o21ba_1 _1801_ (.A1(\gps_channel0.ca_nco.phase_in[8] ),
    .A2(_0334_),
    .B1_N(_0220_),
    .X(_0395_));
 sky130_fd_sc_hd__o21a_1 _1802_ (.A1(net13),
    .A2(_0386_),
    .B1(_0395_),
    .X(_0174_));
 sky130_fd_sc_hd__o21ba_1 _1803_ (.A1(\gps_channel0.ca_nco.phase_in[9] ),
    .A2(_0333_),
    .B1_N(_0220_),
    .X(_0396_));
 sky130_fd_sc_hd__o21a_1 _1804_ (.A1(net14),
    .A2(_0386_),
    .B1(_0396_),
    .X(_0175_));
 sky130_fd_sc_hd__o21ba_1 _1805_ (.A1(\gps_channel0.ca_nco.phase_in[10] ),
    .A2(_0333_),
    .B1_N(_0220_),
    .X(_0397_));
 sky130_fd_sc_hd__o21a_1 _1806_ (.A1(net15),
    .A2(_0385_),
    .B1(_0397_),
    .X(_0176_));
 sky130_fd_sc_hd__o21ba_1 _1807_ (.A1(\gps_channel0.ca_nco.phase_in[11] ),
    .A2(_0333_),
    .B1_N(_0220_),
    .X(_0398_));
 sky130_fd_sc_hd__o21a_1 _1808_ (.A1(net16),
    .A2(_0385_),
    .B1(_0398_),
    .X(_0177_));
 sky130_fd_sc_hd__o21ba_1 _1809_ (.A1(\gps_channel0.ca_nco.phase_in[12] ),
    .A2(_0333_),
    .B1_N(_0220_),
    .X(_0399_));
 sky130_fd_sc_hd__o21a_1 _1810_ (.A1(net17),
    .A2(_0385_),
    .B1(_0399_),
    .X(_0178_));
 sky130_fd_sc_hd__o21ba_1 _1811_ (.A1(\gps_channel0.ca_nco.phase_in[13] ),
    .A2(_0333_),
    .B1_N(_0220_),
    .X(_0400_));
 sky130_fd_sc_hd__o21a_1 _1812_ (.A1(net18),
    .A2(_0385_),
    .B1(_0400_),
    .X(_0179_));
 sky130_fd_sc_hd__o21ba_1 _1813_ (.A1(\gps_channel0.ca_nco.phase_in[14] ),
    .A2(_0333_),
    .B1_N(_0220_),
    .X(_0401_));
 sky130_fd_sc_hd__o21a_1 _1814_ (.A1(net20),
    .A2(_0385_),
    .B1(_0401_),
    .X(_0180_));
 sky130_fd_sc_hd__o21ba_1 _1815_ (.A1(\gps_channel0.ca_nco.phase_in[15] ),
    .A2(_0333_),
    .B1_N(_0220_),
    .X(_0402_));
 sky130_fd_sc_hd__o21a_1 _1816_ (.A1(net21),
    .A2(_0385_),
    .B1(_0402_),
    .X(_0181_));
 sky130_fd_sc_hd__dfxtp_1 _1817_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0030_),
    .Q(\gps_channel0.lo_nco.accumulator[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1818_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0031_),
    .Q(\gps_channel0.lo_nco.accumulator[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1819_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0032_),
    .Q(\gps_channel0.lo_nco.accumulator[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1820_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0033_),
    .Q(\gps_channel0.lo_nco.accumulator[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1821_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0034_),
    .Q(\gps_channel0.lo_nco.accumulator[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1822_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0035_),
    .Q(\gps_channel0.lo_nco.accumulator[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1823_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0036_),
    .Q(\gps_channel0.lo_nco.accumulator[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1824_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0037_),
    .Q(\gps_channel0.lo_nco.accumulator[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1825_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0038_),
    .Q(\gps_channel0.lo_nco.accumulator[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1826_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0039_),
    .Q(\gps_channel0.lo_nco.accumulator[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1827_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0040_),
    .Q(\gps_channel0.lo_nco.accumulator[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1828_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0041_),
    .Q(\gps_channel0.lo_nco.accumulator[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1829_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0042_),
    .Q(\gps_channel0.lo_nco.accumulator[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1830_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0043_),
    .Q(\gps_channel0.lo_nco.accumulator[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1831_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0044_),
    .Q(\gps_channel0.lo_nco.accumulator[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1832_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0045_),
    .Q(\gps_channel0.lo_nco.accumulator[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1833_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0046_),
    .Q(\gps_channel0.ca_nco.accumulator[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1834_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0047_),
    .Q(\gps_channel0.ca_nco.accumulator[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1835_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0048_),
    .Q(\gps_channel0.ca_nco.accumulator[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1836_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0049_),
    .Q(\gps_channel0.ca_nco.accumulator[19] ));
 sky130_fd_sc_hd__dfxtp_1 _1837_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0050_),
    .Q(\gps_channel0.ca_nco.accumulator[20] ));
 sky130_fd_sc_hd__dfxtp_1 _1838_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0051_),
    .Q(\gps_channel0.ca_nco.accumulator[21] ));
 sky130_fd_sc_hd__dfxtp_1 _1839_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0052_),
    .Q(\gps_channel0.ca_nco.accumulator[22] ));
 sky130_fd_sc_hd__dfxtp_1 _1840_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0053_),
    .Q(\gps_channel0.ca_nco.accumulator[23] ));
 sky130_fd_sc_hd__dfxtp_1 _1841_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0054_),
    .Q(\gps_channel0.ca_nco.accumulator[24] ));
 sky130_fd_sc_hd__dfxtp_1 _1842_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0055_),
    .Q(\gps_channel0.ca_nco.accumulator[25] ));
 sky130_fd_sc_hd__dfxtp_1 _1843_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0056_),
    .Q(\gps_channel0.ca_nco.accumulator[26] ));
 sky130_fd_sc_hd__dfxtp_1 _1844_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0057_),
    .Q(\gps_channel0.ca_nco.accumulator[27] ));
 sky130_fd_sc_hd__dfxtp_1 _1845_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0058_),
    .Q(\gps_channel0.ca_nco.accumulator[28] ));
 sky130_fd_sc_hd__dfxtp_1 _1846_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0059_),
    .Q(\gps_channel0.ca_nco.accumulator[29] ));
 sky130_fd_sc_hd__dfxtp_1 _1847_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0060_),
    .Q(\gps_channel0.ca_nco.accumulator[30] ));
 sky130_fd_sc_hd__dfxtp_1 _1848_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0061_),
    .Q(\gps_channel0.ca_nco.accumulator[31] ));
 sky130_fd_sc_hd__dfxtp_1 _1849_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0062_),
    .Q(\gps_channel0.ca_nco.accumulator[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1850_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0063_),
    .Q(\gps_channel0.ca_nco.accumulator[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1851_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0064_),
    .Q(\gps_channel0.ca_nco.accumulator[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1852_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0065_),
    .Q(\gps_channel0.ca_nco.accumulator[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1853_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0066_),
    .Q(\gps_channel0.ca_nco.accumulator[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1854_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0067_),
    .Q(\gps_channel0.ca_nco.accumulator[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1855_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0068_),
    .Q(\gps_channel0.ca_nco.accumulator[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1856_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0069_),
    .Q(\gps_channel0.ca_nco.accumulator[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1857_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0070_),
    .Q(\gps_channel0.ca_nco.accumulator[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1858_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0071_),
    .Q(\gps_channel0.ca_nco.accumulator[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1859_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0072_),
    .Q(\gps_channel0.ca_nco.accumulator[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1860_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0073_),
    .Q(\gps_channel0.ca_nco.accumulator[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1861_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0074_),
    .Q(\gps_channel0.ca_nco.accumulator[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1862_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0075_),
    .Q(\gps_channel0.ca_nco.accumulator[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1863_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0076_),
    .Q(\gps_channel0.ca_nco.accumulator[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1864_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0077_),
    .Q(\gps_channel0.ca_nco.accumulator[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1865_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0078_),
    .Q(\gps_channel0.lo_nco.phase_in[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1866_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0079_),
    .Q(\gps_channel0.lo_nco.phase_in[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1867_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0080_),
    .Q(\gps_channel0.lo_nco.phase_in[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1868_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0081_),
    .Q(\gps_channel0.lo_nco.phase_in[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1869_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0082_),
    .Q(\gps_channel0.lo_nco.phase_in[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1870_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0083_),
    .Q(\gps_channel0.lo_nco.phase_in[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1871_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0084_),
    .Q(\gps_channel0.lo_nco.phase_in[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1872_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0085_),
    .Q(\gps_channel0.lo_nco.phase_in[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1873_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0086_),
    .Q(\gps_channel0.lo_nco.phase_in[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1874_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0087_),
    .Q(\gps_channel0.lo_nco.phase_in[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1875_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0088_),
    .Q(\gps_channel0.lo_nco.phase_in[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1876_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0089_),
    .Q(\gps_channel0.lo_nco.phase_in[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1877_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0090_),
    .Q(\gps_channel0.lo_nco.phase_in[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1878_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0091_),
    .Q(\gps_channel0.lo_nco.phase_in[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1879_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0092_),
    .Q(\gps_channel0.lo_nco.phase_in[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1880_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0093_),
    .Q(\gps_channel0.lo_nco.phase_in[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1881_ (.CLK(_0010_),
    .D(_0000_),
    .Q(\gps_channel0.ca_gen.g2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1882_ (.CLK(_0011_),
    .D(_0001_),
    .Q(\gps_channel0.ca_gen.g2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1883_ (.CLK(_0012_),
    .D(_0002_),
    .Q(\gps_channel0.ca_gen.g2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1884_ (.CLK(_0013_),
    .D(_0003_),
    .Q(\gps_channel0.ca_gen.g2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1885_ (.CLK(_0014_),
    .D(_0004_),
    .Q(\gps_channel0.ca_gen.g2[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1886_ (.CLK(_0015_),
    .D(_0005_),
    .Q(\gps_channel0.ca_gen.g2[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1887_ (.CLK(_0016_),
    .D(_0006_),
    .Q(\gps_channel0.ca_gen.g2[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1888_ (.CLK(_0017_),
    .D(_0007_),
    .Q(\gps_channel0.ca_gen.g2[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1889_ (.CLK(_0018_),
    .D(_0008_),
    .Q(\gps_channel0.ca_gen.g2[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1890_ (.CLK(_0019_),
    .D(_0009_),
    .Q(\gps_channel0.ca_gen.g2[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1891_ (.CLK(_0020_),
    .D(_0094_),
    .Q(\gps_channel0.ca_gen.g1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1892_ (.CLK(_0021_),
    .D(_0095_),
    .Q(\gps_channel0.ca_gen.g1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1893_ (.CLK(_0022_),
    .D(_0096_),
    .Q(\gps_channel0.ca_gen.g1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1894_ (.CLK(_0023_),
    .D(_0097_),
    .Q(\gps_channel0.ca_gen.g1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1895_ (.CLK(_0024_),
    .D(_0098_),
    .Q(\gps_channel0.ca_gen.g1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1896_ (.CLK(_0025_),
    .D(_0099_),
    .Q(\gps_channel0.ca_gen.g1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1897_ (.CLK(_0026_),
    .D(_0100_),
    .Q(\gps_channel0.ca_gen.g1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1898_ (.CLK(_0027_),
    .D(_0101_),
    .Q(\gps_channel0.ca_gen.g1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1899_ (.CLK(_0028_),
    .D(_0102_),
    .Q(\gps_channel0.ca_gen.g1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1900_ (.CLK(_0029_),
    .D(_0103_),
    .Q(\gps_channel0.ca_gen.g1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1901_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0104_),
    .Q(\gps_channel0.lo_nco.accumulator[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1902_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0105_),
    .Q(\gps_channel0.lo_nco.accumulator[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1903_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0106_),
    .Q(\gps_channel0.lo_nco.accumulator[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1904_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0107_),
    .Q(\gps_channel0.lo_nco.accumulator[19] ));
 sky130_fd_sc_hd__dfxtp_1 _1905_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0108_),
    .Q(\gps_channel0.lo_nco.accumulator[20] ));
 sky130_fd_sc_hd__dfxtp_1 _1906_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0109_),
    .Q(\gps_channel0.lo_nco.accumulator[21] ));
 sky130_fd_sc_hd__dfxtp_1 _1907_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0110_),
    .Q(\gps_channel0.lo_nco.accumulator[22] ));
 sky130_fd_sc_hd__dfxtp_1 _1908_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0111_),
    .Q(\gps_channel0.lo_nco.accumulator[23] ));
 sky130_fd_sc_hd__dfxtp_1 _1909_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0112_),
    .Q(\gps_channel0.lo_nco.accumulator[24] ));
 sky130_fd_sc_hd__dfxtp_1 _1910_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0113_),
    .Q(\gps_channel0.lo_nco.accumulator[25] ));
 sky130_fd_sc_hd__dfxtp_1 _1911_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0114_),
    .Q(\gps_channel0.lo_nco.accumulator[26] ));
 sky130_fd_sc_hd__dfxtp_1 _1912_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0115_),
    .Q(\gps_channel0.lo_nco.accumulator[27] ));
 sky130_fd_sc_hd__dfxtp_1 _1913_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0116_),
    .Q(\gps_channel0.lo_nco.accumulator[28] ));
 sky130_fd_sc_hd__dfxtp_1 _1914_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0117_),
    .Q(\gps_channel0.lo_nco.accumulator[29] ));
 sky130_fd_sc_hd__dfxtp_2 _1915_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0118_),
    .Q(\gps_channel0.lo_nco.accumulator[30] ));
 sky130_fd_sc_hd__dfxtp_4 _1916_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0119_),
    .Q(\gps_channel0.lo_i ));
 sky130_fd_sc_hd__dfxtp_1 _1917_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0120_),
    .Q(\gps_channel0.ca_gen.g2_init[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1918_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0121_),
    .Q(\gps_channel0.ca_gen.g2_init[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1919_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0122_),
    .Q(\gps_channel0.ca_gen.g2_init[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1920_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0123_),
    .Q(\gps_channel0.ca_gen.g2_init[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1921_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0124_),
    .Q(\gps_channel0.ca_gen.g2_init[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1922_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0125_),
    .Q(\gps_channel0.ca_gen.g2_init[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1923_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0126_),
    .Q(\gps_channel0.ca_gen.g2_init[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1924_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0127_),
    .Q(\gps_channel0.ca_gen.g2_init[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1925_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0128_),
    .Q(\gps_channel0.ca_gen.g2_init[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1926_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0129_),
    .Q(\gps_channel0.ca_gen.g2_init[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1927_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0130_),
    .Q(\gps_channel0.ca_nco.phase_sync ));
 sky130_fd_sc_hd__dfxtp_1 _1928_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0131_),
    .Q(\gps_channel0.lo_nco.phase_sync ));
 sky130_fd_sc_hd__dfxtp_1 _1929_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0132_),
    .Q(\gps_channel0.lo_nco.step[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1930_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0133_),
    .Q(\gps_channel0.lo_nco.step[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1931_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0134_),
    .Q(\gps_channel0.lo_nco.step[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1932_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0135_),
    .Q(\gps_channel0.lo_nco.step[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1933_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0136_),
    .Q(\gps_channel0.lo_nco.step[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1934_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0137_),
    .Q(\gps_channel0.lo_nco.step[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1935_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0138_),
    .Q(\gps_channel0.lo_nco.step[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1936_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0139_),
    .Q(\gps_channel0.lo_nco.step[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1937_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0140_),
    .Q(\gps_channel0.lo_nco.step[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1938_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0141_),
    .Q(\gps_channel0.lo_nco.step[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1939_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0142_),
    .Q(\gps_channel0.lo_nco.step[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1940_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0143_),
    .Q(\gps_channel0.lo_nco.step[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1941_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0144_),
    .Q(\gps_channel0.lo_nco.step[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1942_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0145_),
    .Q(\gps_channel0.lo_nco.step[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1943_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0146_),
    .Q(\gps_channel0.lo_nco.step[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1944_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0147_),
    .Q(\gps_channel0.lo_nco.step[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1945_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0148_),
    .Q(\gps_channel0.lo_nco.step[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1946_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0149_),
    .Q(\gps_channel0.ca_nco.step[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1947_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0150_),
    .Q(\gps_channel0.ca_nco.step[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1948_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0151_),
    .Q(\gps_channel0.ca_nco.step[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1949_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0152_),
    .Q(\gps_channel0.ca_nco.step[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1950_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0153_),
    .Q(\gps_channel0.ca_nco.step[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1951_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0154_),
    .Q(\gps_channel0.ca_nco.step[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1952_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0155_),
    .Q(\gps_channel0.ca_nco.step[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1953_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0156_),
    .Q(\gps_channel0.ca_nco.step[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1954_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0157_),
    .Q(\gps_channel0.ca_nco.step[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1955_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0158_),
    .Q(\gps_channel0.ca_nco.step[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1956_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0159_),
    .Q(\gps_channel0.ca_nco.step[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1957_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0160_),
    .Q(\gps_channel0.ca_nco.step[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1958_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0161_),
    .Q(\gps_channel0.ca_nco.step[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1959_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0162_),
    .Q(\gps_channel0.ca_nco.step[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1960_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0163_),
    .Q(\gps_channel0.ca_nco.step[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1961_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0164_),
    .Q(\gps_channel0.ca_nco.step[15] ));
 sky130_fd_sc_hd__dfxtp_2 _1962_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0165_),
    .Q(\gps_channel0.ca_nco.step[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1963_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0166_),
    .Q(\gps_channel0.ca_nco.phase_in[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1964_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0167_),
    .Q(\gps_channel0.ca_nco.phase_in[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1965_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0168_),
    .Q(\gps_channel0.ca_nco.phase_in[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1966_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0169_),
    .Q(\gps_channel0.ca_nco.phase_in[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1967_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0170_),
    .Q(\gps_channel0.ca_nco.phase_in[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1968_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0171_),
    .Q(\gps_channel0.ca_nco.phase_in[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1969_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0172_),
    .Q(\gps_channel0.ca_nco.phase_in[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1970_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0173_),
    .Q(\gps_channel0.ca_nco.phase_in[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1971_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0174_),
    .Q(\gps_channel0.ca_nco.phase_in[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1972_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0175_),
    .Q(\gps_channel0.ca_nco.phase_in[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1973_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0176_),
    .Q(\gps_channel0.ca_nco.phase_in[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1974_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0177_),
    .Q(\gps_channel0.ca_nco.phase_in[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1975_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0178_),
    .Q(\gps_channel0.ca_nco.phase_in[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1976_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0179_),
    .Q(\gps_channel0.ca_nco.phase_in[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1977_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0180_),
    .Q(\gps_channel0.ca_nco.phase_in[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1978_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0181_),
    .Q(\gps_channel0.ca_nco.phase_in[15] ));
 sky130_fd_sc_hd__conb_1 _2077__27 (.LO(net27));
 sky130_fd_sc_hd__conb_1 _2078__28 (.LO(net28));
 sky130_fd_sc_hd__conb_1 _2079__29 (.LO(net29));
 sky130_fd_sc_hd__conb_1 _2080__30 (.LO(net30));
 sky130_fd_sc_hd__conb_1 _2081__31 (.LO(net31));
 sky130_fd_sc_hd__conb_1 _2082__32 (.LO(net32));
 sky130_fd_sc_hd__conb_1 _2092__33 (.LO(net33));
 sky130_fd_sc_hd__conb_1 _2093__34 (.LO(net34));
 sky130_fd_sc_hd__conb_1 _2094__35 (.LO(net35));
 sky130_fd_sc_hd__conb_1 _2095__36 (.LO(net36));
 sky130_fd_sc_hd__conb_1 _2096__37 (.LO(net37));
 sky130_fd_sc_hd__conb_1 _2097__38 (.LO(net38));
 sky130_fd_sc_hd__conb_1 _2098__39 (.LO(net39));
 sky130_fd_sc_hd__conb_1 _2099__40 (.LO(net40));
 sky130_fd_sc_hd__conb_1 _2100__41 (.LO(net41));
 sky130_fd_sc_hd__conb_1 _2101__42 (.LO(net42));
 sky130_fd_sc_hd__conb_1 _2102__43 (.LO(net43));
 sky130_fd_sc_hd__conb_1 _2103__44 (.LO(net44));
 sky130_fd_sc_hd__conb_1 _2104__45 (.LO(net45));
 sky130_fd_sc_hd__conb_1 _2105__46 (.LO(net46));
 sky130_fd_sc_hd__conb_1 _2106__47 (.LO(net47));
 sky130_fd_sc_hd__conb_1 _2107__48 (.LO(net48));
 sky130_fd_sc_hd__conb_1 _2108__49 (.LO(net49));
 sky130_fd_sc_hd__conb_1 _2109__50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 _2110__51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 _2111__52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 _2112__53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 _2113__54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 _2114__55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 _2115__56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 _2116__57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 _2117__58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 _2118__59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 _2119__60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 _2120__61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 _2121__62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 _2122__63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 _2123__64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 _2124__65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 _2125__66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 _2126__67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 _2128__68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 _2130__69 (.LO(net69));
 sky130_fd_sc_hd__conb_1 _2131__70 (.LO(net70));
 sky130_fd_sc_hd__conb_1 _2132__71 (.LO(net71));
 sky130_fd_sc_hd__conb_1 _2133__72 (.LO(net72));
 sky130_fd_sc_hd__conb_1 _2134__73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 _2135__74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 _2136__75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 _2137__76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 _2138__77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 _2139__78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 _2140__79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 _2141__80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 _2142__81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 _2143__82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 _2144__83 (.LO(net83));
 sky130_fd_sc_hd__conb_1 _2145__84 (.LO(net84));
 sky130_fd_sc_hd__conb_1 _2146__85 (.LO(net85));
 sky130_fd_sc_hd__conb_1 _2147__86 (.LO(net86));
 sky130_fd_sc_hd__conb_1 _2148__87 (.LO(net87));
 sky130_fd_sc_hd__conb_1 _2149__88 (.LO(net88));
 sky130_fd_sc_hd__conb_1 _2150__89 (.LO(net89));
 sky130_fd_sc_hd__conb_1 _2151__90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 _2152__91 (.LO(net91));
 sky130_fd_sc_hd__conb_1 _2153__92 (.LO(net92));
 sky130_fd_sc_hd__conb_1 _2154__93 (.LO(net93));
 sky130_fd_sc_hd__conb_1 _2155__94 (.LO(net94));
 sky130_fd_sc_hd__conb_1 _2156__95 (.LO(net95));
 sky130_fd_sc_hd__conb_1 _2157__96 (.LO(net96));
 sky130_fd_sc_hd__conb_1 _2158__97 (.LO(net97));
 sky130_fd_sc_hd__conb_1 _2159__98 (.LO(net98));
 sky130_fd_sc_hd__conb_1 _2160__99 (.LO(net99));
 sky130_fd_sc_hd__conb_1 _2161__100 (.LO(net100));
 sky130_fd_sc_hd__conb_1 _2162__101 (.LO(net101));
 sky130_fd_sc_hd__conb_1 _2163__102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 _2164__103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 _2165__104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 _2166__105 (.LO(net105));
 sky130_fd_sc_hd__conb_1 _2167__106 (.LO(net106));
 sky130_fd_sc_hd__conb_1 _2168__107 (.LO(net107));
 sky130_fd_sc_hd__conb_1 _2169__108 (.LO(net108));
 sky130_fd_sc_hd__conb_1 _2170__109 (.LO(net109));
 sky130_fd_sc_hd__conb_1 _2171__110 (.LO(net110));
 sky130_fd_sc_hd__conb_1 _2172__111 (.LO(net111));
 sky130_fd_sc_hd__conb_1 _2173__112 (.LO(net112));
 sky130_fd_sc_hd__conb_1 _2174__113 (.LO(net113));
 sky130_fd_sc_hd__conb_1 _2175__114 (.LO(net114));
 sky130_fd_sc_hd__conb_1 _2176__115 (.LO(net115));
 sky130_fd_sc_hd__conb_1 _2177__116 (.LO(net116));
 sky130_fd_sc_hd__conb_1 _2178__117 (.LO(net117));
 sky130_fd_sc_hd__conb_1 _2179__118 (.LO(net118));
 sky130_fd_sc_hd__conb_1 _2180__119 (.LO(net119));
 sky130_fd_sc_hd__conb_1 _2181__120 (.LO(net120));
 sky130_fd_sc_hd__conb_1 _2182__121 (.LO(net121));
 sky130_fd_sc_hd__conb_1 _2183__122 (.LO(net122));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__ebufn_8 _2076_ (.A(net26),
    .TE_B(_0751_),
    .Z(la1_data_out[0]));
 sky130_fd_sc_hd__ebufn_8 _2077_ (.A(net27),
    .TE_B(_0752_),
    .Z(la1_data_out[1]));
 sky130_fd_sc_hd__ebufn_8 _2078_ (.A(net28),
    .TE_B(_0753_),
    .Z(la1_data_out[2]));
 sky130_fd_sc_hd__ebufn_8 _2079_ (.A(net29),
    .TE_B(_0754_),
    .Z(la1_data_out[3]));
 sky130_fd_sc_hd__ebufn_8 _2080_ (.A(net30),
    .TE_B(_0755_),
    .Z(la1_data_out[4]));
 sky130_fd_sc_hd__ebufn_8 _2081_ (.A(net31),
    .TE_B(_0756_),
    .Z(la1_data_out[5]));
 sky130_fd_sc_hd__ebufn_8 _2082_ (.A(net32),
    .TE_B(_0757_),
    .Z(la1_data_out[6]));
 sky130_fd_sc_hd__ebufn_8 _2083_ (.A(\gps_channel0.prompt_q ),
    .TE_B(_0758_),
    .Z(la1_data_out[7]));
 sky130_fd_sc_hd__ebufn_8 _2084_ (.A(\gps_channel0.lo_nco.accumulator[28] ),
    .TE_B(_0759_),
    .Z(la1_data_out[8]));
 sky130_fd_sc_hd__ebufn_8 _2085_ (.A(\gps_channel0.lo_nco.accumulator[29] ),
    .TE_B(_0760_),
    .Z(la1_data_out[9]));
 sky130_fd_sc_hd__ebufn_8 _2086_ (.A(\gps_channel0.lo_nco.accumulator[30] ),
    .TE_B(_0761_),
    .Z(la1_data_out[10]));
 sky130_fd_sc_hd__ebufn_8 _2087_ (.A(\gps_channel0.lo_i ),
    .TE_B(_0762_),
    .Z(la1_data_out[11]));
 sky130_fd_sc_hd__ebufn_8 _2088_ (.A(\gps_channel0.ca_nco.accumulator[28] ),
    .TE_B(_0763_),
    .Z(la1_data_out[12]));
 sky130_fd_sc_hd__ebufn_8 _2089_ (.A(\gps_channel0.ca_nco.accumulator[29] ),
    .TE_B(_0764_),
    .Z(la1_data_out[13]));
 sky130_fd_sc_hd__ebufn_8 _2090_ (.A(\gps_channel0.ca_nco.accumulator[30] ),
    .TE_B(_0765_),
    .Z(la1_data_out[14]));
 sky130_fd_sc_hd__ebufn_8 _2091_ (.A(\gps_channel0.ca_nco.accumulator[31] ),
    .TE_B(_0766_),
    .Z(la1_data_out[15]));
 sky130_fd_sc_hd__ebufn_8 _2092_ (.A(net33),
    .TE_B(_0767_),
    .Z(la1_data_out[16]));
 sky130_fd_sc_hd__ebufn_8 _2093_ (.A(net34),
    .TE_B(_0768_),
    .Z(la1_data_out[17]));
 sky130_fd_sc_hd__ebufn_8 _2094_ (.A(net35),
    .TE_B(_0769_),
    .Z(la1_data_out[18]));
 sky130_fd_sc_hd__ebufn_8 _2095_ (.A(net36),
    .TE_B(_0770_),
    .Z(la1_data_out[19]));
 sky130_fd_sc_hd__ebufn_8 _2096_ (.A(net37),
    .TE_B(_0771_),
    .Z(la1_data_out[20]));
 sky130_fd_sc_hd__ebufn_8 _2097_ (.A(net38),
    .TE_B(_0772_),
    .Z(la1_data_out[21]));
 sky130_fd_sc_hd__ebufn_8 _2098_ (.A(net39),
    .TE_B(_0773_),
    .Z(la1_data_out[22]));
 sky130_fd_sc_hd__ebufn_8 _2099_ (.A(net40),
    .TE_B(_0774_),
    .Z(la1_data_out[23]));
 sky130_fd_sc_hd__ebufn_8 _2100_ (.A(net41),
    .TE_B(_0775_),
    .Z(la1_data_out[24]));
 sky130_fd_sc_hd__ebufn_8 _2101_ (.A(net42),
    .TE_B(_0776_),
    .Z(la1_data_out[25]));
 sky130_fd_sc_hd__ebufn_8 _2102_ (.A(net43),
    .TE_B(_0777_),
    .Z(la1_data_out[26]));
 sky130_fd_sc_hd__ebufn_8 _2103_ (.A(net44),
    .TE_B(_0778_),
    .Z(la1_data_out[27]));
 sky130_fd_sc_hd__ebufn_8 _2104_ (.A(net45),
    .TE_B(_0779_),
    .Z(la1_data_out[28]));
 sky130_fd_sc_hd__ebufn_8 _2105_ (.A(net46),
    .TE_B(_0780_),
    .Z(la1_data_out[29]));
 sky130_fd_sc_hd__ebufn_8 _2106_ (.A(net47),
    .TE_B(_0781_),
    .Z(la1_data_out[30]));
 sky130_fd_sc_hd__ebufn_8 _2107_ (.A(net48),
    .TE_B(_0782_),
    .Z(la1_data_out[31]));
 sky130_fd_sc_hd__ebufn_8 _2108_ (.A(net49),
    .TE_B(_0783_),
    .Z(io_out[0]));
 sky130_fd_sc_hd__ebufn_8 _2109_ (.A(net50),
    .TE_B(_0784_),
    .Z(io_out[1]));
 sky130_fd_sc_hd__ebufn_8 _2110_ (.A(net51),
    .TE_B(_0785_),
    .Z(io_out[2]));
 sky130_fd_sc_hd__ebufn_8 _2111_ (.A(net52),
    .TE_B(_0786_),
    .Z(io_out[3]));
 sky130_fd_sc_hd__ebufn_8 _2112_ (.A(net53),
    .TE_B(_0787_),
    .Z(io_out[4]));
 sky130_fd_sc_hd__ebufn_8 _2113_ (.A(net54),
    .TE_B(_0788_),
    .Z(io_out[5]));
 sky130_fd_sc_hd__ebufn_8 _2114_ (.A(net55),
    .TE_B(_0789_),
    .Z(io_out[6]));
 sky130_fd_sc_hd__ebufn_8 _2115_ (.A(net56),
    .TE_B(_0790_),
    .Z(io_out[7]));
 sky130_fd_sc_hd__ebufn_8 _2116_ (.A(net57),
    .TE_B(_0791_),
    .Z(io_out[8]));
 sky130_fd_sc_hd__ebufn_8 _2117_ (.A(net58),
    .TE_B(_0792_),
    .Z(io_out[9]));
 sky130_fd_sc_hd__ebufn_8 _2118_ (.A(net59),
    .TE_B(_0793_),
    .Z(io_out[10]));
 sky130_fd_sc_hd__ebufn_8 _2119_ (.A(net60),
    .TE_B(_0794_),
    .Z(io_out[11]));
 sky130_fd_sc_hd__ebufn_8 _2120_ (.A(net61),
    .TE_B(_0795_),
    .Z(io_out[12]));
 sky130_fd_sc_hd__ebufn_8 _2121_ (.A(net62),
    .TE_B(_0796_),
    .Z(io_out[13]));
 sky130_fd_sc_hd__ebufn_8 _2122_ (.A(net63),
    .TE_B(_0797_),
    .Z(io_out[14]));
 sky130_fd_sc_hd__ebufn_8 _2123_ (.A(net64),
    .TE_B(_0798_),
    .Z(io_out[15]));
 sky130_fd_sc_hd__ebufn_8 _2124_ (.A(net65),
    .TE_B(_0799_),
    .Z(io_out[16]));
 sky130_fd_sc_hd__ebufn_8 _2125_ (.A(net66),
    .TE_B(_0800_),
    .Z(io_out[17]));
 sky130_fd_sc_hd__ebufn_8 _2126_ (.A(net67),
    .TE_B(_0801_),
    .Z(io_out[18]));
 sky130_fd_sc_hd__ebufn_8 _2127_ (.A(\gps_channel0.lo_i ),
    .TE_B(_0802_),
    .Z(io_out[19]));
 sky130_fd_sc_hd__ebufn_8 _2128_ (.A(net68),
    .TE_B(_0803_),
    .Z(io_out[20]));
 sky130_fd_sc_hd__ebufn_8 _2129_ (.A(\gps_channel0.prompt_i ),
    .TE_B(_0804_),
    .Z(io_out[21]));
 sky130_fd_sc_hd__ebufn_8 _2130_ (.A(net69),
    .TE_B(_0805_),
    .Z(io_out[22]));
 sky130_fd_sc_hd__ebufn_8 _2131_ (.A(net70),
    .TE_B(_0806_),
    .Z(io_out[23]));
 sky130_fd_sc_hd__ebufn_8 _2132_ (.A(net71),
    .TE_B(_0807_),
    .Z(io_out[24]));
 sky130_fd_sc_hd__ebufn_8 _2133_ (.A(net72),
    .TE_B(_0808_),
    .Z(io_out[25]));
 sky130_fd_sc_hd__ebufn_8 _2134_ (.A(net73),
    .TE_B(_0809_),
    .Z(io_out[26]));
 sky130_fd_sc_hd__ebufn_8 _2135_ (.A(net74),
    .TE_B(_0810_),
    .Z(io_out[27]));
 sky130_fd_sc_hd__ebufn_8 _2136_ (.A(net75),
    .TE_B(_0811_),
    .Z(io_out[28]));
 sky130_fd_sc_hd__ebufn_8 _2137_ (.A(net76),
    .TE_B(_0812_),
    .Z(io_out[29]));
 sky130_fd_sc_hd__ebufn_8 _2138_ (.A(net77),
    .TE_B(_0813_),
    .Z(io_out[30]));
 sky130_fd_sc_hd__ebufn_8 _2139_ (.A(net78),
    .TE_B(_0814_),
    .Z(io_out[31]));
 sky130_fd_sc_hd__ebufn_8 _2140_ (.A(net79),
    .TE_B(_0815_),
    .Z(io_out[32]));
 sky130_fd_sc_hd__ebufn_8 _2141_ (.A(net80),
    .TE_B(_0816_),
    .Z(io_out[33]));
 sky130_fd_sc_hd__ebufn_8 _2142_ (.A(net81),
    .TE_B(_0817_),
    .Z(io_out[34]));
 sky130_fd_sc_hd__ebufn_8 _2143_ (.A(net82),
    .TE_B(_0818_),
    .Z(io_out[35]));
 sky130_fd_sc_hd__ebufn_8 _2144_ (.A(net83),
    .TE_B(_0819_),
    .Z(io_out[36]));
 sky130_fd_sc_hd__ebufn_8 _2145_ (.A(net84),
    .TE_B(_0820_),
    .Z(io_out[37]));
 sky130_fd_sc_hd__ebufn_8 _2146_ (.A(net85),
    .TE_B(_0821_),
    .Z(io_oeb[0]));
 sky130_fd_sc_hd__ebufn_8 _2147_ (.A(net86),
    .TE_B(_0822_),
    .Z(io_oeb[1]));
 sky130_fd_sc_hd__ebufn_8 _2148_ (.A(net87),
    .TE_B(_0823_),
    .Z(io_oeb[2]));
 sky130_fd_sc_hd__ebufn_8 _2149_ (.A(net88),
    .TE_B(_0824_),
    .Z(io_oeb[3]));
 sky130_fd_sc_hd__ebufn_8 _2150_ (.A(net89),
    .TE_B(_0825_),
    .Z(io_oeb[4]));
 sky130_fd_sc_hd__ebufn_8 _2151_ (.A(net90),
    .TE_B(_0826_),
    .Z(io_oeb[5]));
 sky130_fd_sc_hd__ebufn_8 _2152_ (.A(net91),
    .TE_B(_0827_),
    .Z(io_oeb[6]));
 sky130_fd_sc_hd__ebufn_8 _2153_ (.A(net92),
    .TE_B(_0828_),
    .Z(io_oeb[7]));
 sky130_fd_sc_hd__ebufn_8 _2154_ (.A(net93),
    .TE_B(_0829_),
    .Z(io_oeb[8]));
 sky130_fd_sc_hd__ebufn_8 _2155_ (.A(net94),
    .TE_B(_0830_),
    .Z(io_oeb[9]));
 sky130_fd_sc_hd__ebufn_8 _2156_ (.A(net95),
    .TE_B(_0831_),
    .Z(io_oeb[10]));
 sky130_fd_sc_hd__ebufn_8 _2157_ (.A(net96),
    .TE_B(_0832_),
    .Z(io_oeb[11]));
 sky130_fd_sc_hd__ebufn_8 _2158_ (.A(net97),
    .TE_B(_0833_),
    .Z(io_oeb[12]));
 sky130_fd_sc_hd__ebufn_8 _2159_ (.A(net98),
    .TE_B(_0834_),
    .Z(io_oeb[13]));
 sky130_fd_sc_hd__ebufn_8 _2160_ (.A(net99),
    .TE_B(_0835_),
    .Z(io_oeb[14]));
 sky130_fd_sc_hd__ebufn_8 _2161_ (.A(net100),
    .TE_B(_0836_),
    .Z(io_oeb[15]));
 sky130_fd_sc_hd__ebufn_8 _2162_ (.A(net101),
    .TE_B(_0837_),
    .Z(io_oeb[16]));
 sky130_fd_sc_hd__ebufn_8 _2163_ (.A(net102),
    .TE_B(_0838_),
    .Z(io_oeb[17]));
 sky130_fd_sc_hd__ebufn_8 _2164_ (.A(net103),
    .TE_B(_0839_),
    .Z(io_oeb[18]));
 sky130_fd_sc_hd__ebufn_8 _2165_ (.A(net104),
    .TE_B(_0840_),
    .Z(io_oeb[19]));
 sky130_fd_sc_hd__ebufn_8 _2166_ (.A(net105),
    .TE_B(_0841_),
    .Z(io_oeb[20]));
 sky130_fd_sc_hd__ebufn_8 _2167_ (.A(net106),
    .TE_B(_0842_),
    .Z(io_oeb[21]));
 sky130_fd_sc_hd__ebufn_8 _2168_ (.A(net107),
    .TE_B(_0843_),
    .Z(io_oeb[22]));
 sky130_fd_sc_hd__ebufn_8 _2169_ (.A(net108),
    .TE_B(_0844_),
    .Z(io_oeb[23]));
 sky130_fd_sc_hd__ebufn_8 _2170_ (.A(net109),
    .TE_B(_0845_),
    .Z(io_oeb[24]));
 sky130_fd_sc_hd__ebufn_8 _2171_ (.A(net110),
    .TE_B(_0846_),
    .Z(io_oeb[25]));
 sky130_fd_sc_hd__ebufn_8 _2172_ (.A(net111),
    .TE_B(_0847_),
    .Z(io_oeb[26]));
 sky130_fd_sc_hd__ebufn_8 _2173_ (.A(net112),
    .TE_B(_0848_),
    .Z(io_oeb[27]));
 sky130_fd_sc_hd__ebufn_8 _2174_ (.A(net113),
    .TE_B(_0849_),
    .Z(io_oeb[28]));
 sky130_fd_sc_hd__ebufn_8 _2175_ (.A(net114),
    .TE_B(_0850_),
    .Z(io_oeb[29]));
 sky130_fd_sc_hd__ebufn_8 _2176_ (.A(net115),
    .TE_B(_0851_),
    .Z(io_oeb[30]));
 sky130_fd_sc_hd__ebufn_8 _2177_ (.A(net116),
    .TE_B(_0852_),
    .Z(io_oeb[31]));
 sky130_fd_sc_hd__ebufn_8 _2178_ (.A(net117),
    .TE_B(_0853_),
    .Z(io_oeb[32]));
 sky130_fd_sc_hd__ebufn_8 _2179_ (.A(net118),
    .TE_B(_0854_),
    .Z(io_oeb[33]));
 sky130_fd_sc_hd__ebufn_8 _2180_ (.A(net119),
    .TE_B(_0855_),
    .Z(io_oeb[34]));
 sky130_fd_sc_hd__ebufn_8 _2181_ (.A(net120),
    .TE_B(_0856_),
    .Z(io_oeb[35]));
 sky130_fd_sc_hd__ebufn_8 _2182_ (.A(net121),
    .TE_B(_0857_),
    .Z(io_oeb[36]));
 sky130_fd_sc_hd__ebufn_8 _2183_ (.A(net122),
    .TE_B(_0858_),
    .Z(io_oeb[37]));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(active),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(io_in[23]),
    .X(net2));
 sky130_fd_sc_hd__buf_4 input3 (.A(la1_data_in[0]),
    .X(net3));
 sky130_fd_sc_hd__buf_2 input4 (.A(la1_data_in[16]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input5 (.A(la1_data_in[17]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(la1_data_in[18]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(la1_data_in[19]),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input8 (.A(la1_data_in[1]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(la1_data_in[20]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 input10 (.A(la1_data_in[21]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(la1_data_in[22]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 input12 (.A(la1_data_in[23]),
    .X(net12));
 sky130_fd_sc_hd__buf_2 input13 (.A(la1_data_in[24]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(la1_data_in[25]),
    .X(net14));
 sky130_fd_sc_hd__buf_2 input15 (.A(la1_data_in[26]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(la1_data_in[27]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(la1_data_in[28]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 input18 (.A(la1_data_in[29]),
    .X(net18));
 sky130_fd_sc_hd__buf_2 input19 (.A(la1_data_in[2]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input20 (.A(la1_data_in[30]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(la1_data_in[31]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(la1_data_in[3]),
    .X(net22));
 sky130_fd_sc_hd__buf_2 input23 (.A(la1_data_in[4]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(la1_data_in[5]),
    .X(net24));
 sky130_fd_sc_hd__buf_2 input25 (.A(la1_data_in[6]),
    .X(net25));
 sky130_fd_sc_hd__conb_1 _2076__26 (.LO(net26));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_4_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_5_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_6_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_7_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_8_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_9_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_10_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_11_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_12_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_13_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_14_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_15_0_wb_clk_i));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_514 ();
endmodule

