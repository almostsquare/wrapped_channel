magic
tech sky130B
magscale 1 2
timestamp 1671932820
<< viali >>
rect 17693 47141 17727 47175
rect 32505 47141 32539 47175
rect 42809 47141 42843 47175
rect 3433 47073 3467 47107
rect 9137 47073 9171 47107
rect 14749 47073 14783 47107
rect 47225 47073 47259 47107
rect 2145 47005 2179 47039
rect 2697 47005 2731 47039
rect 3985 47005 4019 47039
rect 5457 47005 5491 47039
rect 6561 47005 6595 47039
rect 7389 47005 7423 47039
rect 9413 47005 9447 47039
rect 12725 47005 12759 47039
rect 13737 47005 13771 47039
rect 14289 47005 14323 47039
rect 17509 47005 17543 47039
rect 19533 47005 19567 47039
rect 22937 47005 22971 47039
rect 24685 47005 24719 47039
rect 25697 47005 25731 47039
rect 30021 47005 30055 47039
rect 32321 47005 32355 47039
rect 33241 47005 33275 47039
rect 38577 47005 38611 47039
rect 40233 47005 40267 47039
rect 41429 47005 41463 47039
rect 42625 47005 42659 47039
rect 45385 47005 45419 47039
rect 47961 47005 47995 47039
rect 4813 46937 4847 46971
rect 6653 46937 6687 46971
rect 14473 46937 14507 46971
rect 19717 46937 19751 46971
rect 25053 46937 25087 46971
rect 45569 46937 45603 46971
rect 5549 46869 5583 46903
rect 48053 46869 48087 46903
rect 6009 46597 6043 46631
rect 47225 46597 47259 46631
rect 4169 46529 4203 46563
rect 11989 46529 12023 46563
rect 22477 46529 22511 46563
rect 24777 46529 24811 46563
rect 32873 46529 32907 46563
rect 39773 46529 39807 46563
rect 42625 46529 42659 46563
rect 47777 46529 47811 46563
rect 1869 46461 1903 46495
rect 2053 46461 2087 46495
rect 2329 46461 2363 46495
rect 4353 46461 4387 46495
rect 12173 46461 12207 46495
rect 12909 46461 12943 46495
rect 14289 46461 14323 46495
rect 14473 46461 14507 46495
rect 14841 46461 14875 46495
rect 22661 46461 22695 46495
rect 23213 46461 23247 46495
rect 24961 46461 24995 46495
rect 25789 46461 25823 46495
rect 28549 46461 28583 46495
rect 29009 46461 29043 46495
rect 29193 46461 29227 46495
rect 29653 46461 29687 46495
rect 33057 46461 33091 46495
rect 33517 46461 33551 46495
rect 36461 46461 36495 46495
rect 37473 46461 37507 46495
rect 37657 46461 37691 46495
rect 37933 46461 37967 46495
rect 39957 46461 39991 46495
rect 40233 46461 40267 46495
rect 42809 46461 42843 46495
rect 43085 46461 43119 46495
rect 45385 46461 45419 46495
rect 45569 46461 45603 46495
rect 7389 46393 7423 46427
rect 6745 46325 6779 46359
rect 8033 46325 8067 46359
rect 17049 46325 17083 46359
rect 35725 46325 35759 46359
rect 47869 46325 47903 46359
rect 7665 46121 7699 46155
rect 12541 46121 12575 46155
rect 13645 46121 13679 46155
rect 14473 46121 14507 46155
rect 22753 46121 22787 46155
rect 29101 46121 29135 46155
rect 33149 46121 33183 46155
rect 38485 46121 38519 46155
rect 45385 46121 45419 46155
rect 45937 46121 45971 46155
rect 1593 45985 1627 46019
rect 2789 45985 2823 46019
rect 5273 45985 5307 46019
rect 5457 45985 5491 46019
rect 5825 45985 5859 46019
rect 15025 45985 15059 46019
rect 15485 45985 15519 46019
rect 35449 45985 35483 46019
rect 36093 45985 36127 46019
rect 40049 45985 40083 46019
rect 40601 45985 40635 46019
rect 46673 45985 46707 46019
rect 48237 45985 48271 46019
rect 4077 45917 4111 45951
rect 7573 45917 7607 45951
rect 12449 45917 12483 45951
rect 13553 45917 13587 45951
rect 14381 45917 14415 45951
rect 22661 45917 22695 45951
rect 24041 45917 24075 45951
rect 24685 45917 24719 45951
rect 29009 45917 29043 45951
rect 29745 45917 29779 45951
rect 33057 45917 33091 45951
rect 38393 45917 38427 45951
rect 45845 45917 45879 45951
rect 46489 45917 46523 45951
rect 1777 45849 1811 45883
rect 4629 45849 4663 45883
rect 15209 45849 15243 45883
rect 24869 45849 24903 45883
rect 26525 45849 26559 45883
rect 29929 45849 29963 45883
rect 31585 45849 31619 45883
rect 35633 45849 35667 45883
rect 40233 45849 40267 45883
rect 15301 45577 15335 45611
rect 24869 45577 24903 45611
rect 25513 45577 25547 45611
rect 29837 45577 29871 45611
rect 35541 45577 35575 45611
rect 40049 45577 40083 45611
rect 2329 45509 2363 45543
rect 6653 45509 6687 45543
rect 7297 45509 7331 45543
rect 36369 45509 36403 45543
rect 41429 45509 41463 45543
rect 47041 45509 47075 45543
rect 4813 45441 4847 45475
rect 6561 45441 6595 45475
rect 7205 45441 7239 45475
rect 14473 45441 14507 45475
rect 15209 45441 15243 45475
rect 24777 45441 24811 45475
rect 25421 45441 25455 45475
rect 29745 45441 29779 45475
rect 35449 45441 35483 45475
rect 36277 45441 36311 45475
rect 39957 45441 39991 45475
rect 41337 45441 41371 45475
rect 45845 45441 45879 45475
rect 46489 45441 46523 45475
rect 46949 45441 46983 45475
rect 2145 45373 2179 45407
rect 2973 45373 3007 45407
rect 5457 45373 5491 45407
rect 10701 45237 10735 45271
rect 47961 45237 47995 45271
rect 6837 44897 6871 44931
rect 10517 44897 10551 44931
rect 11069 44897 11103 44931
rect 40601 44897 40635 44931
rect 46489 44897 46523 44931
rect 48237 44897 48271 44931
rect 1593 44829 1627 44863
rect 2605 44829 2639 44863
rect 3985 44829 4019 44863
rect 6193 44829 6227 44863
rect 40049 44829 40083 44863
rect 3249 44761 3283 44795
rect 10701 44761 10735 44795
rect 46673 44761 46707 44795
rect 1777 44693 1811 44727
rect 5273 44693 5307 44727
rect 10609 44489 10643 44523
rect 47869 44489 47903 44523
rect 4905 44353 4939 44387
rect 10517 44353 10551 44387
rect 20361 44353 20395 44387
rect 47777 44353 47811 44387
rect 2053 44285 2087 44319
rect 2237 44285 2271 44319
rect 2789 44285 2823 44319
rect 5089 44285 5123 44319
rect 20453 44149 20487 44183
rect 29745 43877 29779 43911
rect 2789 43809 2823 43843
rect 4997 43809 5031 43843
rect 20545 43809 20579 43843
rect 22201 43809 22235 43843
rect 1593 43741 1627 43775
rect 4629 43741 4663 43775
rect 20361 43741 20395 43775
rect 30021 43741 30055 43775
rect 30481 43741 30515 43775
rect 30665 43741 30699 43775
rect 1777 43673 1811 43707
rect 29745 43673 29779 43707
rect 29929 43605 29963 43639
rect 30665 43605 30699 43639
rect 2421 43401 2455 43435
rect 19073 43333 19107 43367
rect 25697 43333 25731 43367
rect 30941 43333 30975 43367
rect 1869 43265 1903 43299
rect 2329 43265 2363 43299
rect 3709 43265 3743 43299
rect 25513 43265 25547 43299
rect 25789 43265 25823 43299
rect 25881 43265 25915 43299
rect 29009 43265 29043 43299
rect 30021 43265 30055 43299
rect 30113 43265 30147 43299
rect 31125 43265 31159 43299
rect 32377 43265 32411 43299
rect 32505 43265 32539 43299
rect 32597 43265 32631 43299
rect 33701 43265 33735 43299
rect 34529 43265 34563 43299
rect 47777 43265 47811 43299
rect 3893 43197 3927 43231
rect 17233 43197 17267 43231
rect 17417 43197 17451 43231
rect 29101 43197 29135 43231
rect 30205 43197 30239 43231
rect 30297 43197 30331 43231
rect 33609 43197 33643 43231
rect 34069 43197 34103 43231
rect 34805 43197 34839 43231
rect 29377 43129 29411 43163
rect 34621 43129 34655 43163
rect 26065 43061 26099 43095
rect 29837 43061 29871 43095
rect 31309 43061 31343 43095
rect 32781 43061 32815 43095
rect 34713 43061 34747 43095
rect 47225 43061 47259 43095
rect 47869 43061 47903 43095
rect 17417 42857 17451 42891
rect 27169 42857 27203 42891
rect 22201 42789 22235 42823
rect 29193 42789 29227 42823
rect 32597 42789 32631 42823
rect 33885 42789 33919 42823
rect 2329 42721 2363 42755
rect 3065 42721 3099 42755
rect 5549 42721 5583 42755
rect 23305 42721 23339 42755
rect 27813 42721 27847 42755
rect 29929 42721 29963 42755
rect 30389 42721 30423 42755
rect 34069 42721 34103 42755
rect 46489 42721 46523 42755
rect 48237 42721 48271 42755
rect 1777 42653 1811 42687
rect 2237 42653 2271 42687
rect 4905 42653 4939 42687
rect 17325 42653 17359 42687
rect 19717 42653 19751 42687
rect 20821 42653 20855 42687
rect 22845 42653 22879 42687
rect 23147 42653 23181 42687
rect 25237 42653 25271 42687
rect 27077 42653 27111 42687
rect 27261 42653 27295 42687
rect 30021 42653 30055 42687
rect 31033 42653 31067 42687
rect 31493 42653 31527 42687
rect 31953 42653 31987 42687
rect 32321 42653 32355 42687
rect 32413 42653 32447 42687
rect 33057 42653 33091 42687
rect 33793 42653 33827 42687
rect 35081 42653 35115 42687
rect 5089 42585 5123 42619
rect 19441 42585 19475 42619
rect 21088 42585 21122 42619
rect 22661 42585 22695 42619
rect 22937 42585 22971 42619
rect 23029 42585 23063 42619
rect 25504 42585 25538 42619
rect 28080 42585 28114 42619
rect 30297 42585 30331 42619
rect 31125 42585 31159 42619
rect 31217 42585 31251 42619
rect 31355 42585 31389 42619
rect 34069 42585 34103 42619
rect 35326 42585 35360 42619
rect 46673 42585 46707 42619
rect 1593 42517 1627 42551
rect 19539 42517 19573 42551
rect 19625 42517 19659 42551
rect 26617 42517 26651 42551
rect 29745 42517 29779 42551
rect 30849 42517 30883 42551
rect 33241 42517 33275 42551
rect 36461 42517 36495 42551
rect 5089 42313 5123 42347
rect 17417 42313 17451 42347
rect 20177 42313 20211 42347
rect 23305 42313 23339 42347
rect 24317 42313 24351 42347
rect 25145 42313 25179 42347
rect 30665 42313 30699 42347
rect 32689 42313 32723 42347
rect 34437 42313 34471 42347
rect 29552 42245 29586 42279
rect 31493 42245 31527 42279
rect 32597 42245 32631 42279
rect 33977 42245 34011 42279
rect 34734 42245 34768 42279
rect 4997 42177 5031 42211
rect 15945 42177 15979 42211
rect 17141 42177 17175 42211
rect 17233 42177 17267 42211
rect 19064 42177 19098 42211
rect 22477 42177 22511 42211
rect 23489 42177 23523 42211
rect 23673 42177 23707 42211
rect 23765 42177 23799 42211
rect 24225 42177 24259 42211
rect 24409 42177 24443 42211
rect 24501 42177 24535 42211
rect 25329 42177 25363 42211
rect 26249 42177 26283 42211
rect 27169 42177 27203 42211
rect 29285 42177 29319 42211
rect 31125 42177 31159 42211
rect 31309 42177 31343 42211
rect 32505 42177 32539 42211
rect 33793 42177 33827 42211
rect 34621 42177 34655 42211
rect 34818 42177 34852 42211
rect 34923 42177 34957 42211
rect 35081 42177 35115 42211
rect 35541 42177 35575 42211
rect 35725 42177 35759 42211
rect 47777 42177 47811 42211
rect 16037 42109 16071 42143
rect 16129 42109 16163 42143
rect 18797 42109 18831 42143
rect 22569 42109 22603 42143
rect 25605 42109 25639 42143
rect 26157 42109 26191 42143
rect 33609 42109 33643 42143
rect 22845 42041 22879 42075
rect 26617 42041 26651 42075
rect 32321 42041 32355 42075
rect 15577 41973 15611 42007
rect 25513 41973 25547 42007
rect 27261 41973 27295 42007
rect 32873 41973 32907 42007
rect 35541 41973 35575 42007
rect 47225 41973 47259 42007
rect 47869 41973 47903 42007
rect 16865 41769 16899 41803
rect 17509 41769 17543 41803
rect 17693 41769 17727 41803
rect 19441 41769 19475 41803
rect 21925 41769 21959 41803
rect 31125 41769 31159 41803
rect 31217 41769 31251 41803
rect 33057 41769 33091 41803
rect 35081 41769 35115 41803
rect 23305 41701 23339 41735
rect 25605 41701 25639 41735
rect 31309 41701 31343 41735
rect 35265 41701 35299 41735
rect 15485 41633 15519 41667
rect 19625 41633 19659 41667
rect 20085 41633 20119 41667
rect 20821 41633 20855 41667
rect 21005 41633 21039 41667
rect 22109 41633 22143 41667
rect 24961 41633 24995 41667
rect 33701 41633 33735 41667
rect 46489 41633 46523 41667
rect 46673 41633 46707 41667
rect 48237 41633 48271 41667
rect 2237 41565 2271 41599
rect 14933 41565 14967 41599
rect 19717 41565 19751 41599
rect 19993 41565 20027 41599
rect 20729 41565 20763 41599
rect 20913 41565 20947 41599
rect 21833 41565 21867 41599
rect 23121 41565 23155 41599
rect 23213 41565 23247 41599
rect 23397 41565 23431 41599
rect 23765 41565 23799 41599
rect 25605 41565 25639 41599
rect 25789 41565 25823 41599
rect 26801 41565 26835 41599
rect 26893 41565 26927 41599
rect 27077 41565 27111 41599
rect 27169 41565 27203 41599
rect 31033 41565 31067 41599
rect 31493 41565 31527 41599
rect 32965 41565 32999 41599
rect 33149 41565 33183 41599
rect 33609 41565 33643 41599
rect 33793 41565 33827 41599
rect 34897 41565 34931 41599
rect 35081 41565 35115 41599
rect 46029 41565 46063 41599
rect 15752 41497 15786 41531
rect 17325 41497 17359 41531
rect 22109 41497 22143 41531
rect 24593 41497 24627 41531
rect 24777 41497 24811 41531
rect 25973 41497 26007 41531
rect 14749 41429 14783 41463
rect 17525 41429 17559 41463
rect 20545 41429 20579 41463
rect 26617 41429 26651 41463
rect 30757 41429 30791 41463
rect 15485 41225 15519 41259
rect 19533 41225 19567 41259
rect 23581 41225 23615 41259
rect 27169 41225 27203 41259
rect 33885 41225 33919 41259
rect 14372 41157 14406 41191
rect 19257 41157 19291 41191
rect 22385 41157 22419 41191
rect 23213 41157 23247 41191
rect 24133 41157 24167 41191
rect 27721 41157 27755 41191
rect 35234 41157 35268 41191
rect 2053 41089 2087 41123
rect 16037 41089 16071 41123
rect 16129 41089 16163 41123
rect 16865 41089 16899 41123
rect 17049 41089 17083 41123
rect 17233 41089 17267 41123
rect 17325 41089 17359 41123
rect 19441 41089 19475 41123
rect 19625 41089 19659 41123
rect 20361 41089 20395 41123
rect 22569 41089 22603 41123
rect 23397 41089 23431 41123
rect 23673 41089 23707 41123
rect 24317 41089 24351 41123
rect 24409 41089 24443 41123
rect 27445 41089 27479 41123
rect 29377 41089 29411 41123
rect 33241 41089 33275 41123
rect 34161 41089 34195 41123
rect 45385 41089 45419 41123
rect 2237 41021 2271 41055
rect 2789 41021 2823 41055
rect 14105 41021 14139 41055
rect 27353 41021 27387 41055
rect 27813 41021 27847 41055
rect 33057 41021 33091 41055
rect 33425 41021 33459 41055
rect 34069 41021 34103 41055
rect 34437 41021 34471 41055
rect 34529 41021 34563 41055
rect 34989 41021 35023 41055
rect 45569 41021 45603 41055
rect 46949 41021 46983 41055
rect 24225 40953 24259 40987
rect 16313 40885 16347 40919
rect 19809 40885 19843 40919
rect 20453 40885 20487 40919
rect 22753 40885 22787 40919
rect 29469 40885 29503 40919
rect 36369 40885 36403 40919
rect 47961 40885 47995 40919
rect 2329 40681 2363 40715
rect 15945 40681 15979 40715
rect 17233 40681 17267 40715
rect 22017 40681 22051 40715
rect 23673 40681 23707 40715
rect 33885 40681 33919 40715
rect 45937 40681 45971 40715
rect 30941 40613 30975 40647
rect 33793 40613 33827 40647
rect 17049 40545 17083 40579
rect 20085 40545 20119 40579
rect 25789 40545 25823 40579
rect 33977 40545 34011 40579
rect 46489 40545 46523 40579
rect 2237 40477 2271 40511
rect 16129 40477 16163 40511
rect 16865 40477 16899 40511
rect 17233 40477 17267 40511
rect 19566 40477 19600 40511
rect 19993 40477 20027 40511
rect 20637 40477 20671 40511
rect 22661 40477 22695 40511
rect 22963 40477 22997 40511
rect 23121 40477 23155 40511
rect 23581 40477 23615 40511
rect 23765 40477 23799 40511
rect 24685 40477 24719 40511
rect 25697 40477 25731 40511
rect 26525 40477 26559 40511
rect 26709 40477 26743 40511
rect 27169 40477 27203 40511
rect 30941 40477 30975 40511
rect 31217 40477 31251 40511
rect 32229 40477 32263 40511
rect 33701 40477 33735 40511
rect 45845 40477 45879 40511
rect 16957 40409 16991 40443
rect 20904 40409 20938 40443
rect 22477 40409 22511 40443
rect 22753 40409 22787 40443
rect 22845 40409 22879 40443
rect 25053 40409 25087 40443
rect 27436 40409 27470 40443
rect 46673 40409 46707 40443
rect 48329 40409 48363 40443
rect 19441 40341 19475 40375
rect 19625 40341 19659 40375
rect 26065 40341 26099 40375
rect 26709 40341 26743 40375
rect 28549 40341 28583 40375
rect 31125 40341 31159 40375
rect 32321 40341 32355 40375
rect 19809 40137 19843 40171
rect 27721 40137 27755 40171
rect 32597 40137 32631 40171
rect 27353 40069 27387 40103
rect 27445 40069 27479 40103
rect 30481 40069 30515 40103
rect 32413 40069 32447 40103
rect 18696 40001 18730 40035
rect 22569 40001 22603 40035
rect 22753 40001 22787 40035
rect 27169 40001 27203 40035
rect 27537 40001 27571 40035
rect 28273 40001 28307 40035
rect 30665 40001 30699 40035
rect 32320 40023 32354 40057
rect 32689 40001 32723 40035
rect 47041 40001 47075 40035
rect 47133 40001 47167 40035
rect 18429 39933 18463 39967
rect 22661 39933 22695 39967
rect 32505 39933 32539 39967
rect 28365 39797 28399 39831
rect 30849 39797 30883 39831
rect 47961 39797 47995 39831
rect 26709 39593 26743 39627
rect 30849 39593 30883 39627
rect 32045 39593 32079 39627
rect 27077 39525 27111 39559
rect 27997 39525 28031 39559
rect 33609 39525 33643 39559
rect 14289 39457 14323 39491
rect 20177 39457 20211 39491
rect 27169 39457 27203 39491
rect 27629 39457 27663 39491
rect 29929 39457 29963 39491
rect 33333 39457 33367 39491
rect 46489 39457 46523 39491
rect 48237 39457 48271 39491
rect 26893 39389 26927 39423
rect 27813 39389 27847 39423
rect 29837 39389 29871 39423
rect 30021 39389 30055 39423
rect 30665 39389 30699 39423
rect 30941 39389 30975 39423
rect 31401 39389 31435 39423
rect 31585 39389 31619 39423
rect 32045 39389 32079 39423
rect 32137 39389 32171 39423
rect 33241 39389 33275 39423
rect 14534 39321 14568 39355
rect 19441 39321 19475 39355
rect 46673 39321 46707 39355
rect 15669 39253 15703 39287
rect 30481 39253 30515 39287
rect 31493 39253 31527 39287
rect 32413 39253 32447 39287
rect 13921 39049 13955 39083
rect 19809 39049 19843 39083
rect 20453 39049 20487 39083
rect 30389 39049 30423 39083
rect 31033 39049 31067 39083
rect 32321 39049 32355 39083
rect 47869 39049 47903 39083
rect 1593 38913 1627 38947
rect 14105 38913 14139 38947
rect 14841 38913 14875 38947
rect 15108 38913 15142 38947
rect 17233 38913 17267 38947
rect 17500 38913 17534 38947
rect 19625 38913 19659 38947
rect 20269 38913 20303 38947
rect 22385 38913 22419 38947
rect 24225 38913 24259 38947
rect 24685 38913 24719 38947
rect 25329 38913 25363 38947
rect 26065 38913 26099 38947
rect 29276 38913 29310 38947
rect 30941 38913 30975 38947
rect 32597 38913 32631 38947
rect 32781 38913 32815 38947
rect 33057 38913 33091 38947
rect 34069 38913 34103 38947
rect 35348 38913 35382 38947
rect 47777 38913 47811 38947
rect 14381 38845 14415 38879
rect 19441 38845 19475 38879
rect 22477 38845 22511 38879
rect 23213 38845 23247 38879
rect 24961 38845 24995 38879
rect 26157 38845 26191 38879
rect 29009 38845 29043 38879
rect 33977 38845 34011 38879
rect 35081 38845 35115 38879
rect 23489 38777 23523 38811
rect 25605 38777 25639 38811
rect 26433 38777 26467 38811
rect 1777 38709 1811 38743
rect 14289 38709 14323 38743
rect 16221 38709 16255 38743
rect 18613 38709 18647 38743
rect 22569 38709 22603 38743
rect 22753 38709 22787 38743
rect 23673 38709 23707 38743
rect 26157 38709 26191 38743
rect 32689 38709 32723 38743
rect 32873 38709 32907 38743
rect 34437 38709 34471 38743
rect 36461 38709 36495 38743
rect 14381 38505 14415 38539
rect 22845 38505 22879 38539
rect 24869 38505 24903 38539
rect 25053 38505 25087 38539
rect 29745 38505 29779 38539
rect 32321 38505 32355 38539
rect 32781 38505 32815 38539
rect 35449 38505 35483 38539
rect 23029 38437 23063 38471
rect 28089 38437 28123 38471
rect 34161 38437 34195 38471
rect 20821 38369 20855 38403
rect 32505 38369 32539 38403
rect 33425 38369 33459 38403
rect 34345 38369 34379 38403
rect 14565 38301 14599 38335
rect 14841 38301 14875 38335
rect 15025 38301 15059 38335
rect 15669 38301 15703 38335
rect 15945 38301 15979 38335
rect 16129 38301 16163 38335
rect 16865 38301 16899 38335
rect 17969 38301 18003 38335
rect 18245 38301 18279 38335
rect 18429 38301 18463 38335
rect 23676 38311 23710 38345
rect 23838 38301 23872 38335
rect 23961 38301 23995 38335
rect 24051 38311 24085 38345
rect 24593 38301 24627 38335
rect 27077 38301 27111 38335
rect 27445 38301 27479 38335
rect 28089 38301 28123 38335
rect 28273 38301 28307 38335
rect 29929 38301 29963 38335
rect 30389 38301 30423 38335
rect 30849 38301 30883 38335
rect 32597 38301 32631 38335
rect 33241 38301 33275 38335
rect 33609 38301 33643 38335
rect 34069 38301 34103 38335
rect 34897 38301 34931 38335
rect 35173 38301 35207 38335
rect 35265 38301 35299 38335
rect 47685 38301 47719 38335
rect 17141 38233 17175 38267
rect 19993 38233 20027 38267
rect 21088 38233 21122 38267
rect 22661 38233 22695 38267
rect 25697 38233 25731 38267
rect 26525 38233 26559 38267
rect 27261 38233 27295 38267
rect 27353 38233 27387 38267
rect 30021 38233 30055 38267
rect 30113 38233 30147 38267
rect 30251 38233 30285 38267
rect 31033 38233 31067 38267
rect 32321 38233 32355 38267
rect 34345 38233 34379 38267
rect 35081 38233 35115 38267
rect 15485 38165 15519 38199
rect 17785 38165 17819 38199
rect 20085 38165 20119 38199
rect 22201 38165 22235 38199
rect 22861 38165 22895 38199
rect 23489 38165 23523 38199
rect 27629 38165 27663 38199
rect 31217 38165 31251 38199
rect 33333 38165 33367 38199
rect 33517 38165 33551 38199
rect 15209 37961 15243 37995
rect 17509 37961 17543 37995
rect 19533 37961 19567 37995
rect 25329 37961 25363 37995
rect 28549 37961 28583 37995
rect 30573 37961 30607 37995
rect 32873 37961 32907 37995
rect 22385 37893 22419 37927
rect 27436 37893 27470 37927
rect 34161 37893 34195 37927
rect 12909 37825 12943 37859
rect 15393 37825 15427 37859
rect 15577 37825 15611 37859
rect 17693 37825 17727 37859
rect 17969 37825 18003 37859
rect 19257 37825 19291 37859
rect 20341 37825 20375 37859
rect 22201 37825 22235 37859
rect 22477 37825 22511 37859
rect 22569 37825 22603 37859
rect 23857 37825 23891 37859
rect 25513 37825 25547 37859
rect 25789 37825 25823 37859
rect 25973 37825 26007 37859
rect 26433 37825 26467 37859
rect 26617 37825 26651 37859
rect 30389 37825 30423 37859
rect 30573 37825 30607 37859
rect 32689 37825 32723 37859
rect 32965 37825 32999 37859
rect 33885 37825 33919 37859
rect 34069 37825 34103 37859
rect 34253 37825 34287 37859
rect 47777 37825 47811 37859
rect 15669 37757 15703 37791
rect 17877 37757 17911 37791
rect 20085 37757 20119 37791
rect 23673 37757 23707 37791
rect 23765 37757 23799 37791
rect 23949 37757 23983 37791
rect 27169 37757 27203 37791
rect 22753 37689 22787 37723
rect 12725 37621 12759 37655
rect 21465 37621 21499 37655
rect 23489 37621 23523 37655
rect 26433 37621 26467 37655
rect 32505 37621 32539 37655
rect 34437 37621 34471 37655
rect 47869 37621 47903 37655
rect 17325 37417 17359 37451
rect 18705 37417 18739 37451
rect 22661 37417 22695 37451
rect 23489 37417 23523 37451
rect 27077 37417 27111 37451
rect 27905 37417 27939 37451
rect 33793 37417 33827 37451
rect 25973 37281 26007 37315
rect 26065 37281 26099 37315
rect 27537 37281 27571 37315
rect 48237 37281 48271 37315
rect 1593 37213 1627 37247
rect 12357 37213 12391 37247
rect 12624 37213 12658 37247
rect 16957 37213 16991 37247
rect 17877 37213 17911 37247
rect 18153 37213 18187 37247
rect 18245 37213 18279 37247
rect 18705 37213 18739 37247
rect 18889 37213 18923 37247
rect 20177 37213 20211 37247
rect 21281 37213 21315 37247
rect 21557 37213 21591 37247
rect 21741 37213 21775 37247
rect 22937 37213 22971 37247
rect 23397 37213 23431 37247
rect 23581 37213 23615 37247
rect 24869 37213 24903 37247
rect 25237 37213 25271 37247
rect 25881 37213 25915 37247
rect 26157 37213 26191 37247
rect 27721 37213 27755 37247
rect 33057 37213 33091 37247
rect 33241 37213 33275 37247
rect 33701 37213 33735 37247
rect 33885 37213 33919 37247
rect 34897 37213 34931 37247
rect 46489 37213 46523 37247
rect 17141 37145 17175 37179
rect 19441 37145 19475 37179
rect 22661 37145 22695 37179
rect 22845 37145 22879 37179
rect 25053 37145 25087 37179
rect 26709 37145 26743 37179
rect 26893 37145 26927 37179
rect 32873 37145 32907 37179
rect 35142 37145 35176 37179
rect 46673 37145 46707 37179
rect 1777 37077 1811 37111
rect 13737 37077 13771 37111
rect 21097 37077 21131 37111
rect 25697 37077 25731 37111
rect 36277 37077 36311 37111
rect 13277 36873 13311 36907
rect 13645 36873 13679 36907
rect 13737 36873 13771 36907
rect 15577 36873 15611 36907
rect 15945 36873 15979 36907
rect 20821 36873 20855 36907
rect 22661 36873 22695 36907
rect 26071 36873 26105 36907
rect 29929 36873 29963 36907
rect 32873 36873 32907 36907
rect 33609 36873 33643 36907
rect 18604 36805 18638 36839
rect 20453 36805 20487 36839
rect 25973 36805 26007 36839
rect 20177 36737 20211 36771
rect 20270 36737 20304 36771
rect 20545 36737 20579 36771
rect 20642 36737 20676 36771
rect 22569 36737 22603 36771
rect 22753 36737 22787 36771
rect 24593 36737 24627 36771
rect 26157 36737 26191 36771
rect 26249 36737 26283 36771
rect 28549 36737 28583 36771
rect 28805 36737 28839 36771
rect 32689 36737 32723 36771
rect 32965 36737 32999 36771
rect 33425 36737 33459 36771
rect 33609 36737 33643 36771
rect 13921 36669 13955 36703
rect 16037 36669 16071 36703
rect 16129 36669 16163 36703
rect 18337 36669 18371 36703
rect 25329 36669 25363 36703
rect 19717 36533 19751 36567
rect 32505 36533 32539 36567
rect 47961 36533 47995 36567
rect 16589 36329 16623 36363
rect 20177 36329 20211 36363
rect 26341 36329 26375 36363
rect 28273 36329 28307 36363
rect 32321 36329 32355 36363
rect 33977 36329 34011 36363
rect 15485 36193 15519 36227
rect 16405 36193 16439 36227
rect 20637 36193 20671 36227
rect 24685 36193 24719 36227
rect 25421 36193 25455 36227
rect 25513 36193 25547 36227
rect 33425 36193 33459 36227
rect 46489 36193 46523 36227
rect 48237 36193 48271 36227
rect 12357 36125 12391 36159
rect 15209 36125 15243 36159
rect 16313 36125 16347 36159
rect 19441 36125 19475 36159
rect 19625 36125 19659 36159
rect 20361 36125 20395 36159
rect 20545 36125 20579 36159
rect 22201 36125 22235 36159
rect 22385 36125 22419 36159
rect 24593 36125 24627 36159
rect 24777 36125 24811 36159
rect 25605 36125 25639 36159
rect 25697 36125 25731 36159
rect 26249 36125 26283 36159
rect 26433 36125 26467 36159
rect 26893 36125 26927 36159
rect 27077 36125 27111 36159
rect 28457 36125 28491 36159
rect 28733 36125 28767 36159
rect 30941 36125 30975 36159
rect 32965 36125 32999 36159
rect 33057 36125 33091 36159
rect 33885 36125 33919 36159
rect 12624 36057 12658 36091
rect 31208 36057 31242 36091
rect 32781 36057 32815 36091
rect 33149 36057 33183 36091
rect 33267 36057 33301 36091
rect 46673 36057 46707 36091
rect 13737 35989 13771 36023
rect 14841 35989 14875 36023
rect 15301 35989 15335 36023
rect 19533 35989 19567 36023
rect 22385 35989 22419 36023
rect 25237 35989 25271 36023
rect 26985 35989 27019 36023
rect 28641 35989 28675 36023
rect 12817 35785 12851 35819
rect 13829 35785 13863 35819
rect 13921 35785 13955 35819
rect 16957 35785 16991 35819
rect 18797 35785 18831 35819
rect 23397 35785 23431 35819
rect 25145 35785 25179 35819
rect 26249 35785 26283 35819
rect 33425 35785 33459 35819
rect 47869 35785 47903 35819
rect 14657 35717 14691 35751
rect 15669 35717 15703 35751
rect 25053 35717 25087 35751
rect 25881 35717 25915 35751
rect 30481 35717 30515 35751
rect 33517 35717 33551 35751
rect 13001 35649 13035 35683
rect 14841 35649 14875 35683
rect 15025 35649 15059 35683
rect 16129 35649 16163 35683
rect 16865 35649 16899 35683
rect 17049 35649 17083 35683
rect 17693 35649 17727 35683
rect 17877 35649 17911 35683
rect 17969 35649 18003 35683
rect 18981 35649 19015 35683
rect 19073 35649 19107 35683
rect 19257 35649 19291 35683
rect 19441 35649 19475 35683
rect 20085 35649 20119 35683
rect 22273 35649 22307 35683
rect 26065 35649 26099 35683
rect 28365 35649 28399 35683
rect 28632 35649 28666 35683
rect 30205 35649 30239 35683
rect 32505 35649 32539 35683
rect 33333 35649 33367 35683
rect 33609 35649 33643 35683
rect 47777 35649 47811 35683
rect 14105 35581 14139 35615
rect 16037 35581 16071 35615
rect 19901 35581 19935 35615
rect 22017 35581 22051 35615
rect 25329 35581 25363 35615
rect 32597 35581 32631 35615
rect 32873 35581 32907 35615
rect 13461 35513 13495 35547
rect 17693 35513 17727 35547
rect 19165 35513 19199 35547
rect 16313 35445 16347 35479
rect 20269 35445 20303 35479
rect 24685 35445 24719 35479
rect 29745 35445 29779 35479
rect 15853 35241 15887 35275
rect 17417 35241 17451 35275
rect 19625 35241 19659 35275
rect 22661 35241 22695 35275
rect 25973 35241 26007 35275
rect 13645 35173 13679 35207
rect 17325 35173 17359 35207
rect 19533 35173 19567 35207
rect 15669 35105 15703 35139
rect 19717 35105 19751 35139
rect 21649 35105 21683 35139
rect 27353 35105 27387 35139
rect 13553 35037 13587 35071
rect 13737 35037 13771 35071
rect 14565 35037 14599 35071
rect 14749 35037 14783 35071
rect 15577 35037 15611 35071
rect 17233 35037 17267 35071
rect 17693 35037 17727 35071
rect 18521 35037 18555 35071
rect 18705 35037 18739 35071
rect 19441 35037 19475 35071
rect 21746 35037 21780 35071
rect 22293 35037 22327 35071
rect 22569 35037 22603 35071
rect 23489 35037 23523 35071
rect 24593 35037 24627 35071
rect 27169 35037 27203 35071
rect 27445 35037 27479 35071
rect 28733 35037 28767 35071
rect 29009 35037 29043 35071
rect 29193 35037 29227 35071
rect 30757 35037 30791 35071
rect 31033 35037 31067 35071
rect 21373 34969 21407 35003
rect 21557 34969 21591 35003
rect 21649 34969 21683 35003
rect 23305 34969 23339 35003
rect 24838 34969 24872 35003
rect 30941 34969 30975 35003
rect 14657 34901 14691 34935
rect 16957 34901 16991 34935
rect 17601 34901 17635 34935
rect 18613 34901 18647 34935
rect 22845 34901 22879 34935
rect 23673 34901 23707 34935
rect 26985 34901 27019 34935
rect 28549 34901 28583 34935
rect 30573 34901 30607 34935
rect 15853 34697 15887 34731
rect 22109 34697 22143 34731
rect 23229 34697 23263 34731
rect 23397 34697 23431 34731
rect 24409 34697 24443 34731
rect 25421 34697 25455 34731
rect 28549 34697 28583 34731
rect 29009 34697 29043 34731
rect 23029 34629 23063 34663
rect 27414 34629 27448 34663
rect 30564 34629 30598 34663
rect 1593 34561 1627 34595
rect 14565 34561 14599 34595
rect 14749 34561 14783 34595
rect 15393 34561 15427 34595
rect 22293 34561 22327 34595
rect 22477 34561 22511 34595
rect 22569 34561 22603 34595
rect 24593 34561 24627 34595
rect 25237 34561 25271 34595
rect 26065 34561 26099 34595
rect 26249 34561 26283 34595
rect 27169 34561 27203 34595
rect 29193 34561 29227 34595
rect 30297 34561 30331 34595
rect 14657 34493 14691 34527
rect 25053 34493 25087 34527
rect 26341 34493 26375 34527
rect 29377 34493 29411 34527
rect 29469 34493 29503 34527
rect 25881 34425 25915 34459
rect 1777 34357 1811 34391
rect 15485 34357 15519 34391
rect 23213 34357 23247 34391
rect 31677 34357 31711 34391
rect 13185 34153 13219 34187
rect 21925 34153 21959 34187
rect 22661 34153 22695 34187
rect 26985 34153 27019 34187
rect 30481 34153 30515 34187
rect 31309 34153 31343 34187
rect 11805 34017 11839 34051
rect 15761 34017 15795 34051
rect 20361 34017 20395 34051
rect 15025 33949 15059 33983
rect 15209 33949 15243 33983
rect 15301 33949 15335 33983
rect 20177 33949 20211 33983
rect 20453 33949 20487 33983
rect 21833 33949 21867 33983
rect 22017 33949 22051 33983
rect 22569 33949 22603 33983
rect 22753 33949 22787 33983
rect 27169 33949 27203 33983
rect 27445 33949 27479 33983
rect 27629 33949 27663 33983
rect 29929 33949 29963 33983
rect 30205 33949 30239 33983
rect 30297 33949 30331 33983
rect 31309 33949 31343 33983
rect 31493 33949 31527 33983
rect 12072 33881 12106 33915
rect 16028 33881 16062 33915
rect 30113 33881 30147 33915
rect 14841 33813 14875 33847
rect 17141 33813 17175 33847
rect 19993 33813 20027 33847
rect 11989 33609 12023 33643
rect 14289 33609 14323 33643
rect 16865 33609 16899 33643
rect 20913 33609 20947 33643
rect 19800 33541 19834 33575
rect 12173 33473 12207 33507
rect 12909 33473 12943 33507
rect 13176 33473 13210 33507
rect 14933 33473 14967 33507
rect 15209 33473 15243 33507
rect 15393 33473 15427 33507
rect 17049 33473 17083 33507
rect 17233 33473 17267 33507
rect 18245 33473 18279 33507
rect 19533 33473 19567 33507
rect 31401 33473 31435 33507
rect 35909 33473 35943 33507
rect 12449 33405 12483 33439
rect 17325 33405 17359 33439
rect 18521 33405 18555 33439
rect 31217 33405 31251 33439
rect 36645 33405 36679 33439
rect 12357 33269 12391 33303
rect 14749 33269 14783 33303
rect 18061 33269 18095 33303
rect 18429 33269 18463 33303
rect 31585 33269 31619 33303
rect 47961 33269 47995 33303
rect 12357 33065 12391 33099
rect 14289 33065 14323 33099
rect 16405 33065 16439 33099
rect 20453 33065 20487 33099
rect 22753 33065 22787 33099
rect 25973 33065 26007 33099
rect 28825 33065 28859 33099
rect 31217 33065 31251 33099
rect 31861 32997 31895 33031
rect 14749 32929 14783 32963
rect 17509 32929 17543 32963
rect 24593 32929 24627 32963
rect 28917 32929 28951 32963
rect 46489 32929 46523 32963
rect 2053 32861 2087 32895
rect 2513 32861 2547 32895
rect 12541 32861 12575 32895
rect 12817 32861 12851 32895
rect 13001 32861 13035 32895
rect 14473 32861 14507 32895
rect 14657 32861 14691 32895
rect 16589 32861 16623 32895
rect 16865 32861 16899 32895
rect 17049 32861 17083 32895
rect 17776 32861 17810 32895
rect 20637 32861 20671 32895
rect 20913 32861 20947 32895
rect 21097 32861 21131 32895
rect 21833 32861 21867 32895
rect 22109 32861 22143 32895
rect 22293 32861 22327 32895
rect 22937 32861 22971 32895
rect 23213 32861 23247 32895
rect 28641 32861 28675 32895
rect 31217 32861 31251 32895
rect 31401 32861 31435 32895
rect 32137 32861 32171 32895
rect 24838 32793 24872 32827
rect 31861 32793 31895 32827
rect 46673 32793 46707 32827
rect 48329 32793 48363 32827
rect 2605 32725 2639 32759
rect 18889 32725 18923 32759
rect 21649 32725 21683 32759
rect 23121 32725 23155 32759
rect 28457 32725 28491 32759
rect 32045 32725 32079 32759
rect 15761 32521 15795 32555
rect 18245 32521 18279 32555
rect 23397 32521 23431 32555
rect 23949 32521 23983 32555
rect 47869 32521 47903 32555
rect 2329 32453 2363 32487
rect 31401 32453 31435 32487
rect 2145 32385 2179 32419
rect 18429 32385 18463 32419
rect 18705 32385 18739 32419
rect 18889 32385 18923 32419
rect 22017 32385 22051 32419
rect 22273 32385 22307 32419
rect 24133 32385 24167 32419
rect 24869 32385 24903 32419
rect 25053 32385 25087 32419
rect 25329 32385 25363 32419
rect 25513 32385 25547 32419
rect 27425 32385 27459 32419
rect 29009 32385 29043 32419
rect 29265 32385 29299 32419
rect 31125 32385 31159 32419
rect 31273 32385 31307 32419
rect 31493 32385 31527 32419
rect 31590 32385 31624 32419
rect 32321 32385 32355 32419
rect 32577 32385 32611 32419
rect 47777 32385 47811 32419
rect 2789 32317 2823 32351
rect 15853 32317 15887 32351
rect 16037 32317 16071 32351
rect 24409 32317 24443 32351
rect 27169 32317 27203 32351
rect 31769 32249 31803 32283
rect 15393 32181 15427 32215
rect 24317 32181 24351 32215
rect 28549 32181 28583 32215
rect 30389 32181 30423 32215
rect 33701 32181 33735 32215
rect 21925 31977 21959 32011
rect 23949 31977 23983 32011
rect 25973 31977 26007 32011
rect 28549 31977 28583 32011
rect 31677 31977 31711 32011
rect 32045 31977 32079 32011
rect 32597 31909 32631 31943
rect 1593 31841 1627 31875
rect 20545 31841 20579 31875
rect 23581 31841 23615 31875
rect 24593 31841 24627 31875
rect 32137 31841 32171 31875
rect 1869 31773 1903 31807
rect 12633 31773 12667 31807
rect 16313 31773 16347 31807
rect 16497 31773 16531 31807
rect 22661 31773 22695 31807
rect 22937 31773 22971 31807
rect 23121 31773 23155 31807
rect 23765 31773 23799 31807
rect 24041 31773 24075 31807
rect 24849 31773 24883 31807
rect 26985 31773 27019 31807
rect 27261 31773 27295 31807
rect 27445 31773 27479 31807
rect 28733 31773 28767 31807
rect 29009 31773 29043 31807
rect 29193 31773 29227 31807
rect 31861 31773 31895 31807
rect 32781 31773 32815 31807
rect 32873 31773 32907 31807
rect 20812 31705 20846 31739
rect 32597 31705 32631 31739
rect 12449 31637 12483 31671
rect 16497 31637 16531 31671
rect 22477 31637 22511 31671
rect 26801 31637 26835 31671
rect 13829 31433 13863 31467
rect 14289 31433 14323 31467
rect 21005 31433 21039 31467
rect 22109 31433 22143 31467
rect 24685 31433 24719 31467
rect 27169 31433 27203 31467
rect 31309 31433 31343 31467
rect 12256 31365 12290 31399
rect 4620 31297 4654 31331
rect 8401 31297 8435 31331
rect 11989 31297 12023 31331
rect 14197 31297 14231 31331
rect 15485 31297 15519 31331
rect 16865 31297 16899 31331
rect 17049 31297 17083 31331
rect 17601 31297 17635 31331
rect 17785 31297 17819 31331
rect 21189 31297 21223 31331
rect 22293 31297 22327 31331
rect 24869 31297 24903 31331
rect 25145 31297 25179 31331
rect 25329 31297 25363 31331
rect 27353 31297 27387 31331
rect 29929 31297 29963 31331
rect 30196 31297 30230 31331
rect 32505 31297 32539 31331
rect 4353 31229 4387 31263
rect 14473 31229 14507 31263
rect 15577 31229 15611 31263
rect 15853 31229 15887 31263
rect 21465 31229 21499 31263
rect 22569 31229 22603 31263
rect 27629 31229 27663 31263
rect 32597 31229 32631 31263
rect 32873 31229 32907 31263
rect 17693 31161 17727 31195
rect 5733 31093 5767 31127
rect 8217 31093 8251 31127
rect 13369 31093 13403 31127
rect 16957 31093 16991 31127
rect 21373 31093 21407 31127
rect 22477 31093 22511 31127
rect 27537 31093 27571 31127
rect 5365 30889 5399 30923
rect 6009 30889 6043 30923
rect 12541 30889 12575 30923
rect 17141 30889 17175 30923
rect 18061 30889 18095 30923
rect 32413 30889 32447 30923
rect 15117 30821 15151 30855
rect 16313 30821 16347 30855
rect 16497 30821 16531 30855
rect 17049 30821 17083 30855
rect 17693 30821 17727 30855
rect 18705 30821 18739 30855
rect 7205 30753 7239 30787
rect 9137 30753 9171 30787
rect 14381 30753 14415 30787
rect 16037 30753 16071 30787
rect 17233 30753 17267 30787
rect 19441 30753 19475 30787
rect 5089 30685 5123 30719
rect 6193 30685 6227 30719
rect 7472 30685 7506 30719
rect 12357 30685 12391 30719
rect 12633 30685 12667 30719
rect 13553 30685 13587 30719
rect 13737 30685 13771 30719
rect 14289 30685 14323 30719
rect 14473 30685 14507 30719
rect 15301 30685 15335 30719
rect 15577 30685 15611 30719
rect 16957 30685 16991 30719
rect 18705 30685 18739 30719
rect 18889 30685 18923 30719
rect 28641 30685 28675 30719
rect 28825 30685 28859 30719
rect 30573 30685 30607 30719
rect 30849 30685 30883 30719
rect 31033 30685 31067 30719
rect 32137 30685 32171 30719
rect 32229 30685 32263 30719
rect 9404 30617 9438 30651
rect 19686 30617 19720 30651
rect 5549 30549 5583 30583
rect 8585 30549 8619 30583
rect 10517 30549 10551 30583
rect 12173 30549 12207 30583
rect 13737 30549 13771 30583
rect 15485 30549 15519 30583
rect 18061 30549 18095 30583
rect 18245 30549 18279 30583
rect 20821 30549 20855 30583
rect 28825 30549 28859 30583
rect 30389 30549 30423 30583
rect 6009 30345 6043 30379
rect 9045 30345 9079 30379
rect 9505 30345 9539 30379
rect 24409 30345 24443 30379
rect 30205 30345 30239 30379
rect 6653 30277 6687 30311
rect 17049 30277 17083 30311
rect 17233 30277 17267 30311
rect 17785 30277 17819 30311
rect 18889 30277 18923 30311
rect 18981 30277 19015 30311
rect 22385 30277 22419 30311
rect 22937 30277 22971 30311
rect 23153 30277 23187 30311
rect 24317 30277 24351 30311
rect 27905 30277 27939 30311
rect 5089 30209 5123 30243
rect 5549 30209 5583 30243
rect 6837 30209 6871 30243
rect 7481 30209 7515 30243
rect 8585 30209 8619 30243
rect 9689 30209 9723 30243
rect 12256 30209 12290 30243
rect 15209 30209 15243 30243
rect 15485 30209 15519 30243
rect 16865 30209 16899 30243
rect 17693 30209 17727 30243
rect 17877 30209 17911 30243
rect 18613 30209 18647 30243
rect 18761 30209 18795 30243
rect 19078 30209 19112 30243
rect 22201 30209 22235 30243
rect 22477 30209 22511 30243
rect 26065 30209 26099 30243
rect 26341 30209 26375 30243
rect 26525 30209 26559 30243
rect 28089 30209 28123 30243
rect 28365 30209 28399 30243
rect 29009 30209 29043 30243
rect 30389 30209 30423 30243
rect 30665 30209 30699 30243
rect 47777 30209 47811 30243
rect 7757 30141 7791 30175
rect 11989 30141 12023 30175
rect 28273 30141 28307 30175
rect 29101 30141 29135 30175
rect 7665 30073 7699 30107
rect 19257 30073 19291 30107
rect 4905 30005 4939 30039
rect 5825 30005 5859 30039
rect 7573 30005 7607 30039
rect 8861 30005 8895 30039
rect 13369 30005 13403 30039
rect 15577 30005 15611 30039
rect 15761 30005 15795 30039
rect 22017 30005 22051 30039
rect 23121 30005 23155 30039
rect 23305 30005 23339 30039
rect 25881 30005 25915 30039
rect 29377 30005 29411 30039
rect 30573 30005 30607 30039
rect 47225 30005 47259 30039
rect 47869 30005 47903 30039
rect 12449 29801 12483 29835
rect 15761 29801 15795 29835
rect 20637 29801 20671 29835
rect 22109 29801 22143 29835
rect 23121 29801 23155 29835
rect 30113 29801 30147 29835
rect 15853 29733 15887 29767
rect 20913 29733 20947 29767
rect 22753 29733 22787 29767
rect 6929 29665 6963 29699
rect 15485 29665 15519 29699
rect 21649 29665 21683 29699
rect 25421 29665 25455 29699
rect 46489 29665 46523 29699
rect 46673 29665 46707 29699
rect 4353 29597 4387 29631
rect 4620 29597 4654 29631
rect 12633 29597 12667 29631
rect 12909 29597 12943 29631
rect 13093 29597 13127 29631
rect 15945 29597 15979 29631
rect 16221 29597 16255 29631
rect 20361 29597 20395 29631
rect 20729 29597 20763 29631
rect 21373 29597 21407 29631
rect 21557 29597 21591 29631
rect 21741 29597 21775 29631
rect 21925 29597 21959 29631
rect 23857 29597 23891 29631
rect 24041 29597 24075 29631
rect 24777 29597 24811 29631
rect 27353 29597 27387 29631
rect 29929 29597 29963 29631
rect 7196 29529 7230 29563
rect 23121 29529 23155 29563
rect 24593 29529 24627 29563
rect 25688 29529 25722 29563
rect 27620 29529 27654 29563
rect 29745 29529 29779 29563
rect 48329 29529 48363 29563
rect 5733 29461 5767 29495
rect 8309 29461 8343 29495
rect 16129 29461 16163 29495
rect 23305 29461 23339 29495
rect 23949 29461 23983 29495
rect 24961 29461 24995 29495
rect 26801 29461 26835 29495
rect 28733 29461 28767 29495
rect 7297 29257 7331 29291
rect 7665 29257 7699 29291
rect 8677 29257 8711 29291
rect 17065 29257 17099 29291
rect 25697 29257 25731 29291
rect 26157 29257 26191 29291
rect 27997 29257 28031 29291
rect 28089 29257 28123 29291
rect 28825 29257 28859 29291
rect 29285 29257 29319 29291
rect 16129 29189 16163 29223
rect 16865 29189 16899 29223
rect 21005 29189 21039 29223
rect 23581 29189 23615 29223
rect 5181 29121 5215 29155
rect 7481 29121 7515 29155
rect 7757 29121 7791 29155
rect 8217 29121 8251 29155
rect 15945 29121 15979 29155
rect 16221 29121 16255 29155
rect 22385 29121 22419 29155
rect 22661 29121 22695 29155
rect 23213 29121 23247 29155
rect 23361 29121 23395 29155
rect 23489 29121 23523 29155
rect 23719 29121 23753 29155
rect 24317 29121 24351 29155
rect 24573 29121 24607 29155
rect 26341 29121 26375 29155
rect 26525 29121 26559 29155
rect 29193 29121 29227 29155
rect 30849 29121 30883 29155
rect 47777 29121 47811 29155
rect 15761 29053 15795 29087
rect 22477 29053 22511 29087
rect 22569 29053 22603 29087
rect 26617 29053 26651 29087
rect 28181 29053 28215 29087
rect 29377 29053 29411 29087
rect 31125 29053 31159 29087
rect 21281 28985 21315 29019
rect 21465 28985 21499 29019
rect 23857 28985 23891 29019
rect 31033 28985 31067 29019
rect 5457 28917 5491 28951
rect 5641 28917 5675 28951
rect 8309 28917 8343 28951
rect 17049 28917 17083 28951
rect 17233 28917 17267 28951
rect 22201 28917 22235 28951
rect 27629 28917 27663 28951
rect 30665 28917 30699 28951
rect 47225 28917 47259 28951
rect 47869 28917 47903 28951
rect 9229 28713 9263 28747
rect 23581 28713 23615 28747
rect 27537 28713 27571 28747
rect 28457 28713 28491 28747
rect 32137 28713 32171 28747
rect 15485 28577 15519 28611
rect 15669 28577 15703 28611
rect 21005 28577 21039 28611
rect 30757 28577 30791 28611
rect 46489 28577 46523 28611
rect 48237 28577 48271 28611
rect 5181 28509 5215 28543
rect 9137 28509 9171 28543
rect 13461 28509 13495 28543
rect 13645 28509 13679 28543
rect 15393 28509 15427 28543
rect 15577 28509 15611 28543
rect 16405 28509 16439 28543
rect 16681 28509 16715 28543
rect 17509 28509 17543 28543
rect 22109 28509 22143 28543
rect 22385 28509 22419 28543
rect 23489 28509 23523 28543
rect 23673 28509 23707 28543
rect 27721 28509 27755 28543
rect 28365 28509 28399 28543
rect 28549 28509 28583 28543
rect 31013 28509 31047 28543
rect 36553 28509 36587 28543
rect 17776 28441 17810 28475
rect 37381 28441 37415 28475
rect 46673 28441 46707 28475
rect 4997 28373 5031 28407
rect 13553 28373 13587 28407
rect 15209 28373 15243 28407
rect 16221 28373 16255 28407
rect 16589 28373 16623 28407
rect 18889 28373 18923 28407
rect 20453 28373 20487 28407
rect 20821 28373 20855 28407
rect 20913 28373 20947 28407
rect 22207 28373 22241 28407
rect 22293 28373 22327 28407
rect 13369 28169 13403 28203
rect 15301 28169 15335 28203
rect 17601 28169 17635 28203
rect 18889 28169 18923 28203
rect 20821 28169 20855 28203
rect 22109 28169 22143 28203
rect 30665 28169 30699 28203
rect 4620 28101 4654 28135
rect 7941 28101 7975 28135
rect 14565 28101 14599 28135
rect 17417 28101 17451 28135
rect 18521 28101 18555 28135
rect 18613 28101 18647 28135
rect 21373 28101 21407 28135
rect 4353 28033 4387 28067
rect 8953 28033 8987 28067
rect 13461 28033 13495 28067
rect 14749 28033 14783 28067
rect 14841 28033 14875 28067
rect 15577 28033 15611 28067
rect 15666 28033 15700 28067
rect 15761 28036 15795 28070
rect 15945 28033 15979 28067
rect 17049 28033 17083 28067
rect 18245 28033 18279 28067
rect 18393 28033 18427 28067
rect 18751 28033 18785 28067
rect 19708 28033 19742 28067
rect 21281 28033 21315 28067
rect 21465 28033 21499 28067
rect 22293 28033 22327 28067
rect 22385 28033 22419 28067
rect 22661 28033 22695 28067
rect 24593 28033 24627 28067
rect 30849 28033 30883 28067
rect 31125 28033 31159 28067
rect 31309 28033 31343 28067
rect 47777 28033 47811 28067
rect 8861 27965 8895 27999
rect 13645 27965 13679 27999
rect 19441 27965 19475 27999
rect 22569 27965 22603 27999
rect 24869 27965 24903 27999
rect 9321 27897 9355 27931
rect 24409 27897 24443 27931
rect 5733 27829 5767 27863
rect 8033 27829 8067 27863
rect 13001 27829 13035 27863
rect 14565 27829 14599 27863
rect 17417 27829 17451 27863
rect 24777 27829 24811 27863
rect 47225 27829 47259 27863
rect 47869 27829 47903 27863
rect 4813 27625 4847 27659
rect 5733 27625 5767 27659
rect 8401 27625 8435 27659
rect 19993 27625 20027 27659
rect 14381 27557 14415 27591
rect 15393 27557 15427 27591
rect 18153 27557 18187 27591
rect 21005 27557 21039 27591
rect 26617 27557 26651 27591
rect 29101 27557 29135 27591
rect 4997 27489 5031 27523
rect 12081 27489 12115 27523
rect 14841 27489 14875 27523
rect 15761 27489 15795 27523
rect 16957 27489 16991 27523
rect 46489 27489 46523 27523
rect 48237 27489 48271 27523
rect 4537 27421 4571 27455
rect 5457 27421 5491 27455
rect 6561 27421 6595 27455
rect 8125 27421 8159 27455
rect 14565 27421 14599 27455
rect 14657 27421 14691 27455
rect 14933 27421 14967 27455
rect 15577 27421 15611 27455
rect 15669 27421 15703 27455
rect 15853 27421 15887 27455
rect 16589 27421 16623 27455
rect 17417 27421 17451 27455
rect 17601 27421 17635 27455
rect 18061 27421 18095 27455
rect 18245 27421 18279 27455
rect 20177 27421 20211 27455
rect 20913 27421 20947 27455
rect 21097 27421 21131 27455
rect 24593 27421 24627 27455
rect 26433 27421 26467 27455
rect 28917 27421 28951 27455
rect 29193 27421 29227 27455
rect 31217 27421 31251 27455
rect 33609 27421 33643 27455
rect 34897 27421 34931 27455
rect 35081 27421 35115 27455
rect 35725 27421 35759 27455
rect 35909 27421 35943 27455
rect 38117 27421 38151 27455
rect 12348 27353 12382 27387
rect 16773 27353 16807 27387
rect 24860 27353 24894 27387
rect 31462 27353 31496 27387
rect 35265 27353 35299 27387
rect 38384 27353 38418 27387
rect 46673 27353 46707 27387
rect 5917 27285 5951 27319
rect 6377 27285 6411 27319
rect 8585 27285 8619 27319
rect 13461 27285 13495 27319
rect 17601 27285 17635 27319
rect 25973 27285 26007 27319
rect 28733 27285 28767 27319
rect 32597 27285 32631 27319
rect 33425 27285 33459 27319
rect 35817 27285 35851 27319
rect 39497 27285 39531 27319
rect 5733 27081 5767 27115
rect 7389 27081 7423 27115
rect 9413 27081 9447 27115
rect 12541 27081 12575 27115
rect 14565 27081 14599 27115
rect 16037 27081 16071 27115
rect 17325 27081 17359 27115
rect 24409 27081 24443 27115
rect 28549 27081 28583 27115
rect 36001 27081 36035 27115
rect 38577 27081 38611 27115
rect 4620 27013 4654 27047
rect 8278 27013 8312 27047
rect 26617 27013 26651 27047
rect 29254 27013 29288 27047
rect 35265 27013 35299 27047
rect 4353 26945 4387 26979
rect 6745 26945 6779 26979
rect 7573 26945 7607 26979
rect 12725 26945 12759 26979
rect 13553 26945 13587 26979
rect 13737 26945 13771 26979
rect 14381 26945 14415 26979
rect 15945 26945 15979 26979
rect 17233 26945 17267 26979
rect 20545 26945 20579 26979
rect 20729 26945 20763 26979
rect 22477 26945 22511 26979
rect 24593 26945 24627 26979
rect 24869 26945 24903 26979
rect 25053 26945 25087 26979
rect 25881 26945 25915 26979
rect 26341 26945 26375 26979
rect 27169 26945 27203 26979
rect 27425 26945 27459 26979
rect 29009 26945 29043 26979
rect 31309 26945 31343 26979
rect 31585 26945 31619 26979
rect 31769 26945 31803 26979
rect 33508 26945 33542 26979
rect 35081 26945 35115 26979
rect 35909 26945 35943 26979
rect 36093 26945 36127 26979
rect 37657 26945 37691 26979
rect 37933 26945 37967 26979
rect 38117 26945 38151 26979
rect 38761 26945 38795 26979
rect 39037 26945 39071 26979
rect 8033 26877 8067 26911
rect 14197 26877 14231 26911
rect 20821 26877 20855 26911
rect 22753 26877 22787 26911
rect 33241 26877 33275 26911
rect 37473 26877 37507 26911
rect 6561 26741 6595 26775
rect 20361 26741 20395 26775
rect 22293 26741 22327 26775
rect 22661 26741 22695 26775
rect 30389 26741 30423 26775
rect 31125 26741 31159 26775
rect 34621 26741 34655 26775
rect 35449 26741 35483 26775
rect 38945 26741 38979 26775
rect 47961 26741 47995 26775
rect 8493 26537 8527 26571
rect 13553 26537 13587 26571
rect 17969 26537 18003 26571
rect 21097 26537 21131 26571
rect 23397 26537 23431 26571
rect 24961 26537 24995 26571
rect 31033 26537 31067 26571
rect 6653 26469 6687 26503
rect 18429 26469 18463 26503
rect 25697 26469 25731 26503
rect 26525 26469 26559 26503
rect 28549 26469 28583 26503
rect 39405 26469 39439 26503
rect 19717 26401 19751 26435
rect 32781 26401 32815 26435
rect 35173 26401 35207 26435
rect 37933 26401 37967 26435
rect 46489 26401 46523 26435
rect 48237 26401 48271 26435
rect 5273 26333 5307 26367
rect 5540 26333 5574 26367
rect 7113 26333 7147 26367
rect 13461 26333 13495 26367
rect 13645 26333 13679 26367
rect 16589 26333 16623 26367
rect 18613 26333 18647 26367
rect 18705 26333 18739 26367
rect 19984 26333 20018 26367
rect 22017 26333 22051 26367
rect 24685 26333 24719 26367
rect 25513 26333 25547 26367
rect 27353 26333 27387 26367
rect 27629 26333 27663 26367
rect 27813 26333 27847 26367
rect 28733 26333 28767 26367
rect 29009 26333 29043 26367
rect 29193 26333 29227 26367
rect 31953 26333 31987 26367
rect 33333 26333 33367 26367
rect 35081 26333 35115 26367
rect 36369 26333 36403 26367
rect 36553 26333 36587 26367
rect 38117 26333 38151 26367
rect 38393 26333 38427 26367
rect 38577 26333 38611 26367
rect 39221 26333 39255 26367
rect 39497 26333 39531 26367
rect 7380 26265 7414 26299
rect 16856 26265 16890 26299
rect 18429 26265 18463 26299
rect 22284 26265 22318 26299
rect 26341 26265 26375 26299
rect 29745 26265 29779 26299
rect 34069 26265 34103 26299
rect 36737 26265 36771 26299
rect 46673 26265 46707 26299
rect 27169 26197 27203 26231
rect 35449 26197 35483 26231
rect 39037 26197 39071 26231
rect 7757 25993 7791 26027
rect 17877 25993 17911 26027
rect 20545 25993 20579 26027
rect 22477 25993 22511 26027
rect 26065 25993 26099 26027
rect 27169 25993 27203 26027
rect 31309 25993 31343 26027
rect 33517 25993 33551 26027
rect 33977 25993 34011 26027
rect 34713 25993 34747 26027
rect 35173 25993 35207 26027
rect 40693 25993 40727 26027
rect 47869 25993 47903 26027
rect 25881 25925 25915 25959
rect 35081 25925 35115 25959
rect 36001 25925 36035 25959
rect 36201 25925 36235 25959
rect 39558 25925 39592 25959
rect 2237 25857 2271 25891
rect 6837 25857 6871 25891
rect 7941 25857 7975 25891
rect 12725 25857 12759 25891
rect 13001 25857 13035 25891
rect 13185 25857 13219 25891
rect 15669 25857 15703 25891
rect 15945 25857 15979 25891
rect 16129 25857 16163 25891
rect 18061 25857 18095 25891
rect 20729 25857 20763 25891
rect 21005 25857 21039 25891
rect 21189 25857 21223 25891
rect 22661 25857 22695 25891
rect 22937 25857 22971 25891
rect 23121 25857 23155 25891
rect 25697 25857 25731 25891
rect 27353 25857 27387 25891
rect 28181 25857 28215 25891
rect 30113 25857 30147 25891
rect 31493 25857 31527 25891
rect 31781 25857 31815 25891
rect 32321 25857 32355 25891
rect 33885 25857 33919 25891
rect 38301 25857 38335 25891
rect 38577 25857 38611 25891
rect 38761 25857 38795 25891
rect 47777 25857 47811 25891
rect 7297 25789 7331 25823
rect 18337 25789 18371 25823
rect 27629 25789 27663 25823
rect 34161 25789 34195 25823
rect 35357 25789 35391 25823
rect 39313 25789 39347 25823
rect 2329 25653 2363 25687
rect 6929 25653 6963 25687
rect 12541 25653 12575 25687
rect 15485 25653 15519 25687
rect 18245 25653 18279 25687
rect 27537 25653 27571 25687
rect 28273 25653 28307 25687
rect 30297 25653 30331 25687
rect 31677 25653 31711 25687
rect 32505 25653 32539 25687
rect 36185 25653 36219 25687
rect 36369 25653 36403 25687
rect 38117 25653 38151 25687
rect 47225 25653 47259 25687
rect 13461 25449 13495 25483
rect 16221 25449 16255 25483
rect 18797 25449 18831 25483
rect 25697 25449 25731 25483
rect 32505 25449 32539 25483
rect 1777 25313 1811 25347
rect 2789 25313 2823 25347
rect 12081 25313 12115 25347
rect 18889 25313 18923 25347
rect 23673 25313 23707 25347
rect 24961 25313 24995 25347
rect 36461 25313 36495 25347
rect 46489 25313 46523 25347
rect 48237 25313 48271 25347
rect 1593 25245 1627 25279
rect 14841 25245 14875 25279
rect 16865 25245 16899 25279
rect 17049 25245 17083 25279
rect 17141 25245 17175 25279
rect 18613 25245 18647 25279
rect 19625 25245 19659 25279
rect 19901 25245 19935 25279
rect 20085 25245 20119 25279
rect 21557 25245 21591 25279
rect 25513 25245 25547 25279
rect 27721 25245 27755 25279
rect 30113 25245 30147 25279
rect 30297 25245 30331 25279
rect 30389 25245 30423 25279
rect 31125 25245 31159 25279
rect 35633 25245 35667 25279
rect 35817 25245 35851 25279
rect 36369 25245 36403 25279
rect 36921 25245 36955 25279
rect 37657 25245 37691 25279
rect 12348 25177 12382 25211
rect 15108 25177 15142 25211
rect 16681 25177 16715 25211
rect 19441 25177 19475 25211
rect 23397 25177 23431 25211
rect 24685 25177 24719 25211
rect 31392 25177 31426 25211
rect 36829 25177 36863 25211
rect 37924 25177 37958 25211
rect 46673 25177 46707 25211
rect 18429 25109 18463 25143
rect 21649 25109 21683 25143
rect 27905 25109 27939 25143
rect 29929 25109 29963 25143
rect 39037 25109 39071 25143
rect 12357 24905 12391 24939
rect 19533 24905 19567 24939
rect 21373 24905 21407 24939
rect 31309 24905 31343 24939
rect 38025 24905 38059 24939
rect 18420 24837 18454 24871
rect 23498 24837 23532 24871
rect 29736 24837 29770 24871
rect 36185 24837 36219 24871
rect 2237 24769 2271 24803
rect 12541 24769 12575 24803
rect 13829 24769 13863 24803
rect 14096 24769 14130 24803
rect 15853 24769 15887 24803
rect 16129 24769 16163 24803
rect 16313 24769 16347 24803
rect 21189 24769 21223 24803
rect 21465 24769 21499 24803
rect 22201 24769 22235 24803
rect 22385 24769 22419 24803
rect 23121 24769 23155 24803
rect 23765 24769 23799 24803
rect 24317 24769 24351 24803
rect 25412 24769 25446 24803
rect 27353 24769 27387 24803
rect 27629 24769 27663 24803
rect 31493 24769 31527 24803
rect 32321 24769 32355 24803
rect 32505 24769 32539 24803
rect 32781 24769 32815 24803
rect 32882 24769 32916 24803
rect 33609 24769 33643 24803
rect 33885 24769 33919 24803
rect 34069 24769 34103 24803
rect 35817 24769 35851 24803
rect 36001 24769 36035 24803
rect 36277 24769 36311 24803
rect 36737 24769 36771 24803
rect 36921 24769 36955 24803
rect 38209 24769 38243 24803
rect 47041 24769 47075 24803
rect 47133 24769 47167 24803
rect 48145 24769 48179 24803
rect 12817 24701 12851 24735
rect 18153 24701 18187 24735
rect 22477 24701 22511 24735
rect 24409 24701 24443 24735
rect 25145 24701 25179 24735
rect 29469 24701 29503 24735
rect 31677 24701 31711 24735
rect 31769 24701 31803 24735
rect 38485 24701 38519 24735
rect 15209 24633 15243 24667
rect 21189 24633 21223 24667
rect 26525 24633 26559 24667
rect 12725 24565 12759 24599
rect 15669 24565 15703 24599
rect 22017 24565 22051 24599
rect 23489 24565 23523 24599
rect 24501 24565 24535 24599
rect 24685 24565 24719 24599
rect 27169 24565 27203 24599
rect 27537 24565 27571 24599
rect 30849 24565 30883 24599
rect 33425 24565 33459 24599
rect 36737 24565 36771 24599
rect 38393 24565 38427 24599
rect 48237 24565 48271 24599
rect 14381 24361 14415 24395
rect 23213 24361 23247 24395
rect 23673 24361 23707 24395
rect 29837 24361 29871 24395
rect 14749 24293 14783 24327
rect 24593 24293 24627 24327
rect 25789 24293 25823 24327
rect 33701 24293 33735 24327
rect 25145 24225 25179 24259
rect 27077 24225 27111 24259
rect 40049 24225 40083 24259
rect 14565 24157 14599 24191
rect 14841 24157 14875 24191
rect 17141 24157 17175 24191
rect 18153 24157 18187 24191
rect 20637 24157 20671 24191
rect 20904 24157 20938 24191
rect 23121 24157 23155 24191
rect 23397 24157 23431 24191
rect 26065 24157 26099 24191
rect 27333 24157 27367 24191
rect 30021 24157 30055 24191
rect 30297 24157 30331 24191
rect 30481 24157 30515 24191
rect 32321 24157 32355 24191
rect 36369 24157 36403 24191
rect 36461 24157 36495 24191
rect 39497 24157 39531 24191
rect 18521 24089 18555 24123
rect 25789 24089 25823 24123
rect 25973 24089 26007 24123
rect 32588 24089 32622 24123
rect 40294 24089 40328 24123
rect 16957 24021 16991 24055
rect 22017 24021 22051 24055
rect 24961 24021 24995 24055
rect 25053 24021 25087 24055
rect 28457 24021 28491 24055
rect 36369 24021 36403 24055
rect 39313 24021 39347 24055
rect 41429 24021 41463 24055
rect 17509 23817 17543 23851
rect 25053 23817 25087 23851
rect 25697 23817 25731 23851
rect 27537 23817 27571 23851
rect 32597 23817 32631 23851
rect 39405 23817 39439 23851
rect 39773 23817 39807 23851
rect 39865 23817 39899 23851
rect 41153 23817 41187 23851
rect 11897 23749 11931 23783
rect 17049 23749 17083 23783
rect 18797 23749 18831 23783
rect 19809 23749 19843 23783
rect 24685 23749 24719 23783
rect 24869 23749 24903 23783
rect 17969 23681 18003 23715
rect 19993 23681 20027 23715
rect 22477 23681 22511 23715
rect 24133 23681 24167 23715
rect 25605 23681 25639 23715
rect 25789 23681 25823 23715
rect 27721 23681 27755 23715
rect 27997 23681 28031 23715
rect 28181 23681 28215 23715
rect 29561 23681 29595 23715
rect 29745 23681 29779 23715
rect 32781 23681 32815 23715
rect 33793 23681 33827 23715
rect 34049 23681 34083 23715
rect 36461 23681 36495 23715
rect 36645 23681 36679 23715
rect 40785 23681 40819 23715
rect 46305 23681 46339 23715
rect 29837 23613 29871 23647
rect 33057 23613 33091 23647
rect 39957 23613 39991 23647
rect 40693 23613 40727 23647
rect 17417 23545 17451 23579
rect 32965 23545 32999 23579
rect 12173 23477 12207 23511
rect 20177 23477 20211 23511
rect 22661 23477 22695 23511
rect 23949 23477 23983 23511
rect 24869 23477 24903 23511
rect 29377 23477 29411 23511
rect 35173 23477 35207 23511
rect 36553 23477 36587 23511
rect 46397 23477 46431 23511
rect 17693 23273 17727 23307
rect 18061 23273 18095 23307
rect 22753 23273 22787 23307
rect 24869 23273 24903 23307
rect 29745 23273 29779 23307
rect 40325 23273 40359 23307
rect 27629 23205 27663 23239
rect 11069 23137 11103 23171
rect 14289 23137 14323 23171
rect 18613 23137 18647 23171
rect 19441 23137 19475 23171
rect 39221 23137 39255 23171
rect 47593 23137 47627 23171
rect 10149 23069 10183 23103
rect 14565 23069 14599 23103
rect 16037 23069 16071 23103
rect 18521 23069 18555 23103
rect 21465 23069 21499 23103
rect 24685 23069 24719 23103
rect 27445 23069 27479 23103
rect 29929 23069 29963 23103
rect 30205 23069 30239 23103
rect 30389 23069 30423 23103
rect 33885 23069 33919 23103
rect 34161 23069 34195 23103
rect 34345 23069 34379 23103
rect 36369 23069 36403 23103
rect 36553 23069 36587 23103
rect 36645 23069 36679 23103
rect 37473 23069 37507 23103
rect 39129 23069 39163 23103
rect 39313 23069 39347 23103
rect 39405 23069 39439 23103
rect 40233 23069 40267 23103
rect 40417 23069 40451 23103
rect 45937 23069 45971 23103
rect 10333 23001 10367 23035
rect 16304 23001 16338 23035
rect 18429 23001 18463 23035
rect 19708 23001 19742 23035
rect 22569 23001 22603 23035
rect 22785 23001 22819 23035
rect 37105 23001 37139 23035
rect 37289 23001 37323 23035
rect 46121 23001 46155 23035
rect 17417 22933 17451 22967
rect 20821 22933 20855 22967
rect 21281 22933 21315 22967
rect 22937 22933 22971 22967
rect 33701 22933 33735 22967
rect 36185 22933 36219 22967
rect 38945 22933 38979 22967
rect 10517 22729 10551 22763
rect 18245 22729 18279 22763
rect 20177 22729 20211 22763
rect 20545 22729 20579 22763
rect 20637 22729 20671 22763
rect 33609 22729 33643 22763
rect 40509 22729 40543 22763
rect 46121 22729 46155 22763
rect 16865 22661 16899 22695
rect 22201 22661 22235 22695
rect 32505 22661 32539 22695
rect 38853 22661 38887 22695
rect 39497 22661 39531 22695
rect 40417 22661 40451 22695
rect 10425 22593 10459 22627
rect 12532 22593 12566 22627
rect 14197 22593 14231 22627
rect 14453 22593 14487 22627
rect 18153 22593 18187 22627
rect 23489 22593 23523 22627
rect 24501 22593 24535 22627
rect 29193 22593 29227 22627
rect 29460 22593 29494 22627
rect 31585 22593 31619 22627
rect 31769 22593 31803 22627
rect 32321 22593 32355 22627
rect 33793 22593 33827 22627
rect 34069 22593 34103 22627
rect 35817 22593 35851 22627
rect 36001 22593 36035 22627
rect 36369 22593 36403 22627
rect 38485 22593 38519 22627
rect 38669 22593 38703 22627
rect 39313 22593 39347 22627
rect 39589 22593 39623 22627
rect 39681 22593 39715 22627
rect 40325 22593 40359 22627
rect 40693 22593 40727 22627
rect 43085 22593 43119 22627
rect 43985 22593 44019 22627
rect 46029 22593 46063 22627
rect 12265 22525 12299 22559
rect 18429 22525 18463 22559
rect 20729 22525 20763 22559
rect 23765 22525 23799 22559
rect 33977 22525 34011 22559
rect 36093 22525 36127 22559
rect 36185 22525 36219 22559
rect 42901 22525 42935 22559
rect 43729 22525 43763 22559
rect 17233 22457 17267 22491
rect 17785 22457 17819 22491
rect 31677 22457 31711 22491
rect 39865 22457 39899 22491
rect 13645 22389 13679 22423
rect 15577 22389 15611 22423
rect 17325 22389 17359 22423
rect 22293 22389 22327 22423
rect 23581 22389 23615 22423
rect 24041 22389 24075 22423
rect 24593 22389 24627 22423
rect 30573 22389 30607 22423
rect 32689 22389 32723 22423
rect 36553 22389 36587 22423
rect 40417 22389 40451 22423
rect 41521 22389 41555 22423
rect 43269 22389 43303 22423
rect 45109 22389 45143 22423
rect 12357 22185 12391 22219
rect 14289 22185 14323 22219
rect 32781 22185 32815 22219
rect 38577 22185 38611 22219
rect 39497 22185 39531 22219
rect 40233 22185 40267 22219
rect 13553 22117 13587 22151
rect 20637 22117 20671 22151
rect 21189 22117 21223 22151
rect 33149 22117 33183 22151
rect 13277 22049 13311 22083
rect 15761 22049 15795 22083
rect 15853 22049 15887 22083
rect 20729 22049 20763 22083
rect 21741 22049 21775 22083
rect 33701 22049 33735 22083
rect 41337 22049 41371 22083
rect 44281 22049 44315 22083
rect 46397 22049 46431 22083
rect 46673 22049 46707 22083
rect 2237 21981 2271 22015
rect 12541 21981 12575 22015
rect 13185 21981 13219 22015
rect 14473 21981 14507 22015
rect 15669 21981 15703 22015
rect 17417 21981 17451 22015
rect 22569 21981 22603 22015
rect 23121 21981 23155 22015
rect 23305 21981 23339 22015
rect 24777 21981 24811 22015
rect 25053 21981 25087 22015
rect 25237 21981 25271 22015
rect 26801 21981 26835 22015
rect 27077 21981 27111 22015
rect 27261 21981 27295 22015
rect 30573 21981 30607 22015
rect 32965 21981 32999 22015
rect 33241 21981 33275 22015
rect 33885 21981 33919 22015
rect 34161 21981 34195 22015
rect 34345 21981 34379 22015
rect 36185 21981 36219 22015
rect 38485 21981 38519 22015
rect 38669 21981 38703 22015
rect 39221 21981 39255 22015
rect 39313 21981 39347 22015
rect 43177 21981 43211 22015
rect 45385 21981 45419 22015
rect 46213 21981 46247 22015
rect 17684 21913 17718 21947
rect 20269 21913 20303 21947
rect 25697 21913 25731 21947
rect 25881 21913 25915 21947
rect 30840 21913 30874 21947
rect 36452 21913 36486 21947
rect 40049 21913 40083 21947
rect 40249 21913 40283 21947
rect 41521 21913 41555 21947
rect 15301 21845 15335 21879
rect 18797 21845 18831 21879
rect 21557 21845 21591 21879
rect 21649 21845 21683 21879
rect 22385 21845 22419 21879
rect 23489 21845 23523 21879
rect 24593 21845 24627 21879
rect 26065 21845 26099 21879
rect 26617 21845 26651 21879
rect 31953 21845 31987 21879
rect 37565 21845 37599 21879
rect 40417 21845 40451 21879
rect 43637 21845 43671 21879
rect 44005 21845 44039 21879
rect 44097 21845 44131 21879
rect 45201 21845 45235 21879
rect 13277 21641 13311 21675
rect 13921 21641 13955 21675
rect 17785 21641 17819 21675
rect 21465 21641 21499 21675
rect 25237 21641 25271 21675
rect 31585 21641 31619 21675
rect 40877 21641 40911 21675
rect 42809 21641 42843 21675
rect 43729 21641 43763 21675
rect 45753 21641 45787 21675
rect 14381 21573 14415 21607
rect 15945 21573 15979 21607
rect 24124 21573 24158 21607
rect 33968 21573 34002 21607
rect 39865 21573 39899 21607
rect 44640 21573 44674 21607
rect 2053 21505 2087 21539
rect 9597 21505 9631 21539
rect 10425 21505 10459 21539
rect 12164 21505 12198 21539
rect 14289 21505 14323 21539
rect 17969 21505 18003 21539
rect 20085 21505 20119 21539
rect 20352 21505 20386 21539
rect 23121 21505 23155 21539
rect 23857 21505 23891 21539
rect 25881 21505 25915 21539
rect 26249 21505 26283 21539
rect 27169 21505 27203 21539
rect 27425 21505 27459 21539
rect 29016 21505 29050 21539
rect 29265 21505 29299 21539
rect 30849 21505 30883 21539
rect 31033 21505 31067 21539
rect 31125 21505 31159 21539
rect 31401 21505 31435 21539
rect 32965 21505 32999 21539
rect 33149 21505 33183 21539
rect 33241 21505 33275 21539
rect 33701 21505 33735 21539
rect 39596 21505 39630 21539
rect 39737 21505 39771 21539
rect 39957 21505 39991 21539
rect 40095 21505 40129 21539
rect 40785 21505 40819 21539
rect 42993 21505 43027 21539
rect 43177 21505 43211 21539
rect 43269 21505 43303 21539
rect 43913 21505 43947 21539
rect 44373 21505 44407 21539
rect 47041 21505 47075 21539
rect 2237 21437 2271 21471
rect 2789 21437 2823 21471
rect 9689 21437 9723 21471
rect 11897 21437 11931 21471
rect 14473 21437 14507 21471
rect 16037 21437 16071 21471
rect 16129 21437 16163 21471
rect 26433 21437 26467 21471
rect 31217 21437 31251 21471
rect 9965 21369 9999 21403
rect 32781 21369 32815 21403
rect 35081 21369 35115 21403
rect 10517 21301 10551 21335
rect 15577 21301 15611 21335
rect 23305 21301 23339 21335
rect 28549 21301 28583 21335
rect 30389 21301 30423 21335
rect 40233 21301 40267 21335
rect 47133 21301 47167 21335
rect 47961 21301 47995 21335
rect 2329 21097 2363 21131
rect 12817 21097 12851 21131
rect 16681 21097 16715 21131
rect 24593 21097 24627 21131
rect 27169 21097 27203 21131
rect 28917 21097 28951 21131
rect 34069 21097 34103 21131
rect 41429 21097 41463 21131
rect 42809 21097 42843 21131
rect 43453 21097 43487 21131
rect 43637 21097 43671 21131
rect 10241 20961 10275 20995
rect 10517 20961 10551 20995
rect 13277 20961 13311 20995
rect 13369 20961 13403 20995
rect 23857 20961 23891 20995
rect 42625 20961 42659 20995
rect 44189 20961 44223 20995
rect 46489 20961 46523 20995
rect 46673 20961 46707 20995
rect 48237 20961 48271 20995
rect 2237 20893 2271 20927
rect 4537 20893 4571 20927
rect 10057 20893 10091 20927
rect 15301 20893 15335 20927
rect 19993 20893 20027 20927
rect 24869 20893 24903 20927
rect 24961 20893 24995 20927
rect 25053 20893 25087 20927
rect 25237 20893 25271 20927
rect 26157 20893 26191 20927
rect 28181 20893 28215 20927
rect 28365 20893 28399 20927
rect 28457 20893 28491 20927
rect 28549 20893 28583 20927
rect 28733 20893 28767 20927
rect 32689 20893 32723 20927
rect 32873 20893 32907 20927
rect 33701 20893 33735 20927
rect 37841 20893 37875 20927
rect 38117 20893 38151 20927
rect 38301 20893 38335 20927
rect 40049 20893 40083 20927
rect 40316 20893 40350 20927
rect 42441 20893 42475 20927
rect 42809 20893 42843 20927
rect 44373 20893 44407 20927
rect 15546 20825 15580 20859
rect 23121 20825 23155 20859
rect 27077 20825 27111 20859
rect 32781 20825 32815 20859
rect 33885 20825 33919 20859
rect 42533 20825 42567 20859
rect 43269 20825 43303 20859
rect 13185 20757 13219 20791
rect 19809 20757 19843 20791
rect 26433 20757 26467 20791
rect 37657 20757 37691 20791
rect 43469 20757 43503 20791
rect 44557 20757 44591 20791
rect 12449 20553 12483 20587
rect 15301 20553 15335 20587
rect 24609 20553 24643 20587
rect 24777 20553 24811 20587
rect 27169 20553 27203 20587
rect 29193 20553 29227 20587
rect 33793 20553 33827 20587
rect 19594 20485 19628 20519
rect 24409 20485 24443 20519
rect 25329 20485 25363 20519
rect 28365 20485 28399 20519
rect 4169 20417 4203 20451
rect 10057 20417 10091 20451
rect 12633 20417 12667 20451
rect 18429 20417 18463 20451
rect 23397 20417 23431 20451
rect 23673 20417 23707 20451
rect 27353 20417 27387 20451
rect 27629 20417 27663 20451
rect 28181 20417 28215 20451
rect 29009 20417 29043 20451
rect 29193 20417 29227 20451
rect 29653 20417 29687 20451
rect 29837 20417 29871 20451
rect 31033 20417 31067 20451
rect 31217 20417 31251 20451
rect 33701 20417 33735 20451
rect 33885 20417 33919 20451
rect 34345 20417 34379 20451
rect 34529 20417 34563 20451
rect 37473 20417 37507 20451
rect 37740 20417 37774 20451
rect 40325 20417 40359 20451
rect 40785 20417 40819 20451
rect 46765 20417 46799 20451
rect 4353 20349 4387 20383
rect 4997 20349 5031 20383
rect 10149 20349 10183 20383
rect 10425 20349 10459 20383
rect 15393 20349 15427 20383
rect 15577 20349 15611 20383
rect 19349 20349 19383 20383
rect 23765 20349 23799 20383
rect 28549 20349 28583 20383
rect 31309 20349 31343 20383
rect 40877 20349 40911 20383
rect 20729 20281 20763 20315
rect 14933 20213 14967 20247
rect 18245 20213 18279 20247
rect 24593 20213 24627 20247
rect 25421 20213 25455 20247
rect 27537 20213 27571 20247
rect 29745 20213 29779 20247
rect 30849 20213 30883 20247
rect 34437 20213 34471 20247
rect 38853 20213 38887 20247
rect 46857 20213 46891 20247
rect 47961 20213 47995 20247
rect 4905 20009 4939 20043
rect 15209 20009 15243 20043
rect 22569 20009 22603 20043
rect 28273 20009 28307 20043
rect 34161 20009 34195 20043
rect 37749 20009 37783 20043
rect 40417 20009 40451 20043
rect 10701 19873 10735 19907
rect 18705 19873 18739 19907
rect 20821 19873 20855 19907
rect 30665 19873 30699 19907
rect 34253 19873 34287 19907
rect 35173 19873 35207 19907
rect 38209 19873 38243 19907
rect 41889 19873 41923 19907
rect 44189 19873 44223 19907
rect 46489 19873 46523 19907
rect 46673 19873 46707 19907
rect 48237 19873 48271 19907
rect 4813 19805 4847 19839
rect 9597 19805 9631 19839
rect 10241 19805 10275 19839
rect 15393 19805 15427 19839
rect 16037 19805 16071 19839
rect 17969 19805 18003 19839
rect 20637 19805 20671 19839
rect 22385 19805 22419 19839
rect 22661 19805 22695 19839
rect 23397 19805 23431 19839
rect 23581 19805 23615 19839
rect 28457 19805 28491 19839
rect 28733 19805 28767 19839
rect 30932 19805 30966 19839
rect 32505 19805 32539 19839
rect 33977 19805 34011 19839
rect 35081 19805 35115 19839
rect 35909 19805 35943 19839
rect 37933 19805 37967 19839
rect 38117 19805 38151 19839
rect 40141 19805 40175 19839
rect 42165 19805 42199 19839
rect 44005 19805 44039 19839
rect 44373 19805 44407 19839
rect 9689 19737 9723 19771
rect 10425 19737 10459 19771
rect 20729 19737 20763 19771
rect 23765 19737 23799 19771
rect 24685 19737 24719 19771
rect 24869 19737 24903 19771
rect 32689 19737 32723 19771
rect 33793 19737 33827 19771
rect 36154 19737 36188 19771
rect 44097 19737 44131 19771
rect 15853 19669 15887 19703
rect 20269 19669 20303 19703
rect 22201 19669 22235 19703
rect 28641 19669 28675 19703
rect 32045 19669 32079 19703
rect 32873 19669 32907 19703
rect 35449 19669 35483 19703
rect 37289 19669 37323 19703
rect 43269 19669 43303 19703
rect 44281 19669 44315 19703
rect 13093 19465 13127 19499
rect 18245 19465 18279 19499
rect 19073 19465 19107 19499
rect 20177 19465 20211 19499
rect 28089 19465 28123 19499
rect 28917 19465 28951 19499
rect 29469 19465 29503 19499
rect 31033 19465 31067 19499
rect 35909 19465 35943 19499
rect 36553 19465 36587 19499
rect 40141 19465 40175 19499
rect 43545 19465 43579 19499
rect 44649 19465 44683 19499
rect 17785 19397 17819 19431
rect 18705 19397 18739 19431
rect 18889 19397 18923 19431
rect 19717 19397 19751 19431
rect 22753 19397 22787 19431
rect 37473 19397 37507 19431
rect 37657 19397 37691 19431
rect 43729 19397 43763 19431
rect 9965 19329 9999 19363
rect 11713 19329 11747 19363
rect 11969 19329 12003 19363
rect 13921 19329 13955 19363
rect 14933 19329 14967 19363
rect 17877 19329 17911 19363
rect 22937 19329 22971 19363
rect 23213 19329 23247 19363
rect 23397 19329 23431 19363
rect 24409 19329 24443 19363
rect 25237 19329 25271 19363
rect 25504 19329 25538 19363
rect 27169 19329 27203 19363
rect 27353 19329 27387 19363
rect 27813 19329 27847 19363
rect 28549 19329 28583 19363
rect 28733 19329 28767 19363
rect 29377 19329 29411 19363
rect 29561 19329 29595 19363
rect 31217 19329 31251 19363
rect 31493 19329 31527 19363
rect 31677 19329 31711 19363
rect 33885 19329 33919 19363
rect 34253 19329 34287 19363
rect 35173 19329 35207 19363
rect 35357 19329 35391 19363
rect 35725 19329 35759 19363
rect 36461 19329 36495 19363
rect 36645 19329 36679 19363
rect 39957 19329 39991 19363
rect 41889 19329 41923 19363
rect 41981 19329 42015 19363
rect 43361 19329 43395 19363
rect 43821 19329 43855 19363
rect 44465 19329 44499 19363
rect 44741 19329 44775 19363
rect 47041 19329 47075 19363
rect 10057 19261 10091 19295
rect 10333 19261 10367 19295
rect 14013 19261 14047 19295
rect 14841 19261 14875 19295
rect 17693 19261 17727 19295
rect 28089 19261 28123 19295
rect 33793 19261 33827 19295
rect 35449 19261 35483 19295
rect 35541 19261 35575 19295
rect 39773 19261 39807 19295
rect 43453 19261 43487 19295
rect 15301 19193 15335 19227
rect 17233 19193 17267 19227
rect 20085 19193 20119 19227
rect 26617 19193 26651 19227
rect 14197 19125 14231 19159
rect 24685 19125 24719 19159
rect 27169 19125 27203 19159
rect 27905 19125 27939 19159
rect 34161 19125 34195 19159
rect 34437 19125 34471 19159
rect 37841 19125 37875 19159
rect 43177 19125 43211 19159
rect 44281 19125 44315 19159
rect 47133 19125 47167 19159
rect 47961 19125 47995 19159
rect 11713 18921 11747 18955
rect 23213 18921 23247 18955
rect 26801 18921 26835 18955
rect 28365 18921 28399 18955
rect 28733 18921 28767 18955
rect 31401 18921 31435 18955
rect 35265 18921 35299 18955
rect 39037 18921 39071 18955
rect 42625 18921 42659 18955
rect 13001 18853 13035 18887
rect 24961 18853 24995 18887
rect 12725 18785 12759 18819
rect 26341 18785 26375 18819
rect 42993 18785 43027 18819
rect 46489 18785 46523 18819
rect 46673 18785 46707 18819
rect 48237 18785 48271 18819
rect 2237 18717 2271 18751
rect 11897 18717 11931 18751
rect 12633 18717 12667 18751
rect 14933 18717 14967 18751
rect 15200 18717 15234 18751
rect 16957 18717 16991 18751
rect 21833 18717 21867 18751
rect 24777 18717 24811 18751
rect 25053 18717 25087 18751
rect 26065 18717 26099 18751
rect 26249 18717 26283 18751
rect 26433 18717 26467 18751
rect 26617 18717 26651 18751
rect 27537 18717 27571 18751
rect 27813 18717 27847 18751
rect 28273 18717 28307 18751
rect 30297 18717 30331 18751
rect 30481 18717 30515 18751
rect 30573 18717 30607 18751
rect 33885 18717 33919 18751
rect 33977 18717 34011 18751
rect 34989 18717 35023 18751
rect 35081 18717 35115 18751
rect 35725 18717 35759 18751
rect 35909 18717 35943 18751
rect 38853 18717 38887 18751
rect 39129 18717 39163 18751
rect 40785 18717 40819 18751
rect 42809 18717 42843 18751
rect 42901 18717 42935 18751
rect 43085 18717 43119 18751
rect 44097 18717 44131 18751
rect 44281 18717 44315 18751
rect 44373 18717 44407 18751
rect 44465 18717 44499 18751
rect 17224 18649 17258 18683
rect 22100 18649 22134 18683
rect 31125 18649 31159 18683
rect 33701 18649 33735 18683
rect 41153 18649 41187 18683
rect 16313 18581 16347 18615
rect 18337 18581 18371 18615
rect 24593 18581 24627 18615
rect 27353 18581 27387 18615
rect 27721 18581 27755 18615
rect 30113 18581 30147 18615
rect 33977 18581 34011 18615
rect 35909 18581 35943 18615
rect 38669 18581 38703 18615
rect 44649 18581 44683 18615
rect 12265 18377 12299 18411
rect 15945 18377 15979 18411
rect 22293 18377 22327 18411
rect 36645 18377 36679 18411
rect 38485 18377 38519 18411
rect 41797 18377 41831 18411
rect 43653 18377 43687 18411
rect 43821 18377 43855 18411
rect 46213 18377 46247 18411
rect 12633 18309 12667 18343
rect 23664 18309 23698 18343
rect 26525 18309 26559 18343
rect 30634 18309 30668 18343
rect 33793 18309 33827 18343
rect 37657 18309 37691 18343
rect 42717 18309 42751 18343
rect 43453 18309 43487 18343
rect 45078 18309 45112 18343
rect 34023 18275 34057 18309
rect 2053 18241 2087 18275
rect 19073 18241 19107 18275
rect 22477 18241 22511 18275
rect 22753 18241 22787 18275
rect 22937 18241 22971 18275
rect 26433 18241 26467 18275
rect 26617 18241 26651 18275
rect 27721 18241 27755 18275
rect 27905 18241 27939 18275
rect 27997 18241 28031 18275
rect 28549 18241 28583 18275
rect 28641 18241 28675 18275
rect 30389 18241 30423 18275
rect 33241 18241 33275 18275
rect 36461 18241 36495 18275
rect 36737 18241 36771 18275
rect 37473 18241 37507 18275
rect 37749 18241 37783 18275
rect 37877 18241 37911 18275
rect 38669 18241 38703 18275
rect 38945 18241 38979 18275
rect 39129 18241 39163 18275
rect 40684 18241 40718 18275
rect 42625 18241 42659 18275
rect 42993 18241 43027 18275
rect 44833 18241 44867 18275
rect 46765 18241 46799 18275
rect 47777 18241 47811 18275
rect 2237 18173 2271 18207
rect 2789 18173 2823 18207
rect 12725 18173 12759 18207
rect 12909 18173 12943 18207
rect 16037 18173 16071 18207
rect 16129 18173 16163 18207
rect 19165 18173 19199 18207
rect 19257 18173 19291 18207
rect 23397 18173 23431 18207
rect 32965 18173 32999 18207
rect 33057 18173 33091 18207
rect 33149 18173 33183 18207
rect 40417 18173 40451 18207
rect 42809 18173 42843 18207
rect 24777 18105 24811 18139
rect 27813 18105 27847 18139
rect 28917 18105 28951 18139
rect 31769 18105 31803 18139
rect 34161 18105 34195 18139
rect 47869 18105 47903 18139
rect 15577 18037 15611 18071
rect 18705 18037 18739 18071
rect 27537 18037 27571 18071
rect 28733 18037 28767 18071
rect 32781 18037 32815 18071
rect 33977 18037 34011 18071
rect 36461 18037 36495 18071
rect 37473 18037 37507 18071
rect 42993 18037 43027 18071
rect 43637 18037 43671 18071
rect 46857 18037 46891 18071
rect 2329 17833 2363 17867
rect 12909 17833 12943 17867
rect 23581 17833 23615 17867
rect 28825 17833 28859 17867
rect 30849 17833 30883 17867
rect 39497 17833 39531 17867
rect 40877 17833 40911 17867
rect 44189 17833 44223 17867
rect 18705 17765 18739 17799
rect 28273 17765 28307 17799
rect 44373 17765 44407 17799
rect 11529 17697 11563 17731
rect 18797 17697 18831 17731
rect 28181 17697 28215 17731
rect 28365 17697 28399 17731
rect 37013 17697 37047 17731
rect 37105 17697 37139 17731
rect 43453 17697 43487 17731
rect 46489 17697 46523 17731
rect 46673 17697 46707 17731
rect 48053 17697 48087 17731
rect 2237 17629 2271 17663
rect 15209 17629 15243 17663
rect 18337 17629 18371 17663
rect 19625 17629 19659 17663
rect 22017 17629 22051 17663
rect 23489 17629 23523 17663
rect 28089 17629 28123 17663
rect 29101 17629 29135 17663
rect 31033 17629 31067 17663
rect 31309 17629 31343 17663
rect 31493 17629 31527 17663
rect 35541 17629 35575 17663
rect 35633 17629 35667 17663
rect 36001 17629 36035 17663
rect 36921 17629 36955 17663
rect 37197 17629 37231 17663
rect 38117 17629 38151 17663
rect 38384 17629 38418 17663
rect 41061 17629 41095 17663
rect 41705 17629 41739 17663
rect 41889 17629 41923 17663
rect 41981 17629 42015 17663
rect 43177 17629 43211 17663
rect 11796 17561 11830 17595
rect 22753 17561 22787 17595
rect 28825 17561 28859 17595
rect 35725 17561 35759 17595
rect 35843 17561 35877 17595
rect 44005 17561 44039 17595
rect 15025 17493 15059 17527
rect 19441 17493 19475 17527
rect 29009 17493 29043 17527
rect 35357 17493 35391 17527
rect 36737 17493 36771 17527
rect 41521 17493 41555 17527
rect 42809 17493 42843 17527
rect 43269 17493 43303 17527
rect 44205 17493 44239 17527
rect 12081 17289 12115 17323
rect 19809 17289 19843 17323
rect 26249 17289 26283 17323
rect 35817 17289 35851 17323
rect 41797 17289 41831 17323
rect 44925 17289 44959 17323
rect 14556 17221 14590 17255
rect 18696 17221 18730 17255
rect 23296 17221 23330 17255
rect 33885 17221 33919 17255
rect 34621 17221 34655 17255
rect 34821 17221 34855 17255
rect 35449 17221 35483 17255
rect 35649 17221 35683 17255
rect 39405 17221 39439 17255
rect 45569 17221 45603 17255
rect 12265 17153 12299 17187
rect 13461 17153 13495 17187
rect 14289 17153 14323 17187
rect 17049 17153 17083 17187
rect 22201 17153 22235 17187
rect 22477 17153 22511 17187
rect 25237 17153 25271 17187
rect 26157 17153 26191 17187
rect 31033 17153 31067 17187
rect 31309 17153 31343 17187
rect 31493 17153 31527 17187
rect 34069 17153 34103 17187
rect 34161 17153 34195 17187
rect 36553 17153 36587 17187
rect 37729 17153 37763 17187
rect 39313 17153 39347 17187
rect 39497 17153 39531 17187
rect 41613 17153 41647 17187
rect 42717 17153 42751 17187
rect 43545 17153 43579 17187
rect 43801 17153 43835 17187
rect 13553 17085 13587 17119
rect 13829 17085 13863 17119
rect 18429 17085 18463 17119
rect 23029 17085 23063 17119
rect 25329 17085 25363 17119
rect 25513 17085 25547 17119
rect 36645 17085 36679 17119
rect 36921 17085 36955 17119
rect 37473 17085 37507 17119
rect 41429 17085 41463 17119
rect 45385 17085 45419 17119
rect 46857 17085 46891 17119
rect 33885 17017 33919 17051
rect 2329 16949 2363 16983
rect 15669 16949 15703 16983
rect 16865 16949 16899 16983
rect 22017 16949 22051 16983
rect 22385 16949 22419 16983
rect 24409 16949 24443 16983
rect 24869 16949 24903 16983
rect 30849 16949 30883 16983
rect 34805 16949 34839 16983
rect 34989 16949 35023 16983
rect 35633 16949 35667 16983
rect 38853 16949 38887 16983
rect 42993 16949 43027 16983
rect 47961 16949 47995 16983
rect 12725 16745 12759 16779
rect 23489 16745 23523 16779
rect 26249 16745 26283 16779
rect 27813 16745 27847 16779
rect 35265 16745 35299 16779
rect 36737 16745 36771 16779
rect 36829 16745 36863 16779
rect 43453 16745 43487 16779
rect 38301 16677 38335 16711
rect 1593 16609 1627 16643
rect 2789 16609 2823 16643
rect 13185 16609 13219 16643
rect 13369 16609 13403 16643
rect 16405 16609 16439 16643
rect 20821 16609 20855 16643
rect 25053 16609 25087 16643
rect 25237 16609 25271 16643
rect 26893 16609 26927 16643
rect 27905 16609 27939 16643
rect 30297 16609 30331 16643
rect 32137 16609 32171 16643
rect 36921 16609 36955 16643
rect 46489 16609 46523 16643
rect 48237 16609 48271 16643
rect 21088 16541 21122 16575
rect 23673 16541 23707 16575
rect 25881 16541 25915 16575
rect 27077 16541 27111 16575
rect 27261 16541 27295 16575
rect 27353 16541 27387 16575
rect 27813 16541 27847 16575
rect 34069 16541 34103 16575
rect 34345 16541 34379 16575
rect 35725 16541 35759 16575
rect 35909 16541 35943 16575
rect 36645 16541 36679 16575
rect 38025 16541 38059 16575
rect 43637 16541 43671 16575
rect 1777 16473 1811 16507
rect 16672 16473 16706 16507
rect 26065 16473 26099 16507
rect 30564 16473 30598 16507
rect 32404 16473 32438 16507
rect 34253 16473 34287 16507
rect 34897 16473 34931 16507
rect 35081 16473 35115 16507
rect 35817 16473 35851 16507
rect 46673 16473 46707 16507
rect 13093 16405 13127 16439
rect 17785 16405 17819 16439
rect 22201 16405 22235 16439
rect 24593 16405 24627 16439
rect 24961 16405 24995 16439
rect 28181 16405 28215 16439
rect 31677 16405 31711 16439
rect 33517 16405 33551 16439
rect 34167 16405 34201 16439
rect 2605 16201 2639 16235
rect 13461 16201 13495 16235
rect 17141 16201 17175 16235
rect 17509 16201 17543 16235
rect 18705 16201 18739 16235
rect 22017 16201 22051 16235
rect 26249 16201 26283 16235
rect 32321 16201 32355 16235
rect 34923 16201 34957 16235
rect 42825 16201 42859 16235
rect 47133 16201 47167 16235
rect 14749 16133 14783 16167
rect 18337 16133 18371 16167
rect 25145 16133 25179 16167
rect 34713 16133 34747 16167
rect 42625 16133 42659 16167
rect 2513 16065 2547 16099
rect 12081 16065 12115 16099
rect 12348 16065 12382 16099
rect 14841 16065 14875 16099
rect 18521 16065 18555 16099
rect 19349 16065 19383 16099
rect 22201 16065 22235 16099
rect 22477 16065 22511 16099
rect 22661 16065 22695 16099
rect 24409 16065 24443 16099
rect 24593 16065 24627 16099
rect 25053 16065 25087 16099
rect 25237 16065 25271 16099
rect 25881 16065 25915 16099
rect 27261 16065 27295 16099
rect 27445 16065 27479 16099
rect 27537 16065 27571 16099
rect 27813 16065 27847 16099
rect 31033 16065 31067 16099
rect 31309 16065 31343 16099
rect 31493 16065 31527 16099
rect 32505 16065 32539 16099
rect 32689 16065 32723 16099
rect 32781 16065 32815 16099
rect 33425 16065 33459 16099
rect 33609 16065 33643 16099
rect 35541 16065 35575 16099
rect 40029 16065 40063 16099
rect 41613 16065 41647 16099
rect 41797 16065 41831 16099
rect 47041 16065 47075 16099
rect 14933 15997 14967 16031
rect 17601 15997 17635 16031
rect 17693 15997 17727 16031
rect 25973 15997 26007 16031
rect 27629 15997 27663 16031
rect 27997 15997 28031 16031
rect 33701 15997 33735 16031
rect 35817 15997 35851 16031
rect 39773 15997 39807 16031
rect 47961 15997 47995 16031
rect 41153 15929 41187 15963
rect 42993 15929 43027 15963
rect 14381 15861 14415 15895
rect 19165 15861 19199 15895
rect 24409 15861 24443 15895
rect 30849 15861 30883 15895
rect 33241 15861 33275 15895
rect 34897 15861 34931 15895
rect 35081 15861 35115 15895
rect 35633 15861 35667 15895
rect 35725 15861 35759 15895
rect 41705 15861 41739 15895
rect 42809 15861 42843 15895
rect 12909 15657 12943 15691
rect 18889 15657 18923 15691
rect 26249 15657 26283 15691
rect 30481 15657 30515 15691
rect 30849 15657 30883 15691
rect 39313 15657 39347 15691
rect 28089 15589 28123 15623
rect 2789 15521 2823 15555
rect 15025 15521 15059 15555
rect 15117 15521 15151 15555
rect 17693 15521 17727 15555
rect 19993 15521 20027 15555
rect 22661 15521 22695 15555
rect 25789 15521 25823 15555
rect 27629 15521 27663 15555
rect 30941 15521 30975 15555
rect 40785 15521 40819 15555
rect 41797 15521 41831 15555
rect 41889 15521 41923 15555
rect 42717 15521 42751 15555
rect 46489 15521 46523 15555
rect 48237 15521 48271 15555
rect 1593 15453 1627 15487
rect 13093 15453 13127 15487
rect 13737 15453 13771 15487
rect 17417 15453 17451 15487
rect 19809 15453 19843 15487
rect 19901 15453 19935 15487
rect 25421 15453 25455 15487
rect 25605 15453 25639 15487
rect 26249 15453 26283 15487
rect 26433 15453 26467 15487
rect 26893 15453 26927 15487
rect 27077 15453 27111 15487
rect 27721 15453 27755 15487
rect 28549 15453 28583 15487
rect 28733 15453 28767 15487
rect 30665 15453 30699 15487
rect 34897 15453 34931 15487
rect 35081 15453 35115 15487
rect 35265 15453 35299 15487
rect 37381 15453 37415 15487
rect 37657 15453 37691 15487
rect 39497 15453 39531 15487
rect 41613 15453 41647 15487
rect 41705 15453 41739 15487
rect 1777 15385 1811 15419
rect 14933 15385 14967 15419
rect 18521 15385 18555 15419
rect 18705 15385 18739 15419
rect 22928 15385 22962 15419
rect 26985 15385 27019 15419
rect 35173 15385 35207 15419
rect 40049 15385 40083 15419
rect 42984 15385 43018 15419
rect 46673 15385 46707 15419
rect 13553 15317 13587 15351
rect 14565 15317 14599 15351
rect 17049 15317 17083 15351
rect 17509 15317 17543 15351
rect 19441 15317 19475 15351
rect 24041 15317 24075 15351
rect 28641 15317 28675 15351
rect 35449 15317 35483 15351
rect 37197 15317 37231 15351
rect 37565 15317 37599 15351
rect 41429 15317 41463 15351
rect 44097 15317 44131 15351
rect 2881 15113 2915 15147
rect 15209 15113 15243 15147
rect 17325 15113 17359 15147
rect 19901 15113 19935 15147
rect 27261 15113 27295 15147
rect 35725 15113 35759 15147
rect 40351 15113 40385 15147
rect 43085 15113 43119 15147
rect 47133 15113 47167 15147
rect 14096 15045 14130 15079
rect 16865 15045 16899 15079
rect 18788 15045 18822 15079
rect 34612 15045 34646 15079
rect 37718 15045 37752 15079
rect 40141 15045 40175 15079
rect 43571 15045 43605 15079
rect 2329 14977 2363 15011
rect 2789 14977 2823 15011
rect 3801 14977 3835 15011
rect 13829 14977 13863 15011
rect 16313 14977 16347 15011
rect 18521 14977 18555 15011
rect 23397 14977 23431 15011
rect 23673 14977 23707 15011
rect 23857 14977 23891 15011
rect 27169 14977 27203 15011
rect 27353 14977 27387 15011
rect 28733 14977 28767 15011
rect 29000 14977 29034 15011
rect 32689 14977 32723 15011
rect 32873 14977 32907 15011
rect 37473 14977 37507 15011
rect 43269 14977 43303 15011
rect 43361 14977 43395 15011
rect 43453 14977 43487 15011
rect 43729 14977 43763 15011
rect 44189 14977 44223 15011
rect 47041 14977 47075 15011
rect 47961 14977 47995 15011
rect 3985 14909 4019 14943
rect 5365 14909 5399 14943
rect 32965 14909 32999 14943
rect 34345 14909 34379 14943
rect 44465 14909 44499 14943
rect 17141 14841 17175 14875
rect 16129 14773 16163 14807
rect 23213 14773 23247 14807
rect 30113 14773 30147 14807
rect 32505 14773 32539 14807
rect 38853 14773 38887 14807
rect 40325 14773 40359 14807
rect 40509 14773 40543 14807
rect 44281 14773 44315 14807
rect 44373 14773 44407 14807
rect 4077 14569 4111 14603
rect 17417 14569 17451 14603
rect 23213 14569 23247 14603
rect 23581 14569 23615 14603
rect 25053 14569 25087 14603
rect 26709 14569 26743 14603
rect 29193 14569 29227 14603
rect 38945 14569 38979 14603
rect 41153 14569 41187 14603
rect 44281 14569 44315 14603
rect 44649 14569 44683 14603
rect 30113 14501 30147 14535
rect 2789 14433 2823 14467
rect 23673 14433 23707 14467
rect 27537 14433 27571 14467
rect 33701 14433 33735 14467
rect 43545 14433 43579 14467
rect 43821 14433 43855 14467
rect 44373 14433 44407 14467
rect 1593 14365 1627 14399
rect 3985 14365 4019 14399
rect 16037 14365 16071 14399
rect 23397 14365 23431 14399
rect 24869 14365 24903 14399
rect 25145 14365 25179 14399
rect 26525 14365 26559 14399
rect 27353 14365 27387 14399
rect 27629 14365 27663 14399
rect 28549 14365 28583 14399
rect 28697 14365 28731 14399
rect 29055 14365 29089 14399
rect 29929 14365 29963 14399
rect 30185 14365 30219 14399
rect 31493 14365 31527 14399
rect 31769 14365 31803 14399
rect 31861 14365 31895 14399
rect 32965 14365 32999 14399
rect 37933 14365 37967 14399
rect 38301 14365 38335 14399
rect 38761 14365 38795 14399
rect 40969 14365 41003 14399
rect 43453 14365 43487 14399
rect 44281 14365 44315 14399
rect 1777 14297 1811 14331
rect 16282 14297 16316 14331
rect 26341 14297 26375 14331
rect 28825 14297 28859 14331
rect 28917 14297 28951 14331
rect 31677 14297 31711 14331
rect 40785 14297 40819 14331
rect 24685 14229 24719 14263
rect 27169 14229 27203 14263
rect 29745 14229 29779 14263
rect 32045 14229 32079 14263
rect 2881 14025 2915 14059
rect 25697 14025 25731 14059
rect 28549 14025 28583 14059
rect 31125 14025 31159 14059
rect 38853 14025 38887 14059
rect 40785 14025 40819 14059
rect 44649 14025 44683 14059
rect 46581 14025 46615 14059
rect 30012 13957 30046 13991
rect 32588 13957 32622 13991
rect 2329 13889 2363 13923
rect 2789 13889 2823 13923
rect 21189 13889 21223 13923
rect 22017 13889 22051 13923
rect 22201 13889 22235 13923
rect 22477 13889 22511 13923
rect 22661 13889 22695 13923
rect 24317 13889 24351 13923
rect 24584 13889 24618 13923
rect 26157 13889 26191 13923
rect 26341 13889 26375 13923
rect 27169 13889 27203 13923
rect 27425 13889 27459 13923
rect 29745 13889 29779 13923
rect 37473 13889 37507 13923
rect 37729 13889 37763 13923
rect 39405 13889 39439 13923
rect 39672 13889 39706 13923
rect 41245 13889 41279 13923
rect 41429 13889 41463 13923
rect 41613 13889 41647 13923
rect 41705 13889 41739 13923
rect 43545 13889 43579 13923
rect 43729 13889 43763 13923
rect 43821 13889 43855 13923
rect 44465 13889 44499 13923
rect 45468 13889 45502 13923
rect 47041 13889 47075 13923
rect 21373 13821 21407 13855
rect 21465 13821 21499 13855
rect 26525 13821 26559 13855
rect 32321 13821 32355 13855
rect 44281 13821 44315 13855
rect 45201 13821 45235 13855
rect 21005 13685 21039 13719
rect 33701 13685 33735 13719
rect 43361 13685 43395 13719
rect 47133 13685 47167 13719
rect 47961 13685 47995 13719
rect 22201 13481 22235 13515
rect 23029 13481 23063 13515
rect 24777 13481 24811 13515
rect 27629 13481 27663 13515
rect 30389 13481 30423 13515
rect 32229 13481 32263 13515
rect 33701 13481 33735 13515
rect 37565 13481 37599 13515
rect 45753 13481 45787 13515
rect 23121 13345 23155 13379
rect 40877 13345 40911 13379
rect 46489 13345 46523 13379
rect 46673 13345 46707 13379
rect 48237 13345 48271 13379
rect 20821 13277 20855 13311
rect 21088 13277 21122 13311
rect 22845 13277 22879 13311
rect 24961 13277 24995 13311
rect 25237 13277 25271 13311
rect 25421 13277 25455 13311
rect 27813 13277 27847 13311
rect 28089 13277 28123 13311
rect 28273 13277 28307 13311
rect 30573 13277 30607 13311
rect 30849 13277 30883 13311
rect 31033 13277 31067 13311
rect 32413 13277 32447 13311
rect 32689 13277 32723 13311
rect 32873 13277 32907 13311
rect 33517 13277 33551 13311
rect 33793 13277 33827 13311
rect 37013 13277 37047 13311
rect 37381 13277 37415 13311
rect 38025 13277 38059 13311
rect 38209 13277 38243 13311
rect 40141 13277 40175 13311
rect 41521 13277 41555 13311
rect 41705 13277 41739 13311
rect 41797 13277 41831 13311
rect 42257 13277 42291 13311
rect 42441 13277 42475 13311
rect 43545 13277 43579 13311
rect 43729 13277 43763 13311
rect 44189 13277 44223 13311
rect 44373 13277 44407 13311
rect 45201 13277 45235 13311
rect 45477 13277 45511 13311
rect 45569 13277 45603 13311
rect 37197 13209 37231 13243
rect 37289 13209 37323 13243
rect 42349 13209 42383 13243
rect 43637 13209 43671 13243
rect 45385 13209 45419 13243
rect 22661 13141 22695 13175
rect 33333 13141 33367 13175
rect 38393 13141 38427 13175
rect 41613 13141 41647 13175
rect 44281 13141 44315 13175
rect 22017 12937 22051 12971
rect 40049 12937 40083 12971
rect 41797 12937 41831 12971
rect 42901 12937 42935 12971
rect 45017 12937 45051 12971
rect 33241 12869 33275 12903
rect 40325 12869 40359 12903
rect 22201 12801 22235 12835
rect 22477 12801 22511 12835
rect 22661 12801 22695 12835
rect 32505 12801 32539 12835
rect 33885 12801 33919 12835
rect 34152 12801 34186 12835
rect 36369 12801 36403 12835
rect 37473 12801 37507 12835
rect 37657 12801 37691 12835
rect 40233 12801 40267 12835
rect 40417 12801 40451 12835
rect 40555 12801 40589 12835
rect 41153 12801 41187 12835
rect 41246 12801 41280 12835
rect 41429 12801 41463 12835
rect 41521 12801 41555 12835
rect 41618 12801 41652 12835
rect 42901 12801 42935 12835
rect 43177 12801 43211 12835
rect 44281 12801 44315 12835
rect 44925 12801 44959 12835
rect 45109 12801 45143 12835
rect 47041 12801 47075 12835
rect 36461 12733 36495 12767
rect 36737 12733 36771 12767
rect 40693 12733 40727 12767
rect 44097 12733 44131 12767
rect 37565 12665 37599 12699
rect 42993 12665 43027 12699
rect 35265 12597 35299 12631
rect 44465 12597 44499 12631
rect 47133 12597 47167 12631
rect 47961 12597 47995 12631
rect 34345 12393 34379 12427
rect 37105 12393 37139 12427
rect 40969 12393 41003 12427
rect 42809 12393 42843 12427
rect 43177 12393 43211 12427
rect 43913 12393 43947 12427
rect 36461 12325 36495 12359
rect 44097 12325 44131 12359
rect 20729 12257 20763 12291
rect 36553 12257 36587 12291
rect 46489 12257 46523 12291
rect 46673 12257 46707 12291
rect 48237 12257 48271 12291
rect 2237 12189 2271 12223
rect 20996 12189 21030 12223
rect 22753 12189 22787 12223
rect 23029 12189 23063 12223
rect 23213 12189 23247 12223
rect 25237 12189 25271 12223
rect 25513 12189 25547 12223
rect 25697 12189 25731 12223
rect 26525 12189 26559 12223
rect 33793 12189 33827 12223
rect 34161 12189 34195 12223
rect 36277 12189 36311 12223
rect 37013 12189 37047 12223
rect 37197 12189 37231 12223
rect 41153 12189 41187 12223
rect 41429 12189 41463 12223
rect 42993 12189 43027 12223
rect 43269 12189 43303 12223
rect 26792 12121 26826 12155
rect 33977 12121 34011 12155
rect 34069 12121 34103 12155
rect 43729 12121 43763 12155
rect 22109 12053 22143 12087
rect 22569 12053 22603 12087
rect 25053 12053 25087 12087
rect 27905 12053 27939 12087
rect 36093 12053 36127 12087
rect 41337 12053 41371 12087
rect 43939 12053 43973 12087
rect 29929 11849 29963 11883
rect 30849 11849 30883 11883
rect 33977 11849 34011 11883
rect 43085 11849 43119 11883
rect 37657 11781 37691 11815
rect 2053 11713 2087 11747
rect 22477 11713 22511 11747
rect 22753 11713 22787 11747
rect 22937 11713 22971 11747
rect 24501 11713 24535 11747
rect 24777 11713 24811 11747
rect 24961 11713 24995 11747
rect 25605 11713 25639 11747
rect 27169 11713 27203 11747
rect 27353 11713 27387 11747
rect 27445 11713 27479 11747
rect 27721 11713 27755 11747
rect 27905 11713 27939 11747
rect 28641 11713 28675 11747
rect 28825 11713 28859 11747
rect 29009 11713 29043 11747
rect 29101 11713 29135 11747
rect 29561 11713 29595 11747
rect 29745 11713 29779 11747
rect 30021 11713 30055 11747
rect 30665 11713 30699 11747
rect 30941 11713 30975 11747
rect 32781 11713 32815 11747
rect 33793 11713 33827 11747
rect 33977 11713 34011 11747
rect 36461 11713 36495 11747
rect 37473 11713 37507 11747
rect 38393 11713 38427 11747
rect 42717 11713 42751 11747
rect 43637 11713 43671 11747
rect 43729 11713 43763 11747
rect 44557 11713 44591 11747
rect 44833 11713 44867 11747
rect 2237 11645 2271 11679
rect 2789 11645 2823 11679
rect 25881 11645 25915 11679
rect 27537 11645 27571 11679
rect 32505 11645 32539 11679
rect 32597 11645 32631 11679
rect 32689 11645 32723 11679
rect 36921 11645 36955 11679
rect 38669 11645 38703 11679
rect 42809 11645 42843 11679
rect 43913 11645 43947 11679
rect 44649 11577 44683 11611
rect 44741 11577 44775 11611
rect 22293 11509 22327 11543
rect 24317 11509 24351 11543
rect 25421 11509 25455 11543
rect 25789 11509 25823 11543
rect 30481 11509 30515 11543
rect 32321 11509 32355 11543
rect 36553 11509 36587 11543
rect 37841 11509 37875 11543
rect 38485 11509 38519 11543
rect 38577 11509 38611 11543
rect 42901 11509 42935 11543
rect 43821 11509 43855 11543
rect 44373 11509 44407 11543
rect 2329 11305 2363 11339
rect 29837 11305 29871 11339
rect 32413 11305 32447 11339
rect 36921 11305 36955 11339
rect 43085 11305 43119 11339
rect 44649 11305 44683 11339
rect 26065 11237 26099 11271
rect 37841 11237 37875 11271
rect 21925 11169 21959 11203
rect 35449 11169 35483 11203
rect 43453 11169 43487 11203
rect 44281 11169 44315 11203
rect 2237 11101 2271 11135
rect 3065 11101 3099 11135
rect 3985 11101 4019 11135
rect 12541 11101 12575 11135
rect 13001 11101 13035 11135
rect 24685 11101 24719 11135
rect 27537 11101 27571 11135
rect 27721 11101 27755 11135
rect 28365 11101 28399 11135
rect 28549 11101 28583 11135
rect 29009 11101 29043 11135
rect 29193 11101 29227 11135
rect 29745 11101 29779 11135
rect 30021 11101 30055 11135
rect 31033 11101 31067 11135
rect 33149 11101 33183 11135
rect 33333 11101 33367 11135
rect 33793 11101 33827 11135
rect 33977 11101 34011 11135
rect 35357 11101 35391 11135
rect 36645 11101 36679 11135
rect 36737 11101 36771 11135
rect 37841 11101 37875 11135
rect 38025 11101 38059 11135
rect 38485 11101 38519 11135
rect 38761 11101 38795 11135
rect 39129 11101 39163 11135
rect 43269 11101 43303 11135
rect 43545 11101 43579 11135
rect 44465 11101 44499 11135
rect 45201 11101 45235 11135
rect 45569 11101 45603 11135
rect 22192 11033 22226 11067
rect 24952 11033 24986 11067
rect 28181 11033 28215 11067
rect 29101 11033 29135 11067
rect 29929 11033 29963 11067
rect 31300 11033 31334 11067
rect 45385 11033 45419 11067
rect 45477 11033 45511 11067
rect 4077 10965 4111 10999
rect 13093 10965 13127 10999
rect 23305 10965 23339 10999
rect 27721 10965 27755 10999
rect 33241 10965 33275 10999
rect 33977 10965 34011 10999
rect 35725 10965 35759 10999
rect 45753 10965 45787 10999
rect 22477 10761 22511 10795
rect 25329 10761 25363 10795
rect 30021 10761 30055 10795
rect 33425 10761 33459 10795
rect 38117 10761 38151 10795
rect 38669 10761 38703 10795
rect 40509 10761 40543 10795
rect 47041 10761 47075 10795
rect 2881 10693 2915 10727
rect 12541 10693 12575 10727
rect 31401 10693 31435 10727
rect 35541 10693 35575 10727
rect 36645 10693 36679 10727
rect 45906 10693 45940 10727
rect 22661 10625 22695 10659
rect 23949 10625 23983 10659
rect 24216 10625 24250 10659
rect 27169 10625 27203 10659
rect 27353 10625 27387 10659
rect 27537 10625 27571 10659
rect 27721 10625 27755 10659
rect 28917 10625 28951 10659
rect 29101 10625 29135 10659
rect 29653 10625 29687 10659
rect 30757 10625 30791 10659
rect 30941 10625 30975 10659
rect 31585 10625 31619 10659
rect 32689 10625 32723 10659
rect 32873 10625 32907 10659
rect 33057 10625 33091 10659
rect 33241 10625 33275 10659
rect 35357 10625 35391 10659
rect 35633 10625 35667 10659
rect 35725 10625 35759 10659
rect 36829 10625 36863 10659
rect 36921 10625 36955 10659
rect 37933 10625 37967 10659
rect 38209 10625 38243 10659
rect 38945 10625 38979 10659
rect 39037 10625 39071 10659
rect 39405 10625 39439 10659
rect 40325 10625 40359 10659
rect 40601 10625 40635 10659
rect 41061 10625 41095 10659
rect 41245 10625 41279 10659
rect 41349 10625 41383 10659
rect 44189 10625 44223 10659
rect 44373 10625 44407 10659
rect 44925 10625 44959 10659
rect 45109 10625 45143 10659
rect 45661 10625 45695 10659
rect 2697 10557 2731 10591
rect 3157 10557 3191 10591
rect 12357 10557 12391 10591
rect 14197 10557 14231 10591
rect 22937 10557 22971 10591
rect 27445 10557 27479 10591
rect 29745 10557 29779 10591
rect 32965 10557 32999 10591
rect 39129 10557 39163 10591
rect 44097 10557 44131 10591
rect 44281 10557 44315 10591
rect 30849 10489 30883 10523
rect 37749 10489 37783 10523
rect 22845 10421 22879 10455
rect 27905 10421 27939 10455
rect 29009 10421 29043 10455
rect 29837 10421 29871 10455
rect 31769 10421 31803 10455
rect 35909 10421 35943 10455
rect 36921 10421 36955 10455
rect 39221 10421 39255 10455
rect 40141 10421 40175 10455
rect 41153 10421 41187 10455
rect 43913 10421 43947 10455
rect 45017 10421 45051 10455
rect 24593 10217 24627 10251
rect 27537 10217 27571 10251
rect 29009 10217 29043 10251
rect 29745 10217 29779 10251
rect 30941 10217 30975 10251
rect 33333 10217 33367 10251
rect 36277 10217 36311 10251
rect 42165 10217 42199 10251
rect 45569 10217 45603 10251
rect 24961 10149 24995 10183
rect 29193 10149 29227 10183
rect 30849 10149 30883 10183
rect 31861 10149 31895 10183
rect 34069 10149 34103 10183
rect 41613 10149 41647 10183
rect 44373 10149 44407 10183
rect 21833 10081 21867 10115
rect 25053 10081 25087 10115
rect 26157 10081 26191 10115
rect 28089 10081 28123 10115
rect 31033 10081 31067 10115
rect 31493 10081 31527 10115
rect 33057 10081 33091 10115
rect 34897 10081 34931 10115
rect 43453 10081 43487 10115
rect 43913 10081 43947 10115
rect 2329 10013 2363 10047
rect 24777 10013 24811 10047
rect 26424 10013 26458 10047
rect 27997 10013 28031 10047
rect 28181 10013 28215 10047
rect 29929 10013 29963 10047
rect 30205 10013 30239 10047
rect 30757 10013 30791 10047
rect 31677 10013 31711 10047
rect 31769 10013 31803 10047
rect 31953 10013 31987 10047
rect 32965 10013 32999 10047
rect 33793 10013 33827 10047
rect 35164 10013 35198 10047
rect 38209 10013 38243 10047
rect 38301 10013 38335 10047
rect 38393 10013 38427 10047
rect 38531 10013 38565 10047
rect 38669 10013 38703 10047
rect 39313 10013 39347 10047
rect 40233 10013 40267 10047
rect 42073 10013 42107 10047
rect 43545 10013 43579 10047
rect 43821 10013 43855 10047
rect 44373 10013 44407 10047
rect 44649 10013 44683 10047
rect 45201 10013 45235 10047
rect 22100 9945 22134 9979
rect 28825 9945 28859 9979
rect 29041 9945 29075 9979
rect 30113 9945 30147 9979
rect 39129 9945 39163 9979
rect 40478 9945 40512 9979
rect 45385 9945 45419 9979
rect 23213 9877 23247 9911
rect 34253 9877 34287 9911
rect 38025 9877 38059 9911
rect 39497 9877 39531 9911
rect 43269 9877 43303 9911
rect 44557 9877 44591 9911
rect 22385 9673 22419 9707
rect 30021 9673 30055 9707
rect 32873 9673 32907 9707
rect 44005 9673 44039 9707
rect 40509 9605 40543 9639
rect 42892 9605 42926 9639
rect 44833 9605 44867 9639
rect 2053 9537 2087 9571
rect 22569 9537 22603 9571
rect 22753 9537 22787 9571
rect 22845 9537 22879 9571
rect 27905 9537 27939 9571
rect 28089 9537 28123 9571
rect 28733 9537 28767 9571
rect 29561 9537 29595 9571
rect 31401 9537 31435 9571
rect 32413 9537 32447 9571
rect 35633 9537 35667 9571
rect 37473 9537 37507 9571
rect 37740 9537 37774 9571
rect 39313 9537 39347 9571
rect 39497 9537 39531 9571
rect 40417 9537 40451 9571
rect 40601 9537 40635 9571
rect 40719 9537 40753 9571
rect 40877 9537 40911 9571
rect 41521 9537 41555 9571
rect 42625 9537 42659 9571
rect 44465 9537 44499 9571
rect 2237 9469 2271 9503
rect 2789 9469 2823 9503
rect 27997 9469 28031 9503
rect 28825 9469 28859 9503
rect 31493 9469 31527 9503
rect 35725 9469 35759 9503
rect 36001 9469 36035 9503
rect 40233 9469 40267 9503
rect 41429 9469 41463 9503
rect 41889 9469 41923 9503
rect 31769 9401 31803 9435
rect 39405 9401 39439 9435
rect 45017 9401 45051 9435
rect 29009 9333 29043 9367
rect 29745 9333 29779 9367
rect 31401 9333 31435 9367
rect 32505 9333 32539 9367
rect 38853 9333 38887 9367
rect 44833 9333 44867 9367
rect 2329 9129 2363 9163
rect 32045 9129 32079 9163
rect 39313 9129 39347 9163
rect 48053 9129 48087 9163
rect 44097 9061 44131 9095
rect 43821 8993 43855 9027
rect 2237 8925 2271 8959
rect 31953 8925 31987 8959
rect 32137 8925 32171 8959
rect 39221 8925 39255 8959
rect 39405 8925 39439 8959
rect 43729 8925 43763 8959
rect 47961 8857 47995 8891
rect 47869 8449 47903 8483
rect 48053 8381 48087 8415
rect 2329 7837 2363 7871
rect 2789 7837 2823 7871
rect 2881 7701 2915 7735
rect 2237 7429 2271 7463
rect 2053 7361 2087 7395
rect 2789 7293 2823 7327
rect 47961 7157 47995 7191
rect 2789 6817 2823 6851
rect 46489 6817 46523 6851
rect 48237 6817 48271 6851
rect 1593 6749 1627 6783
rect 1777 6681 1811 6715
rect 46673 6681 46707 6715
rect 2881 6409 2915 6443
rect 47869 6409 47903 6443
rect 2329 6273 2363 6307
rect 2789 6273 2823 6307
rect 39037 6273 39071 6307
rect 46397 6273 46431 6307
rect 47777 6273 47811 6307
rect 39129 6069 39163 6103
rect 45937 6069 45971 6103
rect 46489 6069 46523 6103
rect 47225 6069 47259 6103
rect 46489 5729 46523 5763
rect 48237 5729 48271 5763
rect 1869 5661 1903 5695
rect 2329 5661 2363 5695
rect 3157 5661 3191 5695
rect 9781 5661 9815 5695
rect 10241 5661 10275 5695
rect 39221 5661 39255 5695
rect 46029 5661 46063 5695
rect 46673 5593 46707 5627
rect 2421 5525 2455 5559
rect 10333 5525 10367 5559
rect 39221 5253 39255 5287
rect 45569 5253 45603 5287
rect 47869 5253 47903 5287
rect 39037 5185 39071 5219
rect 44741 5185 44775 5219
rect 47777 5185 47811 5219
rect 1777 5117 1811 5151
rect 2237 5117 2271 5151
rect 2421 5117 2455 5151
rect 2973 5117 3007 5151
rect 40049 5117 40083 5151
rect 45385 5117 45419 5151
rect 47225 5117 47259 5151
rect 44281 4981 44315 5015
rect 44833 4981 44867 5015
rect 47593 4777 47627 4811
rect 1593 4641 1627 4675
rect 1777 4641 1811 4675
rect 2789 4641 2823 4675
rect 9873 4641 9907 4675
rect 10057 4641 10091 4675
rect 10333 4641 10367 4675
rect 45201 4641 45235 4675
rect 45385 4641 45419 4675
rect 45661 4641 45695 4675
rect 4169 4573 4203 4607
rect 4997 4573 5031 4607
rect 5549 4573 5583 4607
rect 43821 4573 43855 4607
rect 44649 4573 44683 4607
rect 47501 4573 47535 4607
rect 48145 4573 48179 4607
rect 6285 4505 6319 4539
rect 43913 4437 43947 4471
rect 48237 4437 48271 4471
rect 43269 4165 43303 4199
rect 2145 4097 2179 4131
rect 2789 4097 2823 4131
rect 2881 4097 2915 4131
rect 6653 4097 6687 4131
rect 10517 4097 10551 4131
rect 19349 4097 19383 4131
rect 39957 4097 39991 4131
rect 41429 4097 41463 4131
rect 43085 4097 43119 4131
rect 47777 4097 47811 4131
rect 3801 4029 3835 4063
rect 3985 4029 4019 4063
rect 4261 4029 4295 4063
rect 20821 4029 20855 4063
rect 22017 4029 22051 4063
rect 22201 4029 22235 4063
rect 22569 4029 22603 4063
rect 44925 4029 44959 4063
rect 45385 4029 45419 4063
rect 45569 4029 45603 4063
rect 47225 4029 47259 4063
rect 2237 3893 2271 3927
rect 6745 3893 6779 3927
rect 7481 3893 7515 3927
rect 10609 3893 10643 3927
rect 13185 3893 13219 3927
rect 17049 3893 17083 3927
rect 18613 3893 18647 3927
rect 19441 3893 19475 3927
rect 20177 3893 20211 3927
rect 25421 3893 25455 3927
rect 26249 3893 26283 3927
rect 27445 3893 27479 3927
rect 40049 3893 40083 3927
rect 40969 3893 41003 3927
rect 41521 3893 41555 3927
rect 47869 3893 47903 3927
rect 2789 3689 2823 3723
rect 3341 3689 3375 3723
rect 22201 3689 22235 3723
rect 6469 3553 6503 3587
rect 10701 3553 10735 3587
rect 10977 3553 11011 3587
rect 16773 3553 16807 3587
rect 17417 3553 17451 3587
rect 19717 3553 19751 3587
rect 19901 3553 19935 3587
rect 20637 3553 20671 3587
rect 25973 3553 26007 3587
rect 26433 3553 26467 3587
rect 40785 3553 40819 3587
rect 40969 3553 41003 3587
rect 41521 3553 41555 3587
rect 44005 3553 44039 3587
rect 45937 3553 45971 3587
rect 46121 3553 46155 3587
rect 47041 3553 47075 3587
rect 1961 3485 1995 3519
rect 3249 3485 3283 3519
rect 4077 3485 4111 3519
rect 4721 3485 4755 3519
rect 5549 3485 5583 3519
rect 6009 3485 6043 3519
rect 8309 3485 8343 3519
rect 10517 3485 10551 3519
rect 13001 3485 13035 3519
rect 16129 3485 16163 3519
rect 22109 3485 22143 3519
rect 24685 3485 24719 3519
rect 25329 3485 25363 3519
rect 28273 3485 28307 3519
rect 32045 3485 32079 3519
rect 32505 3485 32539 3519
rect 40233 3485 40267 3519
rect 43269 3485 43303 3519
rect 44649 3485 44683 3519
rect 45201 3485 45235 3519
rect 2053 3417 2087 3451
rect 4813 3417 4847 3451
rect 6193 3417 6227 3451
rect 16221 3417 16255 3451
rect 16957 3417 16991 3451
rect 25421 3417 25455 3451
rect 26157 3417 26191 3451
rect 4169 3349 4203 3383
rect 8401 3349 8435 3383
rect 13093 3349 13127 3383
rect 24777 3349 24811 3383
rect 28365 3349 28399 3383
rect 32597 3349 32631 3383
rect 45293 3349 45327 3383
rect 2053 3077 2087 3111
rect 4353 3077 4387 3111
rect 7481 3077 7515 3111
rect 13185 3077 13219 3111
rect 24961 3077 24995 3111
rect 27353 3077 27387 3111
rect 32505 3077 32539 3111
rect 40141 3077 40175 3111
rect 45109 3077 45143 3111
rect 1869 3009 1903 3043
rect 7297 3009 7331 3043
rect 10701 3009 10735 3043
rect 13001 3009 13035 3043
rect 17325 3009 17359 3043
rect 19625 3009 19659 3043
rect 24777 3009 24811 3043
rect 27169 3009 27203 3043
rect 32321 3009 32355 3043
rect 39957 3009 39991 3043
rect 42625 3009 42659 3043
rect 44925 3009 44959 3043
rect 48053 3009 48087 3043
rect 2789 2941 2823 2975
rect 4169 2941 4203 2975
rect 5181 2941 5215 2975
rect 7757 2941 7791 2975
rect 13553 2941 13587 2975
rect 17509 2941 17543 2975
rect 19165 2941 19199 2975
rect 19809 2941 19843 2975
rect 21465 2941 21499 2975
rect 25789 2941 25823 2975
rect 27721 2941 27755 2975
rect 32781 2941 32815 2975
rect 40601 2941 40635 2975
rect 42809 2941 42843 2975
rect 43085 2941 43119 2975
rect 45753 2941 45787 2975
rect 6837 2805 6871 2839
rect 48237 2805 48271 2839
rect 1961 2601 1995 2635
rect 14473 2601 14507 2635
rect 18521 2601 18555 2635
rect 19533 2601 19567 2635
rect 41705 2601 41739 2635
rect 47961 2601 47995 2635
rect 11897 2533 11931 2567
rect 44189 2533 44223 2567
rect 3985 2465 4019 2499
rect 4169 2465 4203 2499
rect 4537 2465 4571 2499
rect 6653 2465 6687 2499
rect 7113 2465 7147 2499
rect 20361 2465 20395 2499
rect 45385 2465 45419 2499
rect 45569 2465 45603 2499
rect 46857 2465 46891 2499
rect 11713 2397 11747 2431
rect 14289 2397 14323 2431
rect 18429 2397 18463 2431
rect 19441 2397 19475 2431
rect 20085 2397 20119 2431
rect 38761 2397 38795 2431
rect 41613 2397 41647 2431
rect 1685 2329 1719 2363
rect 2605 2329 2639 2363
rect 6837 2329 6871 2363
rect 29837 2329 29871 2363
rect 44005 2329 44039 2363
rect 2881 2261 2915 2295
rect 29929 2261 29963 2295
rect 38945 2261 38979 2295
<< metal1 >>
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 17681 47175 17739 47181
rect 17681 47141 17693 47175
rect 17727 47172 17739 47175
rect 17954 47172 17960 47184
rect 17727 47144 17960 47172
rect 17727 47141 17739 47144
rect 17681 47135 17739 47141
rect 17954 47132 17960 47144
rect 18012 47132 18018 47184
rect 32214 47132 32220 47184
rect 32272 47172 32278 47184
rect 32493 47175 32551 47181
rect 32493 47172 32505 47175
rect 32272 47144 32505 47172
rect 32272 47132 32278 47144
rect 32493 47141 32505 47144
rect 32539 47141 32551 47175
rect 32493 47135 32551 47141
rect 42797 47175 42855 47181
rect 42797 47141 42809 47175
rect 42843 47172 42855 47175
rect 42886 47172 42892 47184
rect 42843 47144 42892 47172
rect 42843 47141 42855 47144
rect 42797 47135 42855 47141
rect 42886 47132 42892 47144
rect 42944 47132 42950 47184
rect 3421 47107 3479 47113
rect 3421 47073 3433 47107
rect 3467 47104 3479 47107
rect 4154 47104 4160 47116
rect 3467 47076 4160 47104
rect 3467 47073 3479 47076
rect 3421 47067 3479 47073
rect 4154 47064 4160 47076
rect 4212 47064 4218 47116
rect 7190 47104 7196 47116
rect 4816 47076 7196 47104
rect 2130 47036 2136 47048
rect 2091 47008 2136 47036
rect 2130 46996 2136 47008
rect 2188 46996 2194 47048
rect 2685 47039 2743 47045
rect 2685 47005 2697 47039
rect 2731 47036 2743 47039
rect 3973 47039 4031 47045
rect 3973 47036 3985 47039
rect 2731 47008 3985 47036
rect 2731 47005 2743 47008
rect 2685 46999 2743 47005
rect 3973 47005 3985 47008
rect 4019 47036 4031 47039
rect 4062 47036 4068 47048
rect 4019 47008 4068 47036
rect 4019 47005 4031 47008
rect 3973 46999 4031 47005
rect 4062 46996 4068 47008
rect 4120 46996 4126 47048
rect 4816 46980 4844 47076
rect 7190 47064 7196 47076
rect 7248 47064 7254 47116
rect 9030 47064 9036 47116
rect 9088 47104 9094 47116
rect 9125 47107 9183 47113
rect 9125 47104 9137 47107
rect 9088 47076 9137 47104
rect 9088 47064 9094 47076
rect 9125 47073 9137 47076
rect 9171 47073 9183 47107
rect 9125 47067 9183 47073
rect 14182 47064 14188 47116
rect 14240 47104 14246 47116
rect 14737 47107 14795 47113
rect 14737 47104 14749 47107
rect 14240 47076 14749 47104
rect 14240 47064 14246 47076
rect 14737 47073 14749 47076
rect 14783 47073 14795 47107
rect 47210 47104 47216 47116
rect 47171 47076 47216 47104
rect 14737 47067 14795 47073
rect 47210 47064 47216 47076
rect 47268 47064 47274 47116
rect 5350 46996 5356 47048
rect 5408 47036 5414 47048
rect 5445 47039 5503 47045
rect 5445 47036 5457 47039
rect 5408 47008 5457 47036
rect 5408 46996 5414 47008
rect 5445 47005 5457 47008
rect 5491 47005 5503 47039
rect 6546 47036 6552 47048
rect 6507 47008 6552 47036
rect 5445 46999 5503 47005
rect 6546 46996 6552 47008
rect 6604 46996 6610 47048
rect 7374 47036 7380 47048
rect 7335 47008 7380 47036
rect 7374 46996 7380 47008
rect 7432 46996 7438 47048
rect 8846 46996 8852 47048
rect 8904 47036 8910 47048
rect 9401 47039 9459 47045
rect 9401 47036 9413 47039
rect 8904 47008 9413 47036
rect 8904 46996 8910 47008
rect 9401 47005 9413 47008
rect 9447 47005 9459 47039
rect 12710 47036 12716 47048
rect 12671 47008 12716 47036
rect 9401 46999 9459 47005
rect 12710 46996 12716 47008
rect 12768 46996 12774 47048
rect 13725 47039 13783 47045
rect 13725 47005 13737 47039
rect 13771 47036 13783 47039
rect 14277 47039 14335 47045
rect 14277 47036 14289 47039
rect 13771 47008 14289 47036
rect 13771 47005 13783 47008
rect 13725 46999 13783 47005
rect 14277 47005 14289 47008
rect 14323 47005 14335 47039
rect 14277 46999 14335 47005
rect 17402 46996 17408 47048
rect 17460 47036 17466 47048
rect 17497 47039 17555 47045
rect 17497 47036 17509 47039
rect 17460 47008 17509 47036
rect 17460 46996 17466 47008
rect 17497 47005 17509 47008
rect 17543 47005 17555 47039
rect 17497 46999 17555 47005
rect 19334 46996 19340 47048
rect 19392 47036 19398 47048
rect 19521 47039 19579 47045
rect 19521 47036 19533 47039
rect 19392 47008 19533 47036
rect 19392 46996 19398 47008
rect 19521 47005 19533 47008
rect 19567 47005 19579 47039
rect 19521 46999 19579 47005
rect 22462 46996 22468 47048
rect 22520 47036 22526 47048
rect 22925 47039 22983 47045
rect 22925 47036 22937 47039
rect 22520 47008 22937 47036
rect 22520 46996 22526 47008
rect 22925 47005 22937 47008
rect 22971 47005 22983 47039
rect 22925 46999 22983 47005
rect 23842 46996 23848 47048
rect 23900 47036 23906 47048
rect 24673 47039 24731 47045
rect 24673 47036 24685 47039
rect 23900 47008 24685 47036
rect 23900 46996 23906 47008
rect 24673 47005 24685 47008
rect 24719 47005 24731 47039
rect 25682 47036 25688 47048
rect 25643 47008 25688 47036
rect 24673 46999 24731 47005
rect 25682 46996 25688 47008
rect 25740 46996 25746 47048
rect 29730 46996 29736 47048
rect 29788 47036 29794 47048
rect 30009 47039 30067 47045
rect 30009 47036 30021 47039
rect 29788 47008 30021 47036
rect 29788 46996 29794 47008
rect 30009 47005 30021 47008
rect 30055 47005 30067 47039
rect 30009 46999 30067 47005
rect 31754 46996 31760 47048
rect 31812 47036 31818 47048
rect 32309 47039 32367 47045
rect 32309 47036 32321 47039
rect 31812 47008 32321 47036
rect 31812 46996 31818 47008
rect 32309 47005 32321 47008
rect 32355 47005 32367 47039
rect 33226 47036 33232 47048
rect 33187 47008 33232 47036
rect 32309 46999 32367 47005
rect 33226 46996 33232 47008
rect 33284 46996 33290 47048
rect 38565 47039 38623 47045
rect 38565 47005 38577 47039
rect 38611 47036 38623 47039
rect 39758 47036 39764 47048
rect 38611 47008 39764 47036
rect 38611 47005 38623 47008
rect 38565 46999 38623 47005
rect 39758 46996 39764 47008
rect 39816 46996 39822 47048
rect 40218 47036 40224 47048
rect 40179 47008 40224 47036
rect 40218 46996 40224 47008
rect 40276 46996 40282 47048
rect 41414 47036 41420 47048
rect 41375 47008 41420 47036
rect 41414 46996 41420 47008
rect 41472 46996 41478 47048
rect 42518 46996 42524 47048
rect 42576 47036 42582 47048
rect 42613 47039 42671 47045
rect 42613 47036 42625 47039
rect 42576 47008 42625 47036
rect 42576 46996 42582 47008
rect 42613 47005 42625 47008
rect 42659 47005 42671 47039
rect 45370 47036 45376 47048
rect 45331 47008 45376 47036
rect 42613 46999 42671 47005
rect 45370 46996 45376 47008
rect 45428 46996 45434 47048
rect 47949 47039 48007 47045
rect 47949 47005 47961 47039
rect 47995 47036 48007 47039
rect 48958 47036 48964 47048
rect 47995 47008 48964 47036
rect 47995 47005 48007 47008
rect 47949 46999 48007 47005
rect 48958 46996 48964 47008
rect 49016 46996 49022 47048
rect 4798 46968 4804 46980
rect 4759 46940 4804 46968
rect 4798 46928 4804 46940
rect 4856 46928 4862 46980
rect 5626 46928 5632 46980
rect 5684 46968 5690 46980
rect 6641 46971 6699 46977
rect 6641 46968 6653 46971
rect 5684 46940 6653 46968
rect 5684 46928 5690 46940
rect 6641 46937 6653 46940
rect 6687 46937 6699 46971
rect 6641 46931 6699 46937
rect 13814 46928 13820 46980
rect 13872 46968 13878 46980
rect 14461 46971 14519 46977
rect 14461 46968 14473 46971
rect 13872 46940 14473 46968
rect 13872 46928 13878 46940
rect 14461 46937 14473 46940
rect 14507 46937 14519 46971
rect 19702 46968 19708 46980
rect 19663 46940 19708 46968
rect 14461 46931 14519 46937
rect 19702 46928 19708 46940
rect 19760 46928 19766 46980
rect 25041 46971 25099 46977
rect 25041 46937 25053 46971
rect 25087 46968 25099 46971
rect 25406 46968 25412 46980
rect 25087 46940 25412 46968
rect 25087 46937 25099 46940
rect 25041 46931 25099 46937
rect 25406 46928 25412 46940
rect 25464 46928 25470 46980
rect 45554 46928 45560 46980
rect 45612 46968 45618 46980
rect 45612 46940 45657 46968
rect 45612 46928 45618 46940
rect 5534 46900 5540 46912
rect 5495 46872 5540 46900
rect 5534 46860 5540 46872
rect 5592 46860 5598 46912
rect 46382 46860 46388 46912
rect 46440 46900 46446 46912
rect 46934 46900 46940 46912
rect 46440 46872 46940 46900
rect 46440 46860 46446 46872
rect 46934 46860 46940 46872
rect 46992 46860 46998 46912
rect 48038 46900 48044 46912
rect 47999 46872 48044 46900
rect 48038 46860 48044 46872
rect 48096 46860 48102 46912
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 2590 46588 2596 46640
rect 2648 46628 2654 46640
rect 5997 46631 6055 46637
rect 5997 46628 6009 46631
rect 2648 46600 6009 46628
rect 2648 46588 2654 46600
rect 5997 46597 6009 46600
rect 6043 46597 6055 46631
rect 12710 46628 12716 46640
rect 5997 46591 6055 46597
rect 11992 46600 12716 46628
rect 4154 46560 4160 46572
rect 4115 46532 4160 46560
rect 4154 46520 4160 46532
rect 4212 46520 4218 46572
rect 11992 46569 12020 46600
rect 12710 46588 12716 46600
rect 12768 46588 12774 46640
rect 25682 46628 25688 46640
rect 24780 46600 25688 46628
rect 11977 46563 12035 46569
rect 11977 46529 11989 46563
rect 12023 46529 12035 46563
rect 22462 46560 22468 46572
rect 22423 46532 22468 46560
rect 11977 46523 12035 46529
rect 22462 46520 22468 46532
rect 22520 46520 22526 46572
rect 24780 46569 24808 46600
rect 25682 46588 25688 46600
rect 25740 46588 25746 46640
rect 33226 46628 33232 46640
rect 32876 46600 33232 46628
rect 32876 46569 32904 46600
rect 33226 46588 33232 46600
rect 33284 46588 33290 46640
rect 47213 46631 47271 46637
rect 47213 46597 47225 46631
rect 47259 46628 47271 46631
rect 48314 46628 48320 46640
rect 47259 46600 48320 46628
rect 47259 46597 47271 46600
rect 47213 46591 47271 46597
rect 48314 46588 48320 46600
rect 48372 46588 48378 46640
rect 24765 46563 24823 46569
rect 24765 46529 24777 46563
rect 24811 46529 24823 46563
rect 24765 46523 24823 46529
rect 32861 46563 32919 46569
rect 32861 46529 32873 46563
rect 32907 46529 32919 46563
rect 39758 46560 39764 46572
rect 39719 46532 39764 46560
rect 32861 46523 32919 46529
rect 39758 46520 39764 46532
rect 39816 46520 39822 46572
rect 41414 46520 41420 46572
rect 41472 46560 41478 46572
rect 42613 46563 42671 46569
rect 42613 46560 42625 46563
rect 41472 46532 42625 46560
rect 41472 46520 41478 46532
rect 42613 46529 42625 46532
rect 42659 46529 42671 46563
rect 47762 46560 47768 46572
rect 47723 46532 47768 46560
rect 42613 46523 42671 46529
rect 47762 46520 47768 46532
rect 47820 46520 47826 46572
rect 1857 46495 1915 46501
rect 1857 46461 1869 46495
rect 1903 46461 1915 46495
rect 2038 46492 2044 46504
rect 1999 46464 2044 46492
rect 1857 46455 1915 46461
rect 1872 46424 1900 46455
rect 2038 46452 2044 46464
rect 2096 46452 2102 46504
rect 2314 46492 2320 46504
rect 2275 46464 2320 46492
rect 2314 46452 2320 46464
rect 2372 46452 2378 46504
rect 4341 46495 4399 46501
rect 4341 46461 4353 46495
rect 4387 46492 4399 46495
rect 5902 46492 5908 46504
rect 4387 46464 5908 46492
rect 4387 46461 4399 46464
rect 4341 46455 4399 46461
rect 5902 46452 5908 46464
rect 5960 46452 5966 46504
rect 12161 46495 12219 46501
rect 12161 46461 12173 46495
rect 12207 46492 12219 46495
rect 12526 46492 12532 46504
rect 12207 46464 12532 46492
rect 12207 46461 12219 46464
rect 12161 46455 12219 46461
rect 12526 46452 12532 46464
rect 12584 46452 12590 46504
rect 12894 46492 12900 46504
rect 12855 46464 12900 46492
rect 12894 46452 12900 46464
rect 12952 46452 12958 46504
rect 14274 46492 14280 46504
rect 14235 46464 14280 46492
rect 14274 46452 14280 46464
rect 14332 46452 14338 46504
rect 14458 46492 14464 46504
rect 14419 46464 14464 46492
rect 14458 46452 14464 46464
rect 14516 46452 14522 46504
rect 14826 46492 14832 46504
rect 14787 46464 14832 46492
rect 14826 46452 14832 46464
rect 14884 46452 14890 46504
rect 22649 46495 22707 46501
rect 22649 46461 22661 46495
rect 22695 46492 22707 46495
rect 22738 46492 22744 46504
rect 22695 46464 22744 46492
rect 22695 46461 22707 46464
rect 22649 46455 22707 46461
rect 22738 46452 22744 46464
rect 22796 46452 22802 46504
rect 23198 46492 23204 46504
rect 23159 46464 23204 46492
rect 23198 46452 23204 46464
rect 23256 46452 23262 46504
rect 24946 46492 24952 46504
rect 24907 46464 24952 46492
rect 24946 46452 24952 46464
rect 25004 46452 25010 46504
rect 25774 46492 25780 46504
rect 25735 46464 25780 46492
rect 25774 46452 25780 46464
rect 25832 46452 25838 46504
rect 28537 46495 28595 46501
rect 28537 46461 28549 46495
rect 28583 46492 28595 46495
rect 28997 46495 29055 46501
rect 28997 46492 29009 46495
rect 28583 46464 29009 46492
rect 28583 46461 28595 46464
rect 28537 46455 28595 46461
rect 28997 46461 29009 46464
rect 29043 46461 29055 46495
rect 29178 46492 29184 46504
rect 29139 46464 29184 46492
rect 28997 46455 29055 46461
rect 29178 46452 29184 46464
rect 29236 46452 29242 46504
rect 29638 46492 29644 46504
rect 29599 46464 29644 46492
rect 29638 46452 29644 46464
rect 29696 46452 29702 46504
rect 33045 46495 33103 46501
rect 33045 46461 33057 46495
rect 33091 46492 33103 46495
rect 33134 46492 33140 46504
rect 33091 46464 33140 46492
rect 33091 46461 33103 46464
rect 33045 46455 33103 46461
rect 33134 46452 33140 46464
rect 33192 46452 33198 46504
rect 33502 46492 33508 46504
rect 33463 46464 33508 46492
rect 33502 46452 33508 46464
rect 33560 46452 33566 46504
rect 36449 46495 36507 46501
rect 36449 46461 36461 46495
rect 36495 46492 36507 46495
rect 37461 46495 37519 46501
rect 37461 46492 37473 46495
rect 36495 46464 37473 46492
rect 36495 46461 36507 46464
rect 36449 46455 36507 46461
rect 37461 46461 37473 46464
rect 37507 46461 37519 46495
rect 37642 46492 37648 46504
rect 37603 46464 37648 46492
rect 37461 46455 37519 46461
rect 37642 46452 37648 46464
rect 37700 46452 37706 46504
rect 37921 46495 37979 46501
rect 37921 46461 37933 46495
rect 37967 46461 37979 46495
rect 39942 46492 39948 46504
rect 39903 46464 39948 46492
rect 37921 46455 37979 46461
rect 7377 46427 7435 46433
rect 7377 46424 7389 46427
rect 1872 46396 7389 46424
rect 7377 46393 7389 46396
rect 7423 46393 7435 46427
rect 7377 46387 7435 46393
rect 36722 46384 36728 46436
rect 36780 46424 36786 46436
rect 37936 46424 37964 46455
rect 39942 46452 39948 46464
rect 40000 46452 40006 46504
rect 40221 46495 40279 46501
rect 40221 46461 40233 46495
rect 40267 46461 40279 46495
rect 42794 46492 42800 46504
rect 42755 46464 42800 46492
rect 40221 46455 40279 46461
rect 36780 46396 37964 46424
rect 36780 46384 36786 46396
rect 38654 46384 38660 46436
rect 38712 46424 38718 46436
rect 40236 46424 40264 46455
rect 42794 46452 42800 46464
rect 42852 46452 42858 46504
rect 43073 46495 43131 46501
rect 43073 46461 43085 46495
rect 43119 46461 43131 46495
rect 45370 46492 45376 46504
rect 45331 46464 45376 46492
rect 43073 46455 43131 46461
rect 38712 46396 40264 46424
rect 38712 46384 38718 46396
rect 41874 46384 41880 46436
rect 41932 46424 41938 46436
rect 43088 46424 43116 46455
rect 45370 46452 45376 46464
rect 45428 46452 45434 46504
rect 45557 46495 45615 46501
rect 45557 46461 45569 46495
rect 45603 46492 45615 46495
rect 47026 46492 47032 46504
rect 45603 46464 47032 46492
rect 45603 46461 45615 46464
rect 45557 46455 45615 46461
rect 47026 46452 47032 46464
rect 47084 46452 47090 46504
rect 41932 46396 43116 46424
rect 41932 46384 41938 46396
rect 5258 46316 5264 46368
rect 5316 46356 5322 46368
rect 6733 46359 6791 46365
rect 6733 46356 6745 46359
rect 5316 46328 6745 46356
rect 5316 46316 5322 46328
rect 6733 46325 6745 46328
rect 6779 46325 6791 46359
rect 8018 46356 8024 46368
rect 7979 46328 8024 46356
rect 6733 46319 6791 46325
rect 8018 46316 8024 46328
rect 8076 46316 8082 46368
rect 15010 46316 15016 46368
rect 15068 46356 15074 46368
rect 17037 46359 17095 46365
rect 17037 46356 17049 46359
rect 15068 46328 17049 46356
rect 15068 46316 15074 46328
rect 17037 46325 17049 46328
rect 17083 46325 17095 46359
rect 17037 46319 17095 46325
rect 35434 46316 35440 46368
rect 35492 46356 35498 46368
rect 35713 46359 35771 46365
rect 35713 46356 35725 46359
rect 35492 46328 35725 46356
rect 35492 46316 35498 46328
rect 35713 46325 35725 46328
rect 35759 46325 35771 46359
rect 35713 46319 35771 46325
rect 46658 46316 46664 46368
rect 46716 46356 46722 46368
rect 47857 46359 47915 46365
rect 47857 46356 47869 46359
rect 46716 46328 47869 46356
rect 46716 46316 46722 46328
rect 47857 46325 47869 46328
rect 47903 46325 47915 46359
rect 47857 46319 47915 46325
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 2038 46112 2044 46164
rect 2096 46152 2102 46164
rect 7653 46155 7711 46161
rect 7653 46152 7665 46155
rect 2096 46124 7665 46152
rect 2096 46112 2102 46124
rect 7653 46121 7665 46124
rect 7699 46121 7711 46155
rect 12526 46152 12532 46164
rect 12487 46124 12532 46152
rect 7653 46115 7711 46121
rect 12526 46112 12532 46124
rect 12584 46112 12590 46164
rect 13633 46155 13691 46161
rect 13633 46121 13645 46155
rect 13679 46152 13691 46155
rect 13814 46152 13820 46164
rect 13679 46124 13820 46152
rect 13679 46121 13691 46124
rect 13633 46115 13691 46121
rect 13814 46112 13820 46124
rect 13872 46112 13878 46164
rect 14458 46152 14464 46164
rect 14419 46124 14464 46152
rect 14458 46112 14464 46124
rect 14516 46112 14522 46164
rect 22738 46152 22744 46164
rect 22699 46124 22744 46152
rect 22738 46112 22744 46124
rect 22796 46112 22802 46164
rect 29089 46155 29147 46161
rect 29089 46121 29101 46155
rect 29135 46152 29147 46155
rect 29178 46152 29184 46164
rect 29135 46124 29184 46152
rect 29135 46121 29147 46124
rect 29089 46115 29147 46121
rect 29178 46112 29184 46124
rect 29236 46112 29242 46164
rect 33134 46152 33140 46164
rect 33095 46124 33140 46152
rect 33134 46112 33140 46124
rect 33192 46112 33198 46164
rect 38473 46155 38531 46161
rect 38473 46121 38485 46155
rect 38519 46152 38531 46155
rect 39942 46152 39948 46164
rect 38519 46124 39948 46152
rect 38519 46121 38531 46124
rect 38473 46115 38531 46121
rect 39942 46112 39948 46124
rect 40000 46112 40006 46164
rect 45370 46152 45376 46164
rect 45331 46124 45376 46152
rect 45370 46112 45376 46124
rect 45428 46112 45434 46164
rect 45554 46112 45560 46164
rect 45612 46152 45618 46164
rect 45925 46155 45983 46161
rect 45925 46152 45937 46155
rect 45612 46124 45937 46152
rect 45612 46112 45618 46124
rect 45925 46121 45937 46124
rect 45971 46121 45983 46155
rect 45925 46115 45983 46121
rect 8018 46084 8024 46096
rect 1596 46056 8024 46084
rect 1596 46025 1624 46056
rect 8018 46044 8024 46056
rect 8076 46044 8082 46096
rect 41322 46084 41328 46096
rect 12452 46056 41328 46084
rect 1581 46019 1639 46025
rect 1581 45985 1593 46019
rect 1627 45985 1639 46019
rect 2774 46016 2780 46028
rect 2735 45988 2780 46016
rect 1581 45979 1639 45985
rect 2774 45976 2780 45988
rect 2832 45976 2838 46028
rect 5258 46016 5264 46028
rect 5219 45988 5264 46016
rect 5258 45976 5264 45988
rect 5316 45976 5322 46028
rect 5445 46019 5503 46025
rect 5445 45985 5457 46019
rect 5491 46016 5503 46019
rect 5534 46016 5540 46028
rect 5491 45988 5540 46016
rect 5491 45985 5503 45988
rect 5445 45979 5503 45985
rect 5534 45976 5540 45988
rect 5592 45976 5598 46028
rect 5810 46016 5816 46028
rect 5771 45988 5816 46016
rect 5810 45976 5816 45988
rect 5868 45976 5874 46028
rect 12452 45960 12480 46056
rect 41322 46044 41328 46056
rect 41380 46044 41386 46096
rect 15010 46016 15016 46028
rect 14971 45988 15016 46016
rect 15010 45976 15016 45988
rect 15068 45976 15074 46028
rect 15470 46016 15476 46028
rect 15431 45988 15476 46016
rect 15470 45976 15476 45988
rect 15528 45976 15534 46028
rect 19058 45976 19064 46028
rect 19116 46016 19122 46028
rect 35434 46016 35440 46028
rect 19116 45988 35296 46016
rect 35395 45988 35440 46016
rect 19116 45976 19122 45988
rect 4062 45948 4068 45960
rect 4023 45920 4068 45948
rect 4062 45908 4068 45920
rect 4120 45908 4126 45960
rect 6914 45908 6920 45960
rect 6972 45948 6978 45960
rect 7561 45951 7619 45957
rect 7561 45948 7573 45951
rect 6972 45920 7573 45948
rect 6972 45908 6978 45920
rect 7561 45917 7573 45920
rect 7607 45917 7619 45951
rect 7561 45911 7619 45917
rect 1765 45883 1823 45889
rect 1765 45849 1777 45883
rect 1811 45849 1823 45883
rect 4614 45880 4620 45892
rect 4575 45852 4620 45880
rect 1765 45843 1823 45849
rect 1780 45812 1808 45843
rect 4614 45840 4620 45852
rect 4672 45840 4678 45892
rect 4890 45840 4896 45892
rect 4948 45880 4954 45892
rect 5534 45880 5540 45892
rect 4948 45852 5540 45880
rect 4948 45840 4954 45852
rect 5534 45840 5540 45852
rect 5592 45840 5598 45892
rect 7576 45880 7604 45911
rect 12434 45908 12440 45960
rect 12492 45948 12498 45960
rect 13541 45951 13599 45957
rect 12492 45920 12585 45948
rect 12492 45908 12498 45920
rect 13541 45917 13553 45951
rect 13587 45948 13599 45951
rect 14369 45951 14427 45957
rect 14369 45948 14381 45951
rect 13587 45920 14381 45948
rect 13587 45917 13599 45920
rect 13541 45911 13599 45917
rect 14369 45917 14381 45920
rect 14415 45917 14427 45951
rect 22646 45948 22652 45960
rect 22607 45920 22652 45948
rect 14369 45911 14427 45917
rect 13556 45880 13584 45911
rect 7576 45852 13584 45880
rect 7282 45812 7288 45824
rect 1780 45784 7288 45812
rect 7282 45772 7288 45784
rect 7340 45772 7346 45824
rect 14384 45812 14412 45911
rect 22646 45908 22652 45920
rect 22704 45908 22710 45960
rect 24029 45951 24087 45957
rect 24029 45917 24041 45951
rect 24075 45948 24087 45951
rect 24673 45951 24731 45957
rect 24673 45948 24685 45951
rect 24075 45920 24685 45948
rect 24075 45917 24087 45920
rect 24029 45911 24087 45917
rect 24673 45917 24685 45920
rect 24719 45917 24731 45951
rect 24673 45911 24731 45917
rect 28997 45951 29055 45957
rect 28997 45917 29009 45951
rect 29043 45948 29055 45951
rect 29178 45948 29184 45960
rect 29043 45920 29184 45948
rect 29043 45917 29055 45920
rect 28997 45911 29055 45917
rect 29178 45908 29184 45920
rect 29236 45908 29242 45960
rect 29730 45948 29736 45960
rect 29691 45920 29736 45948
rect 29730 45908 29736 45920
rect 29788 45908 29794 45960
rect 32950 45908 32956 45960
rect 33008 45948 33014 45960
rect 33045 45951 33103 45957
rect 33045 45948 33057 45951
rect 33008 45920 33057 45948
rect 33008 45908 33014 45920
rect 33045 45917 33057 45920
rect 33091 45917 33103 45951
rect 33045 45911 33103 45917
rect 15194 45880 15200 45892
rect 15155 45852 15200 45880
rect 15194 45840 15200 45852
rect 15252 45840 15258 45892
rect 24854 45880 24860 45892
rect 24815 45852 24860 45880
rect 24854 45840 24860 45852
rect 24912 45840 24918 45892
rect 25130 45840 25136 45892
rect 25188 45880 25194 45892
rect 26513 45883 26571 45889
rect 26513 45880 26525 45883
rect 25188 45852 26525 45880
rect 25188 45840 25194 45852
rect 26513 45849 26525 45852
rect 26559 45849 26571 45883
rect 29914 45880 29920 45892
rect 29875 45852 29920 45880
rect 26513 45843 26571 45849
rect 29914 45840 29920 45852
rect 29972 45840 29978 45892
rect 30282 45840 30288 45892
rect 30340 45880 30346 45892
rect 31573 45883 31631 45889
rect 31573 45880 31585 45883
rect 30340 45852 31585 45880
rect 30340 45840 30346 45852
rect 31573 45849 31585 45852
rect 31619 45849 31631 45883
rect 31573 45843 31631 45849
rect 34514 45812 34520 45824
rect 14384 45784 34520 45812
rect 34514 45772 34520 45784
rect 34572 45772 34578 45824
rect 35268 45812 35296 45988
rect 35434 45976 35440 45988
rect 35492 45976 35498 46028
rect 36078 46016 36084 46028
rect 36039 45988 36084 46016
rect 36078 45976 36084 45988
rect 36136 45976 36142 46028
rect 40037 46019 40095 46025
rect 40037 45985 40049 46019
rect 40083 46016 40095 46019
rect 40218 46016 40224 46028
rect 40083 45988 40224 46016
rect 40083 45985 40095 45988
rect 40037 45979 40095 45985
rect 40218 45976 40224 45988
rect 40276 45976 40282 46028
rect 40586 46016 40592 46028
rect 40547 45988 40592 46016
rect 40586 45976 40592 45988
rect 40644 45976 40650 46028
rect 46658 46016 46664 46028
rect 46619 45988 46664 46016
rect 46658 45976 46664 45988
rect 46716 45976 46722 46028
rect 48222 46016 48228 46028
rect 48183 45988 48228 46016
rect 48222 45976 48228 45988
rect 48280 45976 48286 46028
rect 38381 45951 38439 45957
rect 38381 45917 38393 45951
rect 38427 45948 38439 45951
rect 38654 45948 38660 45960
rect 38427 45920 38660 45948
rect 38427 45917 38439 45920
rect 38381 45911 38439 45917
rect 38654 45908 38660 45920
rect 38712 45948 38718 45960
rect 39942 45948 39948 45960
rect 38712 45920 39948 45948
rect 38712 45908 38718 45920
rect 39942 45908 39948 45920
rect 40000 45908 40006 45960
rect 45830 45948 45836 45960
rect 45791 45920 45836 45948
rect 45830 45908 45836 45920
rect 45888 45908 45894 45960
rect 46474 45948 46480 45960
rect 46435 45920 46480 45948
rect 46474 45908 46480 45920
rect 46532 45908 46538 45960
rect 35618 45880 35624 45892
rect 35579 45852 35624 45880
rect 35618 45840 35624 45852
rect 35676 45840 35682 45892
rect 40218 45880 40224 45892
rect 40179 45852 40224 45880
rect 40218 45840 40224 45852
rect 40276 45840 40282 45892
rect 46566 45812 46572 45824
rect 35268 45784 46572 45812
rect 46566 45772 46572 45784
rect 46624 45772 46630 45824
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 4614 45568 4620 45620
rect 4672 45608 4678 45620
rect 10042 45608 10048 45620
rect 4672 45580 10048 45608
rect 4672 45568 4678 45580
rect 10042 45568 10048 45580
rect 10100 45568 10106 45620
rect 15194 45568 15200 45620
rect 15252 45608 15258 45620
rect 15289 45611 15347 45617
rect 15289 45608 15301 45611
rect 15252 45580 15301 45608
rect 15252 45568 15258 45580
rect 15289 45577 15301 45580
rect 15335 45577 15347 45611
rect 22646 45608 22652 45620
rect 15289 45571 15347 45577
rect 22066 45580 22652 45608
rect 2317 45543 2375 45549
rect 2317 45509 2329 45543
rect 2363 45540 2375 45543
rect 5626 45540 5632 45552
rect 2363 45512 5632 45540
rect 2363 45509 2375 45512
rect 2317 45503 2375 45509
rect 5626 45500 5632 45512
rect 5684 45500 5690 45552
rect 5902 45500 5908 45552
rect 5960 45540 5966 45552
rect 6641 45543 6699 45549
rect 6641 45540 6653 45543
rect 5960 45512 6653 45540
rect 5960 45500 5966 45512
rect 6641 45509 6653 45512
rect 6687 45509 6699 45543
rect 7282 45540 7288 45552
rect 7243 45512 7288 45540
rect 6641 45503 6699 45509
rect 7282 45500 7288 45512
rect 7340 45500 7346 45552
rect 22066 45540 22094 45580
rect 22646 45568 22652 45580
rect 22704 45608 22710 45620
rect 24854 45608 24860 45620
rect 22704 45580 24716 45608
rect 24815 45580 24860 45608
rect 22704 45568 22710 45580
rect 10336 45512 22094 45540
rect 24688 45540 24716 45580
rect 24854 45568 24860 45580
rect 24912 45568 24918 45620
rect 24946 45568 24952 45620
rect 25004 45608 25010 45620
rect 25501 45611 25559 45617
rect 25501 45608 25513 45611
rect 25004 45580 25513 45608
rect 25004 45568 25010 45580
rect 25501 45577 25513 45580
rect 25547 45577 25559 45611
rect 29825 45611 29883 45617
rect 25501 45571 25559 45577
rect 25608 45580 29776 45608
rect 25608 45540 25636 45580
rect 24688 45512 25636 45540
rect 29748 45540 29776 45580
rect 29825 45577 29837 45611
rect 29871 45608 29883 45611
rect 29914 45608 29920 45620
rect 29871 45580 29920 45608
rect 29871 45577 29883 45580
rect 29825 45571 29883 45577
rect 29914 45568 29920 45580
rect 29972 45568 29978 45620
rect 32950 45608 32956 45620
rect 30024 45580 32956 45608
rect 30024 45540 30052 45580
rect 32950 45568 32956 45580
rect 33008 45568 33014 45620
rect 35529 45611 35587 45617
rect 35529 45577 35541 45611
rect 35575 45608 35587 45611
rect 35618 45608 35624 45620
rect 35575 45580 35624 45608
rect 35575 45577 35587 45580
rect 35529 45571 35587 45577
rect 35618 45568 35624 45580
rect 35676 45568 35682 45620
rect 40037 45611 40095 45617
rect 40037 45577 40049 45611
rect 40083 45608 40095 45611
rect 40218 45608 40224 45620
rect 40083 45580 40224 45608
rect 40083 45577 40095 45580
rect 40037 45571 40095 45577
rect 40218 45568 40224 45580
rect 40276 45568 40282 45620
rect 29748 45512 30052 45540
rect 36357 45543 36415 45549
rect 4801 45475 4859 45481
rect 4801 45441 4813 45475
rect 4847 45472 4859 45475
rect 4890 45472 4896 45484
rect 4847 45444 4896 45472
rect 4847 45441 4859 45444
rect 4801 45435 4859 45441
rect 4890 45432 4896 45444
rect 4948 45432 4954 45484
rect 6549 45475 6607 45481
rect 6549 45472 6561 45475
rect 5460 45444 6561 45472
rect 5460 45416 5488 45444
rect 6549 45441 6561 45444
rect 6595 45472 6607 45475
rect 7190 45472 7196 45484
rect 6595 45444 6914 45472
rect 7103 45444 7196 45472
rect 6595 45441 6607 45444
rect 6549 45435 6607 45441
rect 2133 45407 2191 45413
rect 2133 45373 2145 45407
rect 2179 45373 2191 45407
rect 2958 45404 2964 45416
rect 2919 45376 2964 45404
rect 2133 45367 2191 45373
rect 2148 45336 2176 45367
rect 2958 45364 2964 45376
rect 3016 45364 3022 45416
rect 5442 45404 5448 45416
rect 5403 45376 5448 45404
rect 5442 45364 5448 45376
rect 5500 45364 5506 45416
rect 6886 45404 6914 45444
rect 7190 45432 7196 45444
rect 7248 45472 7254 45484
rect 10336 45472 10364 45512
rect 36357 45509 36369 45543
rect 36403 45540 36415 45543
rect 37642 45540 37648 45552
rect 36403 45512 37648 45540
rect 36403 45509 36415 45512
rect 36357 45503 36415 45509
rect 37642 45500 37648 45512
rect 37700 45500 37706 45552
rect 41417 45543 41475 45549
rect 41417 45509 41429 45543
rect 41463 45540 41475 45543
rect 42794 45540 42800 45552
rect 41463 45512 42800 45540
rect 41463 45509 41475 45512
rect 41417 45503 41475 45509
rect 42794 45500 42800 45512
rect 42852 45500 42858 45552
rect 45922 45500 45928 45552
rect 45980 45540 45986 45552
rect 47026 45540 47032 45552
rect 45980 45512 46612 45540
rect 46987 45512 47032 45540
rect 45980 45500 45986 45512
rect 7248 45444 10364 45472
rect 7248 45432 7254 45444
rect 14274 45432 14280 45484
rect 14332 45472 14338 45484
rect 14461 45475 14519 45481
rect 14461 45472 14473 45475
rect 14332 45444 14473 45472
rect 14332 45432 14338 45444
rect 14461 45441 14473 45444
rect 14507 45441 14519 45475
rect 15194 45472 15200 45484
rect 15155 45444 15200 45472
rect 14461 45435 14519 45441
rect 15194 45432 15200 45444
rect 15252 45432 15258 45484
rect 24765 45475 24823 45481
rect 24765 45472 24777 45475
rect 22066 45444 24777 45472
rect 22066 45404 22094 45444
rect 24765 45441 24777 45444
rect 24811 45472 24823 45475
rect 25409 45475 25467 45481
rect 25409 45472 25421 45475
rect 24811 45444 25421 45472
rect 24811 45441 24823 45444
rect 24765 45435 24823 45441
rect 25409 45441 25421 45444
rect 25455 45472 25467 45475
rect 29178 45472 29184 45484
rect 25455 45444 29184 45472
rect 25455 45441 25467 45444
rect 25409 45435 25467 45441
rect 29178 45432 29184 45444
rect 29236 45432 29242 45484
rect 29730 45472 29736 45484
rect 29691 45444 29736 45472
rect 29730 45432 29736 45444
rect 29788 45432 29794 45484
rect 34514 45432 34520 45484
rect 34572 45472 34578 45484
rect 35437 45475 35495 45481
rect 35437 45472 35449 45475
rect 34572 45444 35449 45472
rect 34572 45432 34578 45444
rect 35437 45441 35449 45444
rect 35483 45472 35495 45475
rect 35618 45472 35624 45484
rect 35483 45444 35624 45472
rect 35483 45441 35495 45444
rect 35437 45435 35495 45441
rect 35618 45432 35624 45444
rect 35676 45432 35682 45484
rect 36265 45475 36323 45481
rect 36265 45441 36277 45475
rect 36311 45472 36323 45475
rect 38654 45472 38660 45484
rect 36311 45444 38660 45472
rect 36311 45441 36323 45444
rect 36265 45435 36323 45441
rect 38654 45432 38660 45444
rect 38712 45432 38718 45484
rect 39942 45472 39948 45484
rect 39855 45444 39948 45472
rect 39942 45432 39948 45444
rect 40000 45472 40006 45484
rect 40586 45472 40592 45484
rect 40000 45444 40592 45472
rect 40000 45432 40006 45444
rect 40586 45432 40592 45444
rect 40644 45432 40650 45484
rect 41322 45472 41328 45484
rect 41283 45444 41328 45472
rect 41322 45432 41328 45444
rect 41380 45432 41386 45484
rect 45462 45432 45468 45484
rect 45520 45472 45526 45484
rect 45833 45475 45891 45481
rect 45833 45472 45845 45475
rect 45520 45444 45845 45472
rect 45520 45432 45526 45444
rect 45833 45441 45845 45444
rect 45879 45441 45891 45475
rect 46474 45472 46480 45484
rect 46435 45444 46480 45472
rect 45833 45435 45891 45441
rect 46474 45432 46480 45444
rect 46532 45432 46538 45484
rect 46584 45472 46612 45512
rect 47026 45500 47032 45512
rect 47084 45500 47090 45552
rect 46937 45475 46995 45481
rect 46937 45472 46949 45475
rect 46584 45444 46949 45472
rect 46937 45441 46949 45444
rect 46983 45472 46995 45475
rect 47762 45472 47768 45484
rect 46983 45444 47768 45472
rect 46983 45441 46995 45444
rect 46937 45435 46995 45441
rect 47762 45432 47768 45444
rect 47820 45432 47826 45484
rect 6886 45376 22094 45404
rect 7374 45336 7380 45348
rect 2148 45308 7380 45336
rect 7374 45296 7380 45308
rect 7432 45296 7438 45348
rect 15194 45296 15200 45348
rect 15252 45336 15258 45348
rect 47762 45336 47768 45348
rect 15252 45308 41414 45336
rect 15252 45296 15258 45308
rect 10502 45228 10508 45280
rect 10560 45268 10566 45280
rect 10689 45271 10747 45277
rect 10689 45268 10701 45271
rect 10560 45240 10701 45268
rect 10560 45228 10566 45240
rect 10689 45237 10701 45240
rect 10735 45237 10747 45271
rect 41386 45268 41414 45308
rect 45526 45308 47768 45336
rect 45526 45268 45554 45308
rect 47762 45296 47768 45308
rect 47820 45296 47826 45348
rect 41386 45240 45554 45268
rect 10689 45231 10747 45237
rect 46474 45228 46480 45280
rect 46532 45268 46538 45280
rect 47949 45271 48007 45277
rect 47949 45268 47961 45271
rect 46532 45240 47961 45268
rect 46532 45228 46538 45240
rect 47949 45237 47961 45240
rect 47995 45237 48007 45271
rect 47949 45231 48007 45237
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 6822 44928 6828 44940
rect 6783 44900 6828 44928
rect 6822 44888 6828 44900
rect 6880 44888 6886 44940
rect 10502 44928 10508 44940
rect 10463 44900 10508 44928
rect 10502 44888 10508 44900
rect 10560 44888 10566 44940
rect 11054 44928 11060 44940
rect 11015 44900 11060 44928
rect 11054 44888 11060 44900
rect 11112 44888 11118 44940
rect 40586 44928 40592 44940
rect 40547 44900 40592 44928
rect 40586 44888 40592 44900
rect 40644 44888 40650 44940
rect 46474 44928 46480 44940
rect 46435 44900 46480 44928
rect 46474 44888 46480 44900
rect 46532 44888 46538 44940
rect 48222 44928 48228 44940
rect 48183 44900 48228 44928
rect 48222 44888 48228 44900
rect 48280 44888 48286 44940
rect 14 44820 20 44872
rect 72 44860 78 44872
rect 1581 44863 1639 44869
rect 1581 44860 1593 44863
rect 72 44832 1593 44860
rect 72 44820 78 44832
rect 1581 44829 1593 44832
rect 1627 44829 1639 44863
rect 1581 44823 1639 44829
rect 2593 44863 2651 44869
rect 2593 44829 2605 44863
rect 2639 44860 2651 44863
rect 3973 44863 4031 44869
rect 3973 44860 3985 44863
rect 2639 44832 3985 44860
rect 2639 44829 2651 44832
rect 2593 44823 2651 44829
rect 3973 44829 3985 44832
rect 4019 44860 4031 44863
rect 4062 44860 4068 44872
rect 4019 44832 4068 44860
rect 4019 44829 4031 44832
rect 3973 44823 4031 44829
rect 4062 44820 4068 44832
rect 4120 44860 4126 44872
rect 4890 44860 4896 44872
rect 4120 44832 4896 44860
rect 4120 44820 4126 44832
rect 4890 44820 4896 44832
rect 4948 44860 4954 44872
rect 6181 44863 6239 44869
rect 6181 44860 6193 44863
rect 4948 44832 6193 44860
rect 4948 44820 4954 44832
rect 6181 44829 6193 44832
rect 6227 44829 6239 44863
rect 40034 44860 40040 44872
rect 39995 44832 40040 44860
rect 6181 44823 6239 44829
rect 40034 44820 40040 44832
rect 40092 44860 40098 44872
rect 45830 44860 45836 44872
rect 40092 44832 45836 44860
rect 40092 44820 40098 44832
rect 45830 44820 45836 44832
rect 45888 44820 45894 44872
rect 3237 44795 3295 44801
rect 3237 44761 3249 44795
rect 3283 44792 3295 44795
rect 3786 44792 3792 44804
rect 3283 44764 3792 44792
rect 3283 44761 3295 44764
rect 3237 44755 3295 44761
rect 3786 44752 3792 44764
rect 3844 44792 3850 44804
rect 5350 44792 5356 44804
rect 3844 44764 5356 44792
rect 3844 44752 3850 44764
rect 5350 44752 5356 44764
rect 5408 44752 5414 44804
rect 10686 44792 10692 44804
rect 10647 44764 10692 44792
rect 10686 44752 10692 44764
rect 10744 44752 10750 44804
rect 46661 44795 46719 44801
rect 46661 44761 46673 44795
rect 46707 44792 46719 44795
rect 47854 44792 47860 44804
rect 46707 44764 47860 44792
rect 46707 44761 46719 44764
rect 46661 44755 46719 44761
rect 47854 44752 47860 44764
rect 47912 44752 47918 44804
rect 1762 44724 1768 44736
rect 1723 44696 1768 44724
rect 1762 44684 1768 44696
rect 1820 44684 1826 44736
rect 5258 44724 5264 44736
rect 5219 44696 5264 44724
rect 5258 44684 5264 44696
rect 5316 44724 5322 44736
rect 12434 44724 12440 44736
rect 5316 44696 12440 44724
rect 5316 44684 5322 44696
rect 12434 44684 12440 44696
rect 12492 44684 12498 44736
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 10597 44523 10655 44529
rect 10597 44489 10609 44523
rect 10643 44520 10655 44523
rect 10686 44520 10692 44532
rect 10643 44492 10692 44520
rect 10643 44489 10655 44492
rect 10597 44483 10655 44489
rect 10686 44480 10692 44492
rect 10744 44480 10750 44532
rect 47854 44520 47860 44532
rect 47815 44492 47860 44520
rect 47854 44480 47860 44492
rect 47912 44480 47918 44532
rect 6886 44424 20392 44452
rect 4890 44384 4896 44396
rect 4851 44356 4896 44384
rect 4890 44344 4896 44356
rect 4948 44344 4954 44396
rect 5350 44344 5356 44396
rect 5408 44384 5414 44396
rect 6886 44384 6914 44424
rect 5408 44356 6914 44384
rect 5408 44344 5414 44356
rect 10042 44344 10048 44396
rect 10100 44384 10106 44396
rect 20364 44393 20392 44424
rect 10505 44387 10563 44393
rect 10505 44384 10517 44387
rect 10100 44356 10517 44384
rect 10100 44344 10106 44356
rect 10505 44353 10517 44356
rect 10551 44353 10563 44387
rect 10505 44347 10563 44353
rect 20349 44387 20407 44393
rect 20349 44353 20361 44387
rect 20395 44384 20407 44387
rect 29730 44384 29736 44396
rect 20395 44356 29736 44384
rect 20395 44353 20407 44356
rect 20349 44347 20407 44353
rect 29730 44344 29736 44356
rect 29788 44344 29794 44396
rect 47762 44384 47768 44396
rect 47723 44356 47768 44384
rect 47762 44344 47768 44356
rect 47820 44344 47826 44396
rect 2041 44319 2099 44325
rect 2041 44285 2053 44319
rect 2087 44285 2099 44319
rect 2041 44279 2099 44285
rect 2225 44319 2283 44325
rect 2225 44285 2237 44319
rect 2271 44316 2283 44319
rect 2314 44316 2320 44328
rect 2271 44288 2320 44316
rect 2271 44285 2283 44288
rect 2225 44279 2283 44285
rect 2056 44248 2084 44279
rect 2314 44276 2320 44288
rect 2372 44276 2378 44328
rect 2774 44316 2780 44328
rect 2735 44288 2780 44316
rect 2774 44276 2780 44288
rect 2832 44276 2838 44328
rect 4798 44276 4804 44328
rect 4856 44316 4862 44328
rect 5077 44319 5135 44325
rect 5077 44316 5089 44319
rect 4856 44288 5089 44316
rect 4856 44276 4862 44288
rect 5077 44285 5089 44288
rect 5123 44316 5135 44319
rect 40034 44316 40040 44328
rect 5123 44288 40040 44316
rect 5123 44285 5135 44288
rect 5077 44279 5135 44285
rect 40034 44276 40040 44288
rect 40092 44276 40098 44328
rect 3050 44248 3056 44260
rect 2056 44220 3056 44248
rect 3050 44208 3056 44220
rect 3108 44208 3114 44260
rect 20441 44183 20499 44189
rect 20441 44149 20453 44183
rect 20487 44180 20499 44183
rect 20530 44180 20536 44192
rect 20487 44152 20536 44180
rect 20487 44149 20499 44152
rect 20441 44143 20499 44149
rect 20530 44140 20536 44152
rect 20588 44140 20594 44192
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 3878 43936 3884 43988
rect 3936 43976 3942 43988
rect 6546 43976 6552 43988
rect 3936 43948 6552 43976
rect 3936 43936 3942 43948
rect 6546 43936 6552 43948
rect 6604 43976 6610 43988
rect 15194 43976 15200 43988
rect 6604 43948 15200 43976
rect 6604 43936 6610 43948
rect 15194 43936 15200 43948
rect 15252 43936 15258 43988
rect 29730 43908 29736 43920
rect 29691 43880 29736 43908
rect 29730 43868 29736 43880
rect 29788 43868 29794 43920
rect 2774 43840 2780 43852
rect 2735 43812 2780 43840
rect 2774 43800 2780 43812
rect 2832 43800 2838 43852
rect 4982 43840 4988 43852
rect 4943 43812 4988 43840
rect 4982 43800 4988 43812
rect 5040 43800 5046 43852
rect 20530 43840 20536 43852
rect 20491 43812 20536 43840
rect 20530 43800 20536 43812
rect 20588 43800 20594 43852
rect 22189 43843 22247 43849
rect 22189 43809 22201 43843
rect 22235 43840 22247 43843
rect 27062 43840 27068 43852
rect 22235 43812 27068 43840
rect 22235 43809 22247 43812
rect 22189 43803 22247 43809
rect 27062 43800 27068 43812
rect 27120 43800 27126 43852
rect 29822 43800 29828 43852
rect 29880 43840 29886 43852
rect 36538 43840 36544 43852
rect 29880 43812 36544 43840
rect 29880 43800 29886 43812
rect 36538 43800 36544 43812
rect 36596 43800 36602 43852
rect 1578 43772 1584 43784
rect 1539 43744 1584 43772
rect 1578 43732 1584 43744
rect 1636 43732 1642 43784
rect 3694 43732 3700 43784
rect 3752 43772 3758 43784
rect 4617 43775 4675 43781
rect 4617 43772 4629 43775
rect 3752 43744 4629 43772
rect 3752 43732 3758 43744
rect 4617 43741 4629 43744
rect 4663 43772 4675 43775
rect 4890 43772 4896 43784
rect 4663 43744 4896 43772
rect 4663 43741 4675 43744
rect 4617 43735 4675 43741
rect 4890 43732 4896 43744
rect 4948 43732 4954 43784
rect 20346 43772 20352 43784
rect 20307 43744 20352 43772
rect 20346 43732 20352 43744
rect 20404 43732 20410 43784
rect 30009 43775 30067 43781
rect 30009 43741 30021 43775
rect 30055 43772 30067 43775
rect 30098 43772 30104 43784
rect 30055 43744 30104 43772
rect 30055 43741 30067 43744
rect 30009 43735 30067 43741
rect 30098 43732 30104 43744
rect 30156 43732 30162 43784
rect 30466 43772 30472 43784
rect 30427 43744 30472 43772
rect 30466 43732 30472 43744
rect 30524 43732 30530 43784
rect 30650 43772 30656 43784
rect 30611 43744 30656 43772
rect 30650 43732 30656 43744
rect 30708 43732 30714 43784
rect 1765 43707 1823 43713
rect 1765 43673 1777 43707
rect 1811 43704 1823 43707
rect 2406 43704 2412 43716
rect 1811 43676 2412 43704
rect 1811 43673 1823 43676
rect 1765 43667 1823 43673
rect 2406 43664 2412 43676
rect 2464 43664 2470 43716
rect 29733 43707 29791 43713
rect 29733 43673 29745 43707
rect 29779 43704 29791 43707
rect 29822 43704 29828 43716
rect 29779 43676 29828 43704
rect 29779 43673 29791 43676
rect 29733 43667 29791 43673
rect 29822 43664 29828 43676
rect 29880 43664 29886 43716
rect 29917 43639 29975 43645
rect 29917 43605 29929 43639
rect 29963 43636 29975 43639
rect 30653 43639 30711 43645
rect 30653 43636 30665 43639
rect 29963 43608 30665 43636
rect 29963 43605 29975 43608
rect 29917 43599 29975 43605
rect 30653 43605 30665 43608
rect 30699 43636 30711 43639
rect 31110 43636 31116 43648
rect 30699 43608 31116 43636
rect 30699 43605 30711 43608
rect 30653 43599 30711 43605
rect 31110 43596 31116 43608
rect 31168 43596 31174 43648
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 2406 43432 2412 43444
rect 2367 43404 2412 43432
rect 2406 43392 2412 43404
rect 2464 43392 2470 43444
rect 30650 43432 30656 43444
rect 29012 43404 30656 43432
rect 4706 43364 4712 43376
rect 2700 43336 4712 43364
rect 2700 43308 2728 43336
rect 4706 43324 4712 43336
rect 4764 43324 4770 43376
rect 19058 43364 19064 43376
rect 19019 43336 19064 43364
rect 19058 43324 19064 43336
rect 19116 43324 19122 43376
rect 25685 43367 25743 43373
rect 25685 43333 25697 43367
rect 25731 43364 25743 43367
rect 27154 43364 27160 43376
rect 25731 43336 27160 43364
rect 25731 43333 25743 43336
rect 25685 43327 25743 43333
rect 27154 43324 27160 43336
rect 27212 43324 27218 43376
rect 29012 43308 29040 43404
rect 30650 43392 30656 43404
rect 30708 43392 30714 43444
rect 32306 43392 32312 43444
rect 32364 43432 32370 43444
rect 32364 43404 32628 43432
rect 32364 43392 32370 43404
rect 30466 43324 30472 43376
rect 30524 43364 30530 43376
rect 30929 43367 30987 43373
rect 30929 43364 30941 43367
rect 30524 43336 30941 43364
rect 30524 43324 30530 43336
rect 30929 43333 30941 43336
rect 30975 43364 30987 43367
rect 31478 43364 31484 43376
rect 30975 43336 31484 43364
rect 30975 43333 30987 43336
rect 30929 43327 30987 43333
rect 31478 43324 31484 43336
rect 31536 43324 31542 43376
rect 1578 43256 1584 43308
rect 1636 43296 1642 43308
rect 1857 43299 1915 43305
rect 1857 43296 1869 43299
rect 1636 43268 1869 43296
rect 1636 43256 1642 43268
rect 1857 43265 1869 43268
rect 1903 43265 1915 43299
rect 1857 43259 1915 43265
rect 2317 43299 2375 43305
rect 2317 43265 2329 43299
rect 2363 43296 2375 43299
rect 2682 43296 2688 43308
rect 2363 43268 2688 43296
rect 2363 43265 2375 43268
rect 2317 43259 2375 43265
rect 2682 43256 2688 43268
rect 2740 43256 2746 43308
rect 3694 43296 3700 43308
rect 3655 43268 3700 43296
rect 3694 43256 3700 43268
rect 3752 43256 3758 43308
rect 25498 43296 25504 43308
rect 25459 43268 25504 43296
rect 25498 43256 25504 43268
rect 25556 43256 25562 43308
rect 25777 43299 25835 43305
rect 25777 43265 25789 43299
rect 25823 43265 25835 43299
rect 25777 43259 25835 43265
rect 25869 43299 25927 43305
rect 25869 43265 25881 43299
rect 25915 43296 25927 43299
rect 26234 43296 26240 43308
rect 25915 43268 26240 43296
rect 25915 43265 25927 43268
rect 25869 43259 25927 43265
rect 3142 43188 3148 43240
rect 3200 43228 3206 43240
rect 3878 43228 3884 43240
rect 3200 43200 3884 43228
rect 3200 43188 3206 43200
rect 3878 43188 3884 43200
rect 3936 43188 3942 43240
rect 17126 43188 17132 43240
rect 17184 43228 17190 43240
rect 17221 43231 17279 43237
rect 17221 43228 17233 43231
rect 17184 43200 17233 43228
rect 17184 43188 17190 43200
rect 17221 43197 17233 43200
rect 17267 43197 17279 43231
rect 17402 43228 17408 43240
rect 17363 43200 17408 43228
rect 17221 43191 17279 43197
rect 17402 43188 17408 43200
rect 17460 43188 17466 43240
rect 25792 43228 25820 43259
rect 26234 43256 26240 43268
rect 26292 43256 26298 43308
rect 28994 43296 29000 43308
rect 28955 43268 29000 43296
rect 28994 43256 29000 43268
rect 29052 43256 29058 43308
rect 29914 43256 29920 43308
rect 29972 43296 29978 43308
rect 30009 43299 30067 43305
rect 30009 43296 30021 43299
rect 29972 43268 30021 43296
rect 29972 43256 29978 43268
rect 30009 43265 30021 43268
rect 30055 43265 30067 43299
rect 30009 43259 30067 43265
rect 30098 43256 30104 43308
rect 30156 43296 30162 43308
rect 30558 43296 30564 43308
rect 30156 43268 30564 43296
rect 30156 43256 30162 43268
rect 30558 43256 30564 43268
rect 30616 43256 30622 43308
rect 30650 43256 30656 43308
rect 30708 43296 30714 43308
rect 31018 43296 31024 43308
rect 30708 43268 31024 43296
rect 30708 43256 30714 43268
rect 31018 43256 31024 43268
rect 31076 43296 31082 43308
rect 31113 43299 31171 43305
rect 31113 43296 31125 43299
rect 31076 43268 31125 43296
rect 31076 43256 31082 43268
rect 31113 43265 31125 43268
rect 31159 43265 31171 43299
rect 31113 43259 31171 43265
rect 31938 43256 31944 43308
rect 31996 43296 32002 43308
rect 32365 43299 32423 43305
rect 32365 43296 32377 43299
rect 31996 43268 32377 43296
rect 31996 43256 32002 43268
rect 32365 43265 32377 43268
rect 32411 43265 32423 43299
rect 32490 43296 32496 43308
rect 32451 43268 32496 43296
rect 32365 43259 32423 43265
rect 32490 43256 32496 43268
rect 32548 43256 32554 43308
rect 32600 43305 32628 43404
rect 32585 43299 32643 43305
rect 32585 43265 32597 43299
rect 32631 43265 32643 43299
rect 33686 43296 33692 43308
rect 33647 43268 33692 43296
rect 32585 43259 32643 43265
rect 33686 43256 33692 43268
rect 33744 43256 33750 43308
rect 34514 43296 34520 43308
rect 34475 43268 34520 43296
rect 34514 43256 34520 43268
rect 34572 43256 34578 43308
rect 36538 43256 36544 43308
rect 36596 43296 36602 43308
rect 47394 43296 47400 43308
rect 36596 43268 47400 43296
rect 36596 43256 36602 43268
rect 47394 43256 47400 43268
rect 47452 43296 47458 43308
rect 47765 43299 47823 43305
rect 47765 43296 47777 43299
rect 47452 43268 47777 43296
rect 47452 43256 47458 43268
rect 47765 43265 47777 43268
rect 47811 43265 47823 43299
rect 47765 43259 47823 43265
rect 26142 43228 26148 43240
rect 25792 43200 26148 43228
rect 26142 43188 26148 43200
rect 26200 43188 26206 43240
rect 29086 43228 29092 43240
rect 29047 43200 29092 43228
rect 29086 43188 29092 43200
rect 29144 43188 29150 43240
rect 30193 43231 30251 43237
rect 30193 43197 30205 43231
rect 30239 43197 30251 43231
rect 30193 43191 30251 43197
rect 29365 43163 29423 43169
rect 29365 43129 29377 43163
rect 29411 43160 29423 43163
rect 29914 43160 29920 43172
rect 29411 43132 29920 43160
rect 29411 43129 29423 43132
rect 29365 43123 29423 43129
rect 29914 43120 29920 43132
rect 29972 43120 29978 43172
rect 30208 43160 30236 43191
rect 30282 43188 30288 43240
rect 30340 43228 30346 43240
rect 30340 43200 31754 43228
rect 30340 43188 30346 43200
rect 31110 43160 31116 43172
rect 30208 43132 31116 43160
rect 31110 43120 31116 43132
rect 31168 43120 31174 43172
rect 31726 43160 31754 43200
rect 33318 43188 33324 43240
rect 33376 43228 33382 43240
rect 33597 43231 33655 43237
rect 33597 43228 33609 43231
rect 33376 43200 33609 43228
rect 33376 43188 33382 43200
rect 33597 43197 33609 43200
rect 33643 43197 33655 43231
rect 33597 43191 33655 43197
rect 34057 43231 34115 43237
rect 34057 43197 34069 43231
rect 34103 43228 34115 43231
rect 34790 43228 34796 43240
rect 34103 43200 34796 43228
rect 34103 43197 34115 43200
rect 34057 43191 34115 43197
rect 34790 43188 34796 43200
rect 34848 43188 34854 43240
rect 33502 43160 33508 43172
rect 31726 43132 33508 43160
rect 33502 43120 33508 43132
rect 33560 43120 33566 43172
rect 34609 43163 34667 43169
rect 34609 43129 34621 43163
rect 34655 43160 34667 43163
rect 35434 43160 35440 43172
rect 34655 43132 35440 43160
rect 34655 43129 34667 43132
rect 34609 43123 34667 43129
rect 35434 43120 35440 43132
rect 35492 43120 35498 43172
rect 26050 43092 26056 43104
rect 26011 43064 26056 43092
rect 26050 43052 26056 43064
rect 26108 43052 26114 43104
rect 29825 43095 29883 43101
rect 29825 43061 29837 43095
rect 29871 43092 29883 43095
rect 30006 43092 30012 43104
rect 29871 43064 30012 43092
rect 29871 43061 29883 43064
rect 29825 43055 29883 43061
rect 30006 43052 30012 43064
rect 30064 43052 30070 43104
rect 31294 43092 31300 43104
rect 31255 43064 31300 43092
rect 31294 43052 31300 43064
rect 31352 43052 31358 43104
rect 32766 43092 32772 43104
rect 32727 43064 32772 43092
rect 32766 43052 32772 43064
rect 32824 43052 32830 43104
rect 34698 43052 34704 43104
rect 34756 43092 34762 43104
rect 47210 43092 47216 43104
rect 34756 43064 34801 43092
rect 47171 43064 47216 43092
rect 34756 43052 34762 43064
rect 47210 43052 47216 43064
rect 47268 43052 47274 43104
rect 47854 43092 47860 43104
rect 47815 43064 47860 43092
rect 47854 43052 47860 43064
rect 47912 43052 47918 43104
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 17402 42888 17408 42900
rect 17363 42860 17408 42888
rect 17402 42848 17408 42860
rect 17460 42848 17466 42900
rect 27154 42888 27160 42900
rect 27115 42860 27160 42888
rect 27154 42848 27160 42860
rect 27212 42848 27218 42900
rect 29914 42848 29920 42900
rect 29972 42888 29978 42900
rect 29972 42860 32904 42888
rect 29972 42848 29978 42860
rect 22189 42823 22247 42829
rect 22189 42789 22201 42823
rect 22235 42789 22247 42823
rect 22189 42783 22247 42789
rect 2314 42752 2320 42764
rect 2275 42724 2320 42752
rect 2314 42712 2320 42724
rect 2372 42712 2378 42764
rect 3050 42752 3056 42764
rect 3011 42724 3056 42752
rect 3050 42712 3056 42724
rect 3108 42712 3114 42764
rect 5534 42752 5540 42764
rect 5495 42724 5540 42752
rect 5534 42712 5540 42724
rect 5592 42712 5598 42764
rect 22204 42752 22232 42783
rect 29086 42780 29092 42832
rect 29144 42820 29150 42832
rect 29181 42823 29239 42829
rect 29181 42820 29193 42823
rect 29144 42792 29193 42820
rect 29144 42780 29150 42792
rect 29181 42789 29193 42792
rect 29227 42820 29239 42823
rect 32585 42823 32643 42829
rect 32585 42820 32597 42823
rect 29227 42792 30328 42820
rect 29227 42789 29239 42792
rect 29181 42783 29239 42789
rect 30300 42764 30328 42792
rect 30944 42792 32597 42820
rect 22554 42752 22560 42764
rect 22204 42724 22560 42752
rect 22554 42712 22560 42724
rect 22612 42752 22618 42764
rect 23293 42755 23351 42761
rect 23293 42752 23305 42755
rect 22612 42724 23305 42752
rect 22612 42712 22618 42724
rect 23293 42721 23305 42724
rect 23339 42721 23351 42755
rect 27522 42752 27528 42764
rect 23293 42715 23351 42721
rect 26988 42724 27528 42752
rect 1765 42687 1823 42693
rect 1765 42653 1777 42687
rect 1811 42653 1823 42687
rect 1765 42647 1823 42653
rect 2225 42687 2283 42693
rect 2225 42653 2237 42687
rect 2271 42684 2283 42687
rect 2406 42684 2412 42696
rect 2271 42656 2412 42684
rect 2271 42653 2283 42656
rect 2225 42647 2283 42653
rect 1780 42616 1808 42647
rect 2406 42644 2412 42656
rect 2464 42684 2470 42696
rect 4614 42684 4620 42696
rect 2464 42656 4620 42684
rect 2464 42644 2470 42656
rect 4614 42644 4620 42656
rect 4672 42644 4678 42696
rect 4893 42687 4951 42693
rect 4893 42653 4905 42687
rect 4939 42653 4951 42687
rect 4893 42647 4951 42653
rect 2866 42616 2872 42628
rect 1780 42588 2872 42616
rect 2866 42576 2872 42588
rect 2924 42576 2930 42628
rect 1581 42551 1639 42557
rect 1581 42517 1593 42551
rect 1627 42548 1639 42551
rect 2130 42548 2136 42560
rect 1627 42520 2136 42548
rect 1627 42517 1639 42520
rect 1581 42511 1639 42517
rect 2130 42508 2136 42520
rect 2188 42508 2194 42560
rect 4908 42548 4936 42647
rect 13998 42644 14004 42696
rect 14056 42684 14062 42696
rect 17313 42687 17371 42693
rect 17313 42684 17325 42687
rect 14056 42656 17325 42684
rect 14056 42644 14062 42656
rect 17313 42653 17325 42656
rect 17359 42653 17371 42687
rect 17313 42647 17371 42653
rect 19518 42644 19524 42696
rect 19576 42684 19582 42696
rect 19705 42687 19763 42693
rect 19705 42684 19717 42687
rect 19576 42656 19717 42684
rect 19576 42644 19582 42656
rect 19705 42653 19717 42656
rect 19751 42653 19763 42687
rect 19705 42647 19763 42653
rect 20622 42644 20628 42696
rect 20680 42684 20686 42696
rect 20809 42687 20867 42693
rect 20809 42684 20821 42687
rect 20680 42656 20821 42684
rect 20680 42644 20686 42656
rect 20809 42653 20821 42656
rect 20855 42653 20867 42687
rect 22830 42684 22836 42696
rect 22791 42656 22836 42684
rect 20809 42647 20867 42653
rect 22830 42644 22836 42656
rect 22888 42644 22894 42696
rect 23106 42644 23112 42696
rect 23164 42693 23170 42696
rect 23164 42687 23193 42693
rect 23181 42653 23193 42687
rect 23164 42647 23193 42653
rect 25225 42687 25283 42693
rect 25225 42653 25237 42687
rect 25271 42684 25283 42687
rect 26988 42684 27016 42724
rect 27522 42712 27528 42724
rect 27580 42752 27586 42764
rect 27801 42755 27859 42761
rect 27801 42752 27813 42755
rect 27580 42724 27813 42752
rect 27580 42712 27586 42724
rect 27801 42721 27813 42724
rect 27847 42721 27859 42755
rect 27801 42715 27859 42721
rect 29730 42712 29736 42764
rect 29788 42752 29794 42764
rect 29917 42755 29975 42761
rect 29917 42752 29929 42755
rect 29788 42724 29929 42752
rect 29788 42712 29794 42724
rect 29917 42721 29929 42724
rect 29963 42721 29975 42755
rect 29917 42715 29975 42721
rect 30282 42712 30288 42764
rect 30340 42752 30346 42764
rect 30377 42755 30435 42761
rect 30377 42752 30389 42755
rect 30340 42724 30389 42752
rect 30340 42712 30346 42724
rect 30377 42721 30389 42724
rect 30423 42721 30435 42755
rect 30377 42715 30435 42721
rect 25271 42656 27016 42684
rect 25271 42653 25283 42656
rect 25225 42647 25283 42653
rect 23164 42644 23170 42647
rect 27062 42644 27068 42696
rect 27120 42684 27126 42696
rect 27246 42684 27252 42696
rect 27120 42656 27165 42684
rect 27207 42656 27252 42684
rect 27120 42644 27126 42656
rect 27246 42644 27252 42656
rect 27304 42644 27310 42696
rect 30006 42644 30012 42696
rect 30064 42684 30070 42696
rect 30064 42656 30109 42684
rect 30064 42644 30070 42656
rect 5074 42616 5080 42628
rect 5035 42588 5080 42616
rect 5074 42576 5080 42588
rect 5132 42576 5138 42628
rect 19429 42619 19487 42625
rect 19429 42585 19441 42619
rect 19475 42616 19487 42619
rect 20346 42616 20352 42628
rect 19475 42588 20352 42616
rect 19475 42585 19487 42588
rect 19429 42579 19487 42585
rect 20346 42576 20352 42588
rect 20404 42576 20410 42628
rect 21076 42619 21134 42625
rect 21076 42585 21088 42619
rect 21122 42616 21134 42619
rect 22649 42619 22707 42625
rect 22649 42616 22661 42619
rect 21122 42588 22661 42616
rect 21122 42585 21134 42588
rect 21076 42579 21134 42585
rect 22649 42585 22661 42588
rect 22695 42585 22707 42619
rect 22649 42579 22707 42585
rect 22925 42619 22983 42625
rect 22925 42585 22937 42619
rect 22971 42585 22983 42619
rect 22925 42579 22983 42585
rect 15194 42548 15200 42560
rect 4908 42520 15200 42548
rect 15194 42508 15200 42520
rect 15252 42548 15258 42560
rect 16114 42548 16120 42560
rect 15252 42520 16120 42548
rect 15252 42508 15258 42520
rect 16114 42508 16120 42520
rect 16172 42508 16178 42560
rect 19334 42508 19340 42560
rect 19392 42548 19398 42560
rect 19527 42551 19585 42557
rect 19527 42548 19539 42551
rect 19392 42520 19539 42548
rect 19392 42508 19398 42520
rect 19527 42517 19539 42520
rect 19573 42517 19585 42551
rect 19527 42511 19585 42517
rect 19613 42551 19671 42557
rect 19613 42517 19625 42551
rect 19659 42548 19671 42551
rect 20162 42548 20168 42560
rect 19659 42520 20168 42548
rect 19659 42517 19671 42520
rect 19613 42511 19671 42517
rect 20162 42508 20168 42520
rect 20220 42508 20226 42560
rect 22940 42548 22968 42579
rect 23014 42576 23020 42628
rect 23072 42616 23078 42628
rect 25492 42619 25550 42625
rect 23072 42588 23117 42616
rect 23072 42576 23078 42588
rect 25492 42585 25504 42619
rect 25538 42616 25550 42619
rect 26050 42616 26056 42628
rect 25538 42588 26056 42616
rect 25538 42585 25550 42588
rect 25492 42579 25550 42585
rect 26050 42576 26056 42588
rect 26108 42576 26114 42628
rect 28068 42619 28126 42625
rect 28068 42585 28080 42619
rect 28114 42616 28126 42619
rect 28114 42588 29776 42616
rect 28114 42585 28126 42588
rect 28068 42579 28126 42585
rect 24302 42548 24308 42560
rect 22940 42520 24308 42548
rect 24302 42508 24308 42520
rect 24360 42508 24366 42560
rect 26142 42508 26148 42560
rect 26200 42548 26206 42560
rect 29748 42557 29776 42588
rect 30190 42576 30196 42628
rect 30248 42616 30254 42628
rect 30285 42619 30343 42625
rect 30285 42616 30297 42619
rect 30248 42588 30297 42616
rect 30248 42576 30254 42588
rect 30285 42585 30297 42588
rect 30331 42585 30343 42619
rect 30285 42579 30343 42585
rect 30558 42576 30564 42628
rect 30616 42616 30622 42628
rect 30944 42616 30972 42792
rect 32585 42789 32597 42792
rect 32631 42789 32643 42823
rect 32585 42783 32643 42789
rect 32766 42752 32772 42764
rect 31036 42724 32772 42752
rect 31036 42693 31064 42724
rect 32766 42712 32772 42724
rect 32824 42712 32830 42764
rect 32876 42752 32904 42860
rect 34514 42848 34520 42900
rect 34572 42888 34578 42900
rect 35342 42888 35348 42900
rect 34572 42860 35348 42888
rect 34572 42848 34578 42860
rect 35342 42848 35348 42860
rect 35400 42848 35406 42900
rect 33318 42780 33324 42832
rect 33376 42820 33382 42832
rect 33873 42823 33931 42829
rect 33873 42820 33885 42823
rect 33376 42792 33885 42820
rect 33376 42780 33382 42792
rect 33873 42789 33885 42792
rect 33919 42789 33931 42823
rect 33873 42783 33931 42789
rect 32876 42724 33088 42752
rect 31021 42687 31079 42693
rect 31021 42653 31033 42687
rect 31067 42653 31079 42687
rect 31478 42684 31484 42696
rect 31439 42656 31484 42684
rect 31021 42647 31079 42653
rect 31478 42644 31484 42656
rect 31536 42644 31542 42696
rect 31938 42684 31944 42696
rect 31899 42656 31944 42684
rect 31938 42644 31944 42656
rect 31996 42644 32002 42696
rect 32306 42684 32312 42696
rect 32267 42656 32312 42684
rect 32306 42644 32312 42656
rect 32364 42644 32370 42696
rect 33060 42693 33088 42724
rect 32401 42687 32459 42693
rect 32401 42653 32413 42687
rect 32447 42653 32459 42687
rect 32401 42647 32459 42653
rect 33045 42687 33103 42693
rect 33045 42653 33057 42687
rect 33091 42653 33103 42687
rect 33045 42647 33103 42653
rect 31113 42619 31171 42625
rect 31113 42616 31125 42619
rect 30616 42588 31125 42616
rect 30616 42576 30622 42588
rect 31113 42585 31125 42588
rect 31159 42585 31171 42619
rect 31113 42579 31171 42585
rect 31202 42576 31208 42628
rect 31260 42616 31266 42628
rect 31386 42625 31392 42628
rect 31343 42619 31392 42625
rect 31260 42588 31305 42616
rect 31260 42576 31266 42588
rect 31343 42585 31355 42619
rect 31389 42585 31392 42619
rect 31343 42579 31392 42585
rect 31386 42576 31392 42579
rect 31444 42576 31450 42628
rect 32416 42616 32444 42647
rect 33410 42644 33416 42696
rect 33468 42684 33474 42696
rect 33781 42687 33839 42693
rect 33781 42684 33793 42687
rect 33468 42656 33793 42684
rect 33468 42644 33474 42656
rect 33781 42653 33793 42656
rect 33827 42653 33839 42687
rect 33888 42684 33916 42783
rect 34057 42755 34115 42761
rect 34057 42721 34069 42755
rect 34103 42752 34115 42755
rect 34238 42752 34244 42764
rect 34103 42724 34244 42752
rect 34103 42721 34115 42724
rect 34057 42715 34115 42721
rect 34238 42712 34244 42724
rect 34296 42712 34302 42764
rect 46477 42755 46535 42761
rect 46477 42721 46489 42755
rect 46523 42752 46535 42755
rect 47210 42752 47216 42764
rect 46523 42724 47216 42752
rect 46523 42721 46535 42724
rect 46477 42715 46535 42721
rect 47210 42712 47216 42724
rect 47268 42712 47274 42764
rect 48222 42752 48228 42764
rect 48183 42724 48228 42752
rect 48222 42712 48228 42724
rect 48280 42712 48286 42764
rect 33888 42656 34376 42684
rect 33781 42647 33839 42653
rect 32490 42616 32496 42628
rect 32403 42588 32496 42616
rect 32490 42576 32496 42588
rect 32548 42616 32554 42628
rect 34057 42619 34115 42625
rect 34057 42616 34069 42619
rect 32548 42588 34069 42616
rect 32548 42576 32554 42588
rect 34057 42585 34069 42588
rect 34103 42585 34115 42619
rect 34057 42579 34115 42585
rect 26605 42551 26663 42557
rect 26605 42548 26617 42551
rect 26200 42520 26617 42548
rect 26200 42508 26206 42520
rect 26605 42517 26617 42520
rect 26651 42517 26663 42551
rect 26605 42511 26663 42517
rect 29733 42551 29791 42557
rect 29733 42517 29745 42551
rect 29779 42517 29791 42551
rect 30834 42548 30840 42560
rect 30795 42520 30840 42548
rect 29733 42511 29791 42517
rect 30834 42508 30840 42520
rect 30892 42508 30898 42560
rect 32674 42508 32680 42560
rect 32732 42548 32738 42560
rect 33229 42551 33287 42557
rect 33229 42548 33241 42551
rect 32732 42520 33241 42548
rect 32732 42508 32738 42520
rect 33229 42517 33241 42520
rect 33275 42517 33287 42551
rect 34348 42548 34376 42656
rect 34790 42644 34796 42696
rect 34848 42684 34854 42696
rect 35069 42687 35127 42693
rect 35069 42684 35081 42687
rect 34848 42656 35081 42684
rect 34848 42644 34854 42656
rect 35069 42653 35081 42656
rect 35115 42653 35127 42687
rect 35069 42647 35127 42653
rect 34422 42576 34428 42628
rect 34480 42616 34486 42628
rect 35314 42619 35372 42625
rect 35314 42616 35326 42619
rect 34480 42588 35326 42616
rect 34480 42576 34486 42588
rect 35314 42585 35326 42588
rect 35360 42585 35372 42619
rect 35314 42579 35372 42585
rect 46661 42619 46719 42625
rect 46661 42585 46673 42619
rect 46707 42616 46719 42619
rect 47854 42616 47860 42628
rect 46707 42588 47860 42616
rect 46707 42585 46719 42588
rect 46661 42579 46719 42585
rect 47854 42576 47860 42588
rect 47912 42576 47918 42628
rect 35066 42548 35072 42560
rect 34348 42520 35072 42548
rect 33229 42511 33287 42517
rect 35066 42508 35072 42520
rect 35124 42548 35130 42560
rect 36449 42551 36507 42557
rect 36449 42548 36461 42551
rect 35124 42520 36461 42548
rect 35124 42508 35130 42520
rect 36449 42517 36461 42520
rect 36495 42517 36507 42551
rect 36449 42511 36507 42517
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 5074 42344 5080 42356
rect 5035 42316 5080 42344
rect 5074 42304 5080 42316
rect 5132 42304 5138 42356
rect 16114 42304 16120 42356
rect 16172 42344 16178 42356
rect 17405 42347 17463 42353
rect 16172 42316 17264 42344
rect 16172 42304 16178 42316
rect 13998 42276 14004 42288
rect 6886 42248 14004 42276
rect 4982 42208 4988 42220
rect 4943 42180 4988 42208
rect 4982 42168 4988 42180
rect 5040 42208 5046 42220
rect 6886 42208 6914 42248
rect 13998 42236 14004 42248
rect 14056 42236 14062 42288
rect 5040 42180 6914 42208
rect 15933 42211 15991 42217
rect 5040 42168 5046 42180
rect 15933 42177 15945 42211
rect 15979 42208 15991 42211
rect 17126 42208 17132 42220
rect 15979 42180 16988 42208
rect 17087 42180 17132 42208
rect 15979 42177 15991 42180
rect 15933 42171 15991 42177
rect 16022 42140 16028 42152
rect 15983 42112 16028 42140
rect 16022 42100 16028 42112
rect 16080 42100 16086 42152
rect 16114 42100 16120 42152
rect 16172 42140 16178 42152
rect 16960 42140 16988 42180
rect 17126 42168 17132 42180
rect 17184 42168 17190 42220
rect 17236 42217 17264 42316
rect 17405 42313 17417 42347
rect 17451 42344 17463 42347
rect 19426 42344 19432 42356
rect 17451 42316 19432 42344
rect 17451 42313 17463 42316
rect 17405 42307 17463 42313
rect 19426 42304 19432 42316
rect 19484 42344 19490 42356
rect 19978 42344 19984 42356
rect 19484 42316 19984 42344
rect 19484 42304 19490 42316
rect 19978 42304 19984 42316
rect 20036 42304 20042 42356
rect 20165 42347 20223 42353
rect 20165 42313 20177 42347
rect 20211 42344 20223 42347
rect 20346 42344 20352 42356
rect 20211 42316 20352 42344
rect 20211 42313 20223 42316
rect 20165 42307 20223 42313
rect 20346 42304 20352 42316
rect 20404 42304 20410 42356
rect 22830 42304 22836 42356
rect 22888 42344 22894 42356
rect 23293 42347 23351 42353
rect 23293 42344 23305 42347
rect 22888 42316 23305 42344
rect 22888 42304 22894 42316
rect 23293 42313 23305 42316
rect 23339 42313 23351 42347
rect 24302 42344 24308 42356
rect 24263 42316 24308 42344
rect 23293 42307 23351 42313
rect 24302 42304 24308 42316
rect 24360 42304 24366 42356
rect 25133 42347 25191 42353
rect 25133 42313 25145 42347
rect 25179 42344 25191 42347
rect 25498 42344 25504 42356
rect 25179 42316 25504 42344
rect 25179 42313 25191 42316
rect 25133 42307 25191 42313
rect 25498 42304 25504 42316
rect 25556 42304 25562 42356
rect 30466 42304 30472 42356
rect 30524 42344 30530 42356
rect 30653 42347 30711 42353
rect 30653 42344 30665 42347
rect 30524 42316 30665 42344
rect 30524 42304 30530 42316
rect 30653 42313 30665 42316
rect 30699 42313 30711 42347
rect 32674 42344 32680 42356
rect 32635 42316 32680 42344
rect 30653 42307 30711 42313
rect 32674 42304 32680 42316
rect 32732 42304 32738 42356
rect 34422 42344 34428 42356
rect 34383 42316 34428 42344
rect 34422 42304 34428 42316
rect 34480 42304 34486 42356
rect 35526 42344 35532 42356
rect 34808 42316 35532 42344
rect 28994 42276 29000 42288
rect 23676 42248 24532 42276
rect 23676 42220 23704 42248
rect 17221 42211 17279 42217
rect 17221 42177 17233 42211
rect 17267 42177 17279 42211
rect 17221 42171 17279 42177
rect 19052 42211 19110 42217
rect 19052 42177 19064 42211
rect 19098 42208 19110 42211
rect 19426 42208 19432 42220
rect 19098 42180 19432 42208
rect 19098 42177 19110 42180
rect 19052 42171 19110 42177
rect 19426 42168 19432 42180
rect 19484 42168 19490 42220
rect 22094 42168 22100 42220
rect 22152 42208 22158 42220
rect 22465 42211 22523 42217
rect 22465 42208 22477 42211
rect 22152 42180 22477 42208
rect 22152 42168 22158 42180
rect 22465 42177 22477 42180
rect 22511 42177 22523 42211
rect 23477 42211 23535 42217
rect 23477 42208 23489 42211
rect 22465 42171 22523 42177
rect 23400 42180 23489 42208
rect 17678 42140 17684 42152
rect 16172 42112 16217 42140
rect 16960 42112 17684 42140
rect 16172 42100 16178 42112
rect 17678 42100 17684 42112
rect 17736 42100 17742 42152
rect 18785 42143 18843 42149
rect 18785 42109 18797 42143
rect 18831 42109 18843 42143
rect 22554 42140 22560 42152
rect 22515 42112 22560 42140
rect 18785 42103 18843 42109
rect 15470 42032 15476 42084
rect 15528 42072 15534 42084
rect 18800 42072 18828 42103
rect 22554 42100 22560 42112
rect 22612 42100 22618 42152
rect 20622 42072 20628 42084
rect 15528 42044 18828 42072
rect 15528 42032 15534 42044
rect 14918 41964 14924 42016
rect 14976 42004 14982 42016
rect 15565 42007 15623 42013
rect 15565 42004 15577 42007
rect 14976 41976 15577 42004
rect 14976 41964 14982 41976
rect 15565 41973 15577 41976
rect 15611 41973 15623 42007
rect 18800 42004 18828 42044
rect 20088 42044 20628 42072
rect 20088 42004 20116 42044
rect 20622 42032 20628 42044
rect 20680 42032 20686 42084
rect 22833 42075 22891 42081
rect 22833 42041 22845 42075
rect 22879 42072 22891 42075
rect 23400 42072 23428 42180
rect 23477 42177 23489 42180
rect 23523 42177 23535 42211
rect 23658 42208 23664 42220
rect 23619 42180 23664 42208
rect 23477 42171 23535 42177
rect 23658 42168 23664 42180
rect 23716 42168 23722 42220
rect 23753 42211 23811 42217
rect 23753 42177 23765 42211
rect 23799 42177 23811 42211
rect 24210 42208 24216 42220
rect 24171 42180 24216 42208
rect 23753 42171 23811 42177
rect 23768 42140 23796 42171
rect 24210 42168 24216 42180
rect 24268 42168 24274 42220
rect 24504 42217 24532 42248
rect 26252 42248 29000 42276
rect 24397 42211 24455 42217
rect 24397 42177 24409 42211
rect 24443 42177 24455 42211
rect 24397 42171 24455 42177
rect 24489 42211 24547 42217
rect 24489 42177 24501 42211
rect 24535 42177 24547 42211
rect 24489 42171 24547 42177
rect 24412 42140 24440 42171
rect 24670 42168 24676 42220
rect 24728 42208 24734 42220
rect 26252 42217 26280 42248
rect 28994 42236 29000 42248
rect 29052 42236 29058 42288
rect 29540 42279 29598 42285
rect 29540 42245 29552 42279
rect 29586 42276 29598 42279
rect 30834 42276 30840 42288
rect 29586 42248 30840 42276
rect 29586 42245 29598 42248
rect 29540 42239 29598 42245
rect 30834 42236 30840 42248
rect 30892 42236 30898 42288
rect 31481 42279 31539 42285
rect 31481 42245 31493 42279
rect 31527 42276 31539 42279
rect 31938 42276 31944 42288
rect 31527 42248 31944 42276
rect 31527 42245 31539 42248
rect 31481 42239 31539 42245
rect 31938 42236 31944 42248
rect 31996 42276 32002 42288
rect 32585 42279 32643 42285
rect 32585 42276 32597 42279
rect 31996 42248 32597 42276
rect 31996 42236 32002 42248
rect 32585 42245 32597 42248
rect 32631 42245 32643 42279
rect 32585 42239 32643 42245
rect 33965 42279 34023 42285
rect 33965 42245 33977 42279
rect 34011 42276 34023 42279
rect 34514 42276 34520 42288
rect 34011 42248 34520 42276
rect 34011 42245 34023 42248
rect 33965 42239 34023 42245
rect 34514 42236 34520 42248
rect 34572 42236 34578 42288
rect 34722 42279 34780 42285
rect 34722 42245 34734 42279
rect 34768 42276 34780 42279
rect 34808 42276 34836 42316
rect 35526 42304 35532 42316
rect 35584 42304 35590 42356
rect 34768 42248 34836 42276
rect 34768 42245 34780 42248
rect 34722 42239 34780 42245
rect 25317 42211 25375 42217
rect 25317 42208 25329 42211
rect 24728 42180 25329 42208
rect 24728 42168 24734 42180
rect 25317 42177 25329 42180
rect 25363 42177 25375 42211
rect 25317 42171 25375 42177
rect 26237 42211 26295 42217
rect 26237 42177 26249 42211
rect 26283 42177 26295 42211
rect 27157 42211 27215 42217
rect 27157 42208 27169 42211
rect 26237 42171 26295 42177
rect 26620 42180 27169 42208
rect 23492 42112 24440 42140
rect 25593 42143 25651 42149
rect 23492 42084 23520 42112
rect 25593 42109 25605 42143
rect 25639 42109 25651 42143
rect 26142 42140 26148 42152
rect 26103 42112 26148 42140
rect 25593 42103 25651 42109
rect 22879 42044 23428 42072
rect 22879 42041 22891 42044
rect 22833 42035 22891 42041
rect 18800 41976 20116 42004
rect 15565 41967 15623 41973
rect 20990 41964 20996 42016
rect 21048 42004 21054 42016
rect 23198 42004 23204 42016
rect 21048 41976 23204 42004
rect 21048 41964 21054 41976
rect 23198 41964 23204 41976
rect 23256 41964 23262 42016
rect 23400 42004 23428 42044
rect 23474 42032 23480 42084
rect 23532 42032 23538 42084
rect 25608 42072 25636 42103
rect 26142 42100 26148 42112
rect 26200 42100 26206 42152
rect 26620 42081 26648 42180
rect 27157 42177 27169 42180
rect 27203 42208 27215 42211
rect 27246 42208 27252 42220
rect 27203 42180 27252 42208
rect 27203 42177 27215 42180
rect 27157 42171 27215 42177
rect 27246 42168 27252 42180
rect 27304 42168 27310 42220
rect 27522 42168 27528 42220
rect 27580 42208 27586 42220
rect 29273 42211 29331 42217
rect 29273 42208 29285 42211
rect 27580 42180 29285 42208
rect 27580 42168 27586 42180
rect 29273 42177 29285 42180
rect 29319 42177 29331 42211
rect 31110 42208 31116 42220
rect 31071 42180 31116 42208
rect 29273 42171 29331 42177
rect 31110 42168 31116 42180
rect 31168 42168 31174 42220
rect 31294 42208 31300 42220
rect 31255 42180 31300 42208
rect 31294 42168 31300 42180
rect 31352 42168 31358 42220
rect 32122 42208 32128 42220
rect 31404 42180 32128 42208
rect 31202 42100 31208 42152
rect 31260 42140 31266 42152
rect 31404 42140 31432 42180
rect 32122 42168 32128 42180
rect 32180 42168 32186 42220
rect 32490 42208 32496 42220
rect 32451 42180 32496 42208
rect 32490 42168 32496 42180
rect 32548 42168 32554 42220
rect 32674 42168 32680 42220
rect 32732 42208 32738 42220
rect 33318 42208 33324 42220
rect 32732 42180 33324 42208
rect 32732 42168 32738 42180
rect 33318 42168 33324 42180
rect 33376 42168 33382 42220
rect 33410 42168 33416 42220
rect 33468 42208 33474 42220
rect 33781 42211 33839 42217
rect 33781 42208 33793 42211
rect 33468 42180 33793 42208
rect 33468 42168 33474 42180
rect 33781 42177 33793 42180
rect 33827 42208 33839 42211
rect 34606 42208 34612 42220
rect 33827 42180 34376 42208
rect 34567 42180 34612 42208
rect 33827 42177 33839 42180
rect 33781 42171 33839 42177
rect 33597 42143 33655 42149
rect 33597 42140 33609 42143
rect 31260 42112 31432 42140
rect 31726 42112 33609 42140
rect 31260 42100 31266 42112
rect 26605 42075 26663 42081
rect 26605 42072 26617 42075
rect 25608 42044 26617 42072
rect 26605 42041 26617 42044
rect 26651 42041 26663 42075
rect 26605 42035 26663 42041
rect 30374 42032 30380 42084
rect 30432 42072 30438 42084
rect 31386 42072 31392 42084
rect 30432 42044 31392 42072
rect 30432 42032 30438 42044
rect 31386 42032 31392 42044
rect 31444 42032 31450 42084
rect 24210 42004 24216 42016
rect 23400 41976 24216 42004
rect 24210 41964 24216 41976
rect 24268 41964 24274 42016
rect 25501 42007 25559 42013
rect 25501 41973 25513 42007
rect 25547 42004 25559 42007
rect 27062 42004 27068 42016
rect 25547 41976 27068 42004
rect 25547 41973 25559 41976
rect 25501 41967 25559 41973
rect 27062 41964 27068 41976
rect 27120 41964 27126 42016
rect 27154 41964 27160 42016
rect 27212 42004 27218 42016
rect 27249 42007 27307 42013
rect 27249 42004 27261 42007
rect 27212 41976 27261 42004
rect 27212 41964 27218 41976
rect 27249 41973 27261 41976
rect 27295 41973 27307 42007
rect 27249 41967 27307 41973
rect 31018 41964 31024 42016
rect 31076 42004 31082 42016
rect 31726 42004 31754 42112
rect 33597 42109 33609 42112
rect 33643 42140 33655 42143
rect 33686 42140 33692 42152
rect 33643 42112 33692 42140
rect 33643 42109 33655 42112
rect 33597 42103 33655 42109
rect 33686 42100 33692 42112
rect 33744 42100 33750 42152
rect 32309 42075 32367 42081
rect 32309 42041 32321 42075
rect 32355 42072 32367 42075
rect 34348 42072 34376 42180
rect 34606 42168 34612 42180
rect 34664 42168 34670 42220
rect 34806 42211 34864 42217
rect 34806 42177 34818 42211
rect 34852 42177 34864 42211
rect 34911 42211 34969 42217
rect 34911 42208 34923 42211
rect 34806 42171 34864 42177
rect 34900 42177 34923 42208
rect 34957 42177 34969 42211
rect 34900 42171 34969 42177
rect 34422 42100 34428 42152
rect 34480 42140 34486 42152
rect 34808 42140 34836 42171
rect 34480 42112 34836 42140
rect 34480 42100 34486 42112
rect 34514 42072 34520 42084
rect 32355 42044 34192 42072
rect 34348 42044 34520 42072
rect 32355 42041 32367 42044
rect 32309 42035 32367 42041
rect 34164 42016 34192 42044
rect 34514 42032 34520 42044
rect 34572 42032 34578 42084
rect 34606 42032 34612 42084
rect 34664 42072 34670 42084
rect 34900 42072 34928 42171
rect 35066 42168 35072 42220
rect 35124 42208 35130 42220
rect 35124 42180 35169 42208
rect 35124 42168 35130 42180
rect 35342 42168 35348 42220
rect 35400 42208 35406 42220
rect 35529 42211 35587 42217
rect 35529 42208 35541 42211
rect 35400 42180 35541 42208
rect 35400 42168 35406 42180
rect 35529 42177 35541 42180
rect 35575 42177 35587 42211
rect 35710 42208 35716 42220
rect 35671 42180 35716 42208
rect 35529 42171 35587 42177
rect 35710 42168 35716 42180
rect 35768 42168 35774 42220
rect 47762 42208 47768 42220
rect 47723 42180 47768 42208
rect 47762 42168 47768 42180
rect 47820 42168 47826 42220
rect 34664 42044 34928 42072
rect 34664 42032 34670 42044
rect 31076 41976 31754 42004
rect 31076 41964 31082 41976
rect 32030 41964 32036 42016
rect 32088 42004 32094 42016
rect 32674 42004 32680 42016
rect 32088 41976 32680 42004
rect 32088 41964 32094 41976
rect 32674 41964 32680 41976
rect 32732 41964 32738 42016
rect 32858 42004 32864 42016
rect 32819 41976 32864 42004
rect 32858 41964 32864 41976
rect 32916 41964 32922 42016
rect 34146 41964 34152 42016
rect 34204 42004 34210 42016
rect 35529 42007 35587 42013
rect 35529 42004 35541 42007
rect 34204 41976 35541 42004
rect 34204 41964 34210 41976
rect 35529 41973 35541 41976
rect 35575 41973 35587 42007
rect 35529 41967 35587 41973
rect 46474 41964 46480 42016
rect 46532 42004 46538 42016
rect 47213 42007 47271 42013
rect 47213 42004 47225 42007
rect 46532 41976 47225 42004
rect 46532 41964 46538 41976
rect 47213 41973 47225 41976
rect 47259 41973 47271 42007
rect 47854 42004 47860 42016
rect 47815 41976 47860 42004
rect 47213 41967 47271 41973
rect 47854 41964 47860 41976
rect 47912 41964 47918 42016
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 16853 41803 16911 41809
rect 16853 41769 16865 41803
rect 16899 41800 16911 41803
rect 17126 41800 17132 41812
rect 16899 41772 17132 41800
rect 16899 41769 16911 41772
rect 16853 41763 16911 41769
rect 17126 41760 17132 41772
rect 17184 41760 17190 41812
rect 17494 41800 17500 41812
rect 17455 41772 17500 41800
rect 17494 41760 17500 41772
rect 17552 41760 17558 41812
rect 17678 41800 17684 41812
rect 17639 41772 17684 41800
rect 17678 41760 17684 41772
rect 17736 41760 17742 41812
rect 19426 41800 19432 41812
rect 19387 41772 19432 41800
rect 19426 41760 19432 41772
rect 19484 41760 19490 41812
rect 21913 41803 21971 41809
rect 21913 41769 21925 41803
rect 21959 41800 21971 41803
rect 22554 41800 22560 41812
rect 21959 41772 22560 41800
rect 21959 41769 21971 41772
rect 21913 41763 21971 41769
rect 22554 41760 22560 41772
rect 22612 41760 22618 41812
rect 23198 41760 23204 41812
rect 23256 41800 23262 41812
rect 30098 41800 30104 41812
rect 23256 41772 30104 41800
rect 23256 41760 23262 41772
rect 30098 41760 30104 41772
rect 30156 41760 30162 41812
rect 30282 41760 30288 41812
rect 30340 41800 30346 41812
rect 31113 41803 31171 41809
rect 31113 41800 31125 41803
rect 30340 41772 31125 41800
rect 30340 41760 30346 41772
rect 31113 41769 31125 41772
rect 31159 41769 31171 41803
rect 31113 41763 31171 41769
rect 31205 41803 31263 41809
rect 31205 41769 31217 41803
rect 31251 41800 31263 41803
rect 31478 41800 31484 41812
rect 31251 41772 31484 41800
rect 31251 41769 31263 41772
rect 31205 41763 31263 41769
rect 31478 41760 31484 41772
rect 31536 41760 31542 41812
rect 32306 41760 32312 41812
rect 32364 41800 32370 41812
rect 33045 41803 33103 41809
rect 33045 41800 33057 41803
rect 32364 41772 33057 41800
rect 32364 41760 32370 41772
rect 33045 41769 33057 41772
rect 33091 41769 33103 41803
rect 33045 41763 33103 41769
rect 34054 41760 34060 41812
rect 34112 41800 34118 41812
rect 35069 41803 35127 41809
rect 35069 41800 35081 41803
rect 34112 41772 35081 41800
rect 34112 41760 34118 41772
rect 35069 41769 35081 41772
rect 35115 41800 35127 41803
rect 35434 41800 35440 41812
rect 35115 41772 35440 41800
rect 35115 41769 35127 41772
rect 35069 41763 35127 41769
rect 35434 41760 35440 41772
rect 35492 41760 35498 41812
rect 17402 41692 17408 41744
rect 17460 41732 17466 41744
rect 20162 41732 20168 41744
rect 17460 41704 20168 41732
rect 17460 41692 17466 41704
rect 20162 41692 20168 41704
rect 20220 41732 20226 41744
rect 23293 41735 23351 41741
rect 23293 41732 23305 41735
rect 20220 41704 23305 41732
rect 20220 41692 20226 41704
rect 15470 41664 15476 41676
rect 15431 41636 15476 41664
rect 15470 41624 15476 41636
rect 15528 41624 15534 41676
rect 19334 41624 19340 41676
rect 19392 41664 19398 41676
rect 19613 41667 19671 41673
rect 19613 41664 19625 41667
rect 19392 41636 19625 41664
rect 19392 41624 19398 41636
rect 19613 41633 19625 41636
rect 19659 41633 19671 41667
rect 20070 41664 20076 41676
rect 19983 41636 20076 41664
rect 19613 41627 19671 41633
rect 20070 41624 20076 41636
rect 20128 41664 20134 41676
rect 20346 41664 20352 41676
rect 20128 41636 20352 41664
rect 20128 41624 20134 41636
rect 20346 41624 20352 41636
rect 20404 41624 20410 41676
rect 20824 41673 20852 41704
rect 23293 41701 23305 41704
rect 23339 41701 23351 41735
rect 25593 41735 25651 41741
rect 25593 41732 25605 41735
rect 23293 41695 23351 41701
rect 25056 41704 25605 41732
rect 20809 41667 20867 41673
rect 20809 41633 20821 41667
rect 20855 41633 20867 41667
rect 20990 41664 20996 41676
rect 20951 41636 20996 41664
rect 20809 41627 20867 41633
rect 20990 41624 20996 41636
rect 21048 41624 21054 41676
rect 22094 41624 22100 41676
rect 22152 41664 22158 41676
rect 24949 41667 25007 41673
rect 24949 41664 24961 41667
rect 22152 41636 22197 41664
rect 23124 41636 24961 41664
rect 22152 41624 22158 41636
rect 2038 41556 2044 41608
rect 2096 41596 2102 41608
rect 2225 41599 2283 41605
rect 2225 41596 2237 41599
rect 2096 41568 2237 41596
rect 2096 41556 2102 41568
rect 2225 41565 2237 41568
rect 2271 41565 2283 41599
rect 14918 41596 14924 41608
rect 14879 41568 14924 41596
rect 2225 41559 2283 41565
rect 14918 41556 14924 41568
rect 14976 41556 14982 41608
rect 19705 41599 19763 41605
rect 19705 41565 19717 41599
rect 19751 41565 19763 41599
rect 19705 41559 19763 41565
rect 19981 41599 20039 41605
rect 19981 41565 19993 41599
rect 20027 41596 20039 41599
rect 20254 41596 20260 41608
rect 20027 41568 20260 41596
rect 20027 41565 20039 41568
rect 19981 41559 20039 41565
rect 15740 41531 15798 41537
rect 15740 41497 15752 41531
rect 15786 41528 15798 41531
rect 15930 41528 15936 41540
rect 15786 41500 15936 41528
rect 15786 41497 15798 41500
rect 15740 41491 15798 41497
rect 15930 41488 15936 41500
rect 15988 41488 15994 41540
rect 17126 41488 17132 41540
rect 17184 41528 17190 41540
rect 17313 41531 17371 41537
rect 17313 41528 17325 41531
rect 17184 41500 17325 41528
rect 17184 41488 17190 41500
rect 17313 41497 17325 41500
rect 17359 41497 17371 41531
rect 17313 41491 17371 41497
rect 14734 41460 14740 41472
rect 14695 41432 14740 41460
rect 14734 41420 14740 41432
rect 14792 41420 14798 41472
rect 17402 41420 17408 41472
rect 17460 41460 17466 41472
rect 17513 41463 17571 41469
rect 17513 41460 17525 41463
rect 17460 41432 17525 41460
rect 17460 41420 17466 41432
rect 17513 41429 17525 41432
rect 17559 41429 17571 41463
rect 17513 41423 17571 41429
rect 19426 41420 19432 41472
rect 19484 41460 19490 41472
rect 19720 41460 19748 41559
rect 20254 41556 20260 41568
rect 20312 41556 20318 41608
rect 20364 41528 20392 41624
rect 20530 41556 20536 41608
rect 20588 41596 20594 41608
rect 20717 41599 20775 41605
rect 20717 41596 20729 41599
rect 20588 41568 20729 41596
rect 20588 41556 20594 41568
rect 20717 41565 20729 41568
rect 20763 41565 20775 41599
rect 20717 41559 20775 41565
rect 20901 41599 20959 41605
rect 20901 41565 20913 41599
rect 20947 41565 20959 41599
rect 21818 41596 21824 41608
rect 21779 41568 21824 41596
rect 20901 41559 20959 41565
rect 20916 41528 20944 41559
rect 21818 41556 21824 41568
rect 21876 41556 21882 41608
rect 23124 41605 23152 41636
rect 24949 41633 24961 41636
rect 24995 41633 25007 41667
rect 24949 41627 25007 41633
rect 23109 41599 23167 41605
rect 23109 41565 23121 41599
rect 23155 41565 23167 41599
rect 23109 41559 23167 41565
rect 23201 41599 23259 41605
rect 23201 41565 23213 41599
rect 23247 41596 23259 41599
rect 23290 41596 23296 41608
rect 23247 41568 23296 41596
rect 23247 41565 23259 41568
rect 23201 41559 23259 41565
rect 23290 41556 23296 41568
rect 23348 41556 23354 41608
rect 23385 41599 23443 41605
rect 23385 41565 23397 41599
rect 23431 41565 23443 41599
rect 23385 41559 23443 41565
rect 23753 41599 23811 41605
rect 23753 41565 23765 41599
rect 23799 41596 23811 41599
rect 24118 41596 24124 41608
rect 23799 41568 24124 41596
rect 23799 41565 23811 41568
rect 23753 41559 23811 41565
rect 20364 41500 20944 41528
rect 22097 41531 22155 41537
rect 22097 41497 22109 41531
rect 22143 41528 22155 41531
rect 23400 41528 23428 41559
rect 24118 41556 24124 41568
rect 24176 41596 24182 41608
rect 25056 41596 25084 41704
rect 25593 41701 25605 41704
rect 25639 41701 25651 41735
rect 25593 41695 25651 41701
rect 31297 41735 31355 41741
rect 31297 41701 31309 41735
rect 31343 41732 31355 41735
rect 32030 41732 32036 41744
rect 31343 41704 32036 41732
rect 31343 41701 31355 41704
rect 31297 41695 31355 41701
rect 32030 41692 32036 41704
rect 32088 41692 32094 41744
rect 32122 41692 32128 41744
rect 32180 41732 32186 41744
rect 34422 41732 34428 41744
rect 32180 41704 34428 41732
rect 32180 41692 32186 41704
rect 34422 41692 34428 41704
rect 34480 41692 34486 41744
rect 35253 41735 35311 41741
rect 35253 41701 35265 41735
rect 35299 41732 35311 41735
rect 35526 41732 35532 41744
rect 35299 41704 35532 41732
rect 35299 41701 35311 41704
rect 35253 41695 35311 41701
rect 35526 41692 35532 41704
rect 35584 41692 35590 41744
rect 26142 41664 26148 41676
rect 25608 41636 26148 41664
rect 25608 41605 25636 41636
rect 26142 41624 26148 41636
rect 26200 41624 26206 41676
rect 29454 41664 29460 41676
rect 26896 41636 29460 41664
rect 24176 41568 25084 41596
rect 25593 41599 25651 41605
rect 24176 41556 24182 41568
rect 25593 41565 25605 41599
rect 25639 41565 25651 41599
rect 25774 41596 25780 41608
rect 25735 41568 25780 41596
rect 25593 41559 25651 41565
rect 25774 41556 25780 41568
rect 25832 41556 25838 41608
rect 26896 41605 26924 41636
rect 29454 41624 29460 41636
rect 29512 41624 29518 41676
rect 33410 41664 33416 41676
rect 31726 41636 33416 41664
rect 26789 41599 26847 41605
rect 26789 41565 26801 41599
rect 26835 41565 26847 41599
rect 26789 41559 26847 41565
rect 26881 41599 26939 41605
rect 26881 41565 26893 41599
rect 26927 41565 26939 41599
rect 26881 41559 26939 41565
rect 22143 41500 23428 41528
rect 22143 41497 22155 41500
rect 22097 41491 22155 41497
rect 24210 41488 24216 41540
rect 24268 41528 24274 41540
rect 24581 41531 24639 41537
rect 24581 41528 24593 41531
rect 24268 41500 24593 41528
rect 24268 41488 24274 41500
rect 24581 41497 24593 41500
rect 24627 41497 24639 41531
rect 24762 41528 24768 41540
rect 24723 41500 24768 41528
rect 24581 41491 24639 41497
rect 24762 41488 24768 41500
rect 24820 41488 24826 41540
rect 25958 41488 25964 41540
rect 26016 41528 26022 41540
rect 26804 41528 26832 41559
rect 26970 41556 26976 41608
rect 27028 41596 27034 41608
rect 27065 41599 27123 41605
rect 27065 41596 27077 41599
rect 27028 41568 27077 41596
rect 27028 41556 27034 41568
rect 27065 41565 27077 41568
rect 27111 41565 27123 41599
rect 27065 41559 27123 41565
rect 27154 41556 27160 41608
rect 27212 41596 27218 41608
rect 27212 41568 27257 41596
rect 27212 41556 27218 41568
rect 30742 41556 30748 41608
rect 30800 41596 30806 41608
rect 31018 41596 31024 41608
rect 30800 41568 31024 41596
rect 30800 41556 30806 41568
rect 31018 41556 31024 41568
rect 31076 41556 31082 41608
rect 31481 41599 31539 41605
rect 31481 41565 31493 41599
rect 31527 41596 31539 41599
rect 31726 41596 31754 41636
rect 33410 41624 33416 41636
rect 33468 41664 33474 41676
rect 33689 41667 33747 41673
rect 33468 41636 33640 41664
rect 33468 41624 33474 41636
rect 31527 41568 31754 41596
rect 31527 41565 31539 41568
rect 31481 41559 31539 41565
rect 32490 41556 32496 41608
rect 32548 41596 32554 41608
rect 33612 41605 33640 41636
rect 33689 41633 33701 41667
rect 33735 41664 33747 41667
rect 35710 41664 35716 41676
rect 33735 41636 35716 41664
rect 33735 41633 33747 41636
rect 33689 41627 33747 41633
rect 35710 41624 35716 41636
rect 35768 41624 35774 41676
rect 46474 41664 46480 41676
rect 46435 41636 46480 41664
rect 46474 41624 46480 41636
rect 46532 41624 46538 41676
rect 46661 41667 46719 41673
rect 46661 41633 46673 41667
rect 46707 41664 46719 41667
rect 47854 41664 47860 41676
rect 46707 41636 47860 41664
rect 46707 41633 46719 41636
rect 46661 41627 46719 41633
rect 47854 41624 47860 41636
rect 47912 41624 47918 41676
rect 48222 41664 48228 41676
rect 48183 41636 48228 41664
rect 48222 41624 48228 41636
rect 48280 41624 48286 41676
rect 32953 41599 33011 41605
rect 32953 41596 32965 41599
rect 32548 41568 32965 41596
rect 32548 41556 32554 41568
rect 32953 41565 32965 41568
rect 32999 41596 33011 41599
rect 33137 41599 33195 41605
rect 32999 41568 33088 41596
rect 32999 41565 33011 41568
rect 32953 41559 33011 41565
rect 27798 41528 27804 41540
rect 26016 41500 26061 41528
rect 26804 41500 27804 41528
rect 26016 41488 26022 41500
rect 27798 41488 27804 41500
rect 27856 41488 27862 41540
rect 20533 41463 20591 41469
rect 20533 41460 20545 41463
rect 19484 41432 20545 41460
rect 19484 41420 19490 41432
rect 20533 41429 20545 41432
rect 20579 41429 20591 41463
rect 20533 41423 20591 41429
rect 24302 41420 24308 41472
rect 24360 41460 24366 41472
rect 26605 41463 26663 41469
rect 26605 41460 26617 41463
rect 24360 41432 26617 41460
rect 24360 41420 24366 41432
rect 26605 41429 26617 41432
rect 26651 41429 26663 41463
rect 26605 41423 26663 41429
rect 30745 41463 30803 41469
rect 30745 41429 30757 41463
rect 30791 41460 30803 41463
rect 30926 41460 30932 41472
rect 30791 41432 30932 41460
rect 30791 41429 30803 41432
rect 30745 41423 30803 41429
rect 30926 41420 30932 41432
rect 30984 41420 30990 41472
rect 33060 41460 33088 41568
rect 33137 41565 33149 41599
rect 33183 41565 33195 41599
rect 33137 41559 33195 41565
rect 33597 41599 33655 41605
rect 33597 41565 33609 41599
rect 33643 41565 33655 41599
rect 33778 41596 33784 41608
rect 33739 41568 33784 41596
rect 33597 41559 33655 41565
rect 33152 41528 33180 41559
rect 33778 41556 33784 41568
rect 33836 41556 33842 41608
rect 34698 41556 34704 41608
rect 34756 41596 34762 41608
rect 34885 41599 34943 41605
rect 34885 41596 34897 41599
rect 34756 41568 34897 41596
rect 34756 41556 34762 41568
rect 34885 41565 34897 41568
rect 34931 41565 34943 41599
rect 34885 41559 34943 41565
rect 35069 41599 35127 41605
rect 35069 41565 35081 41599
rect 35115 41596 35127 41599
rect 35342 41596 35348 41608
rect 35115 41568 35348 41596
rect 35115 41565 35127 41568
rect 35069 41559 35127 41565
rect 35342 41556 35348 41568
rect 35400 41556 35406 41608
rect 46014 41596 46020 41608
rect 45975 41568 46020 41596
rect 46014 41556 46020 41568
rect 46072 41556 46078 41608
rect 34054 41528 34060 41540
rect 33152 41500 34060 41528
rect 34054 41488 34060 41500
rect 34112 41488 34118 41540
rect 34716 41460 34744 41556
rect 33060 41432 34744 41460
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 15194 41216 15200 41268
rect 15252 41256 15258 41268
rect 15473 41259 15531 41265
rect 15473 41256 15485 41259
rect 15252 41228 15485 41256
rect 15252 41216 15258 41228
rect 15473 41225 15485 41228
rect 15519 41225 15531 41259
rect 15473 41219 15531 41225
rect 19521 41259 19579 41265
rect 19521 41225 19533 41259
rect 19567 41256 19579 41259
rect 20162 41256 20168 41268
rect 19567 41228 20168 41256
rect 19567 41225 19579 41228
rect 19521 41219 19579 41225
rect 20162 41216 20168 41228
rect 20220 41216 20226 41268
rect 23290 41216 23296 41268
rect 23348 41256 23354 41268
rect 23569 41259 23627 41265
rect 23569 41256 23581 41259
rect 23348 41228 23581 41256
rect 23348 41216 23354 41228
rect 23569 41225 23581 41228
rect 23615 41256 23627 41259
rect 24302 41256 24308 41268
rect 23615 41228 24308 41256
rect 23615 41225 23627 41228
rect 23569 41219 23627 41225
rect 24302 41216 24308 41228
rect 24360 41216 24366 41268
rect 27062 41216 27068 41268
rect 27120 41256 27126 41268
rect 27157 41259 27215 41265
rect 27157 41256 27169 41259
rect 27120 41228 27169 41256
rect 27120 41216 27126 41228
rect 27157 41225 27169 41228
rect 27203 41225 27215 41259
rect 27157 41219 27215 41225
rect 30098 41216 30104 41268
rect 30156 41256 30162 41268
rect 31202 41256 31208 41268
rect 30156 41228 31208 41256
rect 30156 41216 30162 41228
rect 31202 41216 31208 41228
rect 31260 41216 31266 41268
rect 33873 41259 33931 41265
rect 33873 41225 33885 41259
rect 33919 41225 33931 41259
rect 33873 41219 33931 41225
rect 14360 41191 14418 41197
rect 14360 41157 14372 41191
rect 14406 41188 14418 41191
rect 14734 41188 14740 41200
rect 14406 41160 14740 41188
rect 14406 41157 14418 41160
rect 14360 41151 14418 41157
rect 14734 41148 14740 41160
rect 14792 41148 14798 41200
rect 19245 41191 19303 41197
rect 19245 41157 19257 41191
rect 19291 41188 19303 41191
rect 20070 41188 20076 41200
rect 19291 41160 20076 41188
rect 19291 41157 19303 41160
rect 19245 41151 19303 41157
rect 20070 41148 20076 41160
rect 20128 41148 20134 41200
rect 20530 41188 20536 41200
rect 20180 41160 20536 41188
rect 2038 41120 2044 41132
rect 1999 41092 2044 41120
rect 2038 41080 2044 41092
rect 2096 41080 2102 41132
rect 16022 41120 16028 41132
rect 15983 41092 16028 41120
rect 16022 41080 16028 41092
rect 16080 41080 16086 41132
rect 16117 41123 16175 41129
rect 16117 41089 16129 41123
rect 16163 41120 16175 41123
rect 16853 41123 16911 41129
rect 16853 41120 16865 41123
rect 16163 41092 16865 41120
rect 16163 41089 16175 41092
rect 16117 41083 16175 41089
rect 16853 41089 16865 41092
rect 16899 41089 16911 41123
rect 17034 41120 17040 41132
rect 16995 41092 17040 41120
rect 16853 41083 16911 41089
rect 17034 41080 17040 41092
rect 17092 41080 17098 41132
rect 17221 41123 17279 41129
rect 17221 41089 17233 41123
rect 17267 41089 17279 41123
rect 17221 41083 17279 41089
rect 2225 41055 2283 41061
rect 2225 41021 2237 41055
rect 2271 41052 2283 41055
rect 2314 41052 2320 41064
rect 2271 41024 2320 41052
rect 2271 41021 2283 41024
rect 2225 41015 2283 41021
rect 2314 41012 2320 41024
rect 2372 41012 2378 41064
rect 2774 41052 2780 41064
rect 2735 41024 2780 41052
rect 2774 41012 2780 41024
rect 2832 41012 2838 41064
rect 14090 41052 14096 41064
rect 14051 41024 14096 41052
rect 14090 41012 14096 41024
rect 14148 41012 14154 41064
rect 17236 41052 17264 41083
rect 17310 41080 17316 41132
rect 17368 41120 17374 41132
rect 19429 41123 19487 41129
rect 17368 41092 17413 41120
rect 17368 41080 17374 41092
rect 19429 41089 19441 41123
rect 19475 41089 19487 41123
rect 19429 41083 19487 41089
rect 19613 41123 19671 41129
rect 19613 41089 19625 41123
rect 19659 41120 19671 41123
rect 19978 41120 19984 41132
rect 19659 41092 19984 41120
rect 19659 41089 19671 41092
rect 19613 41083 19671 41089
rect 17494 41052 17500 41064
rect 17236 41024 17500 41052
rect 17494 41012 17500 41024
rect 17552 41052 17558 41064
rect 19242 41052 19248 41064
rect 17552 41024 19248 41052
rect 17552 41012 17558 41024
rect 19242 41012 19248 41024
rect 19300 41052 19306 41064
rect 19444 41052 19472 41083
rect 19978 41080 19984 41092
rect 20036 41120 20042 41132
rect 20180 41120 20208 41160
rect 20530 41148 20536 41160
rect 20588 41148 20594 41200
rect 21818 41148 21824 41200
rect 21876 41188 21882 41200
rect 22373 41191 22431 41197
rect 22373 41188 22385 41191
rect 21876 41160 22385 41188
rect 21876 41148 21882 41160
rect 22373 41157 22385 41160
rect 22419 41157 22431 41191
rect 22373 41151 22431 41157
rect 23201 41191 23259 41197
rect 23201 41157 23213 41191
rect 23247 41188 23259 41191
rect 23474 41188 23480 41200
rect 23247 41160 23480 41188
rect 23247 41157 23259 41160
rect 23201 41151 23259 41157
rect 23474 41148 23480 41160
rect 23532 41148 23538 41200
rect 24118 41188 24124 41200
rect 23676 41160 24124 41188
rect 20346 41120 20352 41132
rect 20036 41092 20208 41120
rect 20307 41092 20352 41120
rect 20036 41080 20042 41092
rect 20346 41080 20352 41092
rect 20404 41080 20410 41132
rect 22094 41080 22100 41132
rect 22152 41120 22158 41132
rect 22557 41123 22615 41129
rect 22557 41120 22569 41123
rect 22152 41092 22569 41120
rect 22152 41080 22158 41092
rect 22557 41089 22569 41092
rect 22603 41120 22615 41123
rect 22830 41120 22836 41132
rect 22603 41092 22836 41120
rect 22603 41089 22615 41092
rect 22557 41083 22615 41089
rect 22830 41080 22836 41092
rect 22888 41080 22894 41132
rect 22922 41080 22928 41132
rect 22980 41120 22986 41132
rect 23676 41129 23704 41160
rect 24118 41148 24124 41160
rect 24176 41148 24182 41200
rect 25774 41148 25780 41200
rect 25832 41188 25838 41200
rect 27709 41191 27767 41197
rect 27709 41188 27721 41191
rect 25832 41160 27721 41188
rect 25832 41148 25838 41160
rect 27709 41157 27721 41160
rect 27755 41157 27767 41191
rect 33888 41188 33916 41219
rect 35222 41191 35280 41197
rect 35222 41188 35234 41191
rect 33888 41160 35234 41188
rect 27709 41151 27767 41157
rect 35222 41157 35234 41160
rect 35268 41157 35280 41191
rect 46014 41188 46020 41200
rect 35222 41151 35280 41157
rect 45388 41160 46020 41188
rect 23385 41123 23443 41129
rect 22980 41092 23336 41120
rect 22980 41080 22986 41092
rect 23308 41052 23336 41092
rect 23385 41089 23397 41123
rect 23431 41120 23443 41123
rect 23661 41123 23719 41129
rect 23431 41092 23612 41120
rect 23431 41089 23443 41092
rect 23385 41083 23443 41089
rect 23584 41052 23612 41092
rect 23661 41089 23673 41123
rect 23707 41089 23719 41123
rect 24302 41120 24308 41132
rect 24263 41092 24308 41120
rect 23661 41083 23719 41089
rect 24302 41080 24308 41092
rect 24360 41080 24366 41132
rect 24397 41123 24455 41129
rect 24397 41089 24409 41123
rect 24443 41120 24455 41123
rect 24762 41120 24768 41132
rect 24443 41092 24768 41120
rect 24443 41089 24455 41092
rect 24397 41083 24455 41089
rect 23750 41052 23756 41064
rect 19300 41024 22094 41052
rect 23308 41024 23428 41052
rect 23584 41024 23756 41052
rect 19300 41012 19306 41024
rect 22066 40984 22094 41024
rect 23400 40984 23428 41024
rect 23750 41012 23756 41024
rect 23808 41052 23814 41064
rect 24412 41052 24440 41083
rect 24762 41080 24768 41092
rect 24820 41080 24826 41132
rect 26970 41080 26976 41132
rect 27028 41120 27034 41132
rect 27433 41123 27491 41129
rect 27433 41120 27445 41123
rect 27028 41092 27445 41120
rect 27028 41080 27034 41092
rect 27433 41089 27445 41092
rect 27479 41089 27491 41123
rect 27433 41083 27491 41089
rect 29365 41123 29423 41129
rect 29365 41089 29377 41123
rect 29411 41120 29423 41123
rect 30926 41120 30932 41132
rect 29411 41092 30932 41120
rect 29411 41089 29423 41092
rect 29365 41083 29423 41089
rect 30926 41080 30932 41092
rect 30984 41080 30990 41132
rect 33229 41123 33287 41129
rect 33229 41089 33241 41123
rect 33275 41089 33287 41123
rect 33229 41083 33287 41089
rect 23808 41024 24440 41052
rect 23808 41012 23814 41024
rect 26786 41012 26792 41064
rect 26844 41052 26850 41064
rect 27341 41055 27399 41061
rect 27341 41052 27353 41055
rect 26844 41024 27353 41052
rect 26844 41012 26850 41024
rect 27341 41021 27353 41024
rect 27387 41021 27399 41055
rect 27341 41015 27399 41021
rect 27801 41055 27859 41061
rect 27801 41021 27813 41055
rect 27847 41052 27859 41055
rect 28442 41052 28448 41064
rect 27847 41024 28448 41052
rect 27847 41021 27859 41024
rect 27801 41015 27859 41021
rect 24213 40987 24271 40993
rect 24213 40984 24225 40987
rect 22066 40956 23152 40984
rect 23400 40956 24225 40984
rect 16114 40876 16120 40928
rect 16172 40916 16178 40928
rect 16301 40919 16359 40925
rect 16301 40916 16313 40919
rect 16172 40888 16313 40916
rect 16172 40876 16178 40888
rect 16301 40885 16313 40888
rect 16347 40885 16359 40919
rect 16301 40879 16359 40885
rect 19797 40919 19855 40925
rect 19797 40885 19809 40919
rect 19843 40916 19855 40919
rect 20070 40916 20076 40928
rect 19843 40888 20076 40916
rect 19843 40885 19855 40888
rect 19797 40879 19855 40885
rect 20070 40876 20076 40888
rect 20128 40876 20134 40928
rect 20438 40916 20444 40928
rect 20399 40888 20444 40916
rect 20438 40876 20444 40888
rect 20496 40876 20502 40928
rect 22738 40916 22744 40928
rect 22699 40888 22744 40916
rect 22738 40876 22744 40888
rect 22796 40876 22802 40928
rect 23124 40916 23152 40956
rect 24213 40953 24225 40956
rect 24259 40953 24271 40987
rect 24213 40947 24271 40953
rect 25682 40944 25688 40996
rect 25740 40984 25746 40996
rect 25958 40984 25964 40996
rect 25740 40956 25964 40984
rect 25740 40944 25746 40956
rect 25958 40944 25964 40956
rect 26016 40984 26022 40996
rect 27816 40984 27844 41015
rect 28442 41012 28448 41024
rect 28500 41012 28506 41064
rect 33042 41052 33048 41064
rect 33003 41024 33048 41052
rect 33042 41012 33048 41024
rect 33100 41012 33106 41064
rect 26016 40956 27844 40984
rect 33244 40984 33272 41083
rect 33870 41080 33876 41132
rect 33928 41120 33934 41132
rect 34149 41123 34207 41129
rect 34149 41120 34161 41123
rect 33928 41092 34161 41120
rect 33928 41080 33934 41092
rect 34149 41089 34161 41092
rect 34195 41089 34207 41123
rect 34606 41120 34612 41132
rect 34149 41083 34207 41089
rect 34440 41092 34612 41120
rect 33413 41055 33471 41061
rect 33413 41021 33425 41055
rect 33459 41052 33471 41055
rect 34054 41052 34060 41064
rect 33459 41024 34060 41052
rect 33459 41021 33471 41024
rect 33413 41015 33471 41021
rect 34054 41012 34060 41024
rect 34112 41012 34118 41064
rect 34440 41061 34468 41092
rect 34606 41080 34612 41092
rect 34664 41080 34670 41132
rect 45388 41129 45416 41160
rect 46014 41148 46020 41160
rect 46072 41148 46078 41200
rect 45373 41123 45431 41129
rect 45373 41089 45385 41123
rect 45419 41089 45431 41123
rect 45373 41083 45431 41089
rect 34425 41055 34483 41061
rect 34425 41021 34437 41055
rect 34471 41021 34483 41055
rect 34425 41015 34483 41021
rect 34146 40984 34152 40996
rect 33244 40956 34152 40984
rect 26016 40944 26022 40956
rect 34146 40944 34152 40956
rect 34204 40944 34210 40996
rect 24670 40916 24676 40928
rect 23124 40888 24676 40916
rect 24670 40876 24676 40888
rect 24728 40876 24734 40928
rect 29454 40916 29460 40928
rect 29415 40888 29460 40916
rect 29454 40876 29460 40888
rect 29512 40876 29518 40928
rect 30190 40876 30196 40928
rect 30248 40916 30254 40928
rect 34330 40916 34336 40928
rect 30248 40888 34336 40916
rect 30248 40876 30254 40888
rect 34330 40876 34336 40888
rect 34388 40916 34394 40928
rect 34440 40916 34468 41015
rect 34514 41012 34520 41064
rect 34572 41052 34578 41064
rect 34572 41024 34665 41052
rect 34572 41012 34578 41024
rect 34790 41012 34796 41064
rect 34848 41052 34854 41064
rect 34977 41055 35035 41061
rect 34977 41052 34989 41055
rect 34848 41024 34989 41052
rect 34848 41012 34854 41024
rect 34977 41021 34989 41024
rect 35023 41021 35035 41055
rect 34977 41015 35035 41021
rect 45557 41055 45615 41061
rect 45557 41021 45569 41055
rect 45603 41052 45615 41055
rect 45922 41052 45928 41064
rect 45603 41024 45928 41052
rect 45603 41021 45615 41024
rect 45557 41015 45615 41021
rect 45922 41012 45928 41024
rect 45980 41012 45986 41064
rect 46934 41052 46940 41064
rect 46895 41024 46940 41052
rect 46934 41012 46940 41024
rect 46992 41012 46998 41064
rect 34388 40888 34468 40916
rect 34532 40916 34560 41012
rect 36357 40919 36415 40925
rect 36357 40916 36369 40919
rect 34532 40888 36369 40916
rect 34388 40876 34394 40888
rect 36357 40885 36369 40888
rect 36403 40885 36415 40919
rect 36357 40879 36415 40885
rect 46474 40876 46480 40928
rect 46532 40916 46538 40928
rect 47949 40919 48007 40925
rect 47949 40916 47961 40919
rect 46532 40888 47961 40916
rect 46532 40876 46538 40888
rect 47949 40885 47961 40888
rect 47995 40885 48007 40919
rect 47949 40879 48007 40885
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 2314 40712 2320 40724
rect 2275 40684 2320 40712
rect 2314 40672 2320 40684
rect 2372 40672 2378 40724
rect 15930 40712 15936 40724
rect 15891 40684 15936 40712
rect 15930 40672 15936 40684
rect 15988 40672 15994 40724
rect 16022 40672 16028 40724
rect 16080 40712 16086 40724
rect 17221 40715 17279 40721
rect 17221 40712 17233 40715
rect 16080 40684 17233 40712
rect 16080 40672 16086 40684
rect 17221 40681 17233 40684
rect 17267 40681 17279 40715
rect 17221 40675 17279 40681
rect 21818 40672 21824 40724
rect 21876 40712 21882 40724
rect 22005 40715 22063 40721
rect 22005 40712 22017 40715
rect 21876 40684 22017 40712
rect 21876 40672 21882 40684
rect 22005 40681 22017 40684
rect 22051 40681 22063 40715
rect 22005 40675 22063 40681
rect 22922 40672 22928 40724
rect 22980 40672 22986 40724
rect 23014 40672 23020 40724
rect 23072 40712 23078 40724
rect 23198 40712 23204 40724
rect 23072 40684 23204 40712
rect 23072 40672 23078 40684
rect 23198 40672 23204 40684
rect 23256 40672 23262 40724
rect 23661 40715 23719 40721
rect 23661 40681 23673 40715
rect 23707 40712 23719 40715
rect 23750 40712 23756 40724
rect 23707 40684 23756 40712
rect 23707 40681 23719 40684
rect 23661 40675 23719 40681
rect 23750 40672 23756 40684
rect 23808 40672 23814 40724
rect 30282 40712 30288 40724
rect 23860 40684 30288 40712
rect 22940 40644 22968 40672
rect 22664 40616 22968 40644
rect 16942 40536 16948 40588
rect 17000 40576 17006 40588
rect 17037 40579 17095 40585
rect 17037 40576 17049 40579
rect 17000 40548 17049 40576
rect 17000 40536 17006 40548
rect 17037 40545 17049 40548
rect 17083 40545 17095 40579
rect 17310 40576 17316 40588
rect 17037 40539 17095 40545
rect 17144 40548 17316 40576
rect 2225 40511 2283 40517
rect 2225 40477 2237 40511
rect 2271 40508 2283 40511
rect 2590 40508 2596 40520
rect 2271 40480 2596 40508
rect 2271 40477 2283 40480
rect 2225 40471 2283 40477
rect 2590 40468 2596 40480
rect 2648 40468 2654 40520
rect 16114 40508 16120 40520
rect 16075 40480 16120 40508
rect 16114 40468 16120 40480
rect 16172 40468 16178 40520
rect 16853 40511 16911 40517
rect 16853 40477 16865 40511
rect 16899 40508 16911 40511
rect 17144 40508 17172 40548
rect 17310 40536 17316 40548
rect 17368 40536 17374 40588
rect 20070 40576 20076 40588
rect 20031 40548 20076 40576
rect 20070 40536 20076 40548
rect 20128 40536 20134 40588
rect 16899 40480 17172 40508
rect 17221 40511 17279 40517
rect 16899 40477 16911 40480
rect 16853 40471 16911 40477
rect 17221 40477 17233 40511
rect 17267 40477 17279 40511
rect 17221 40471 17279 40477
rect 16945 40443 17003 40449
rect 16945 40409 16957 40443
rect 16991 40440 17003 40443
rect 17034 40440 17040 40452
rect 16991 40412 17040 40440
rect 16991 40409 17003 40412
rect 16945 40403 17003 40409
rect 17034 40400 17040 40412
rect 17092 40400 17098 40452
rect 17236 40440 17264 40471
rect 19426 40468 19432 40520
rect 19484 40508 19490 40520
rect 19554 40511 19612 40517
rect 19554 40508 19566 40511
rect 19484 40480 19566 40508
rect 19484 40468 19490 40480
rect 19554 40477 19566 40480
rect 19600 40477 19612 40511
rect 19554 40471 19612 40477
rect 19981 40511 20039 40517
rect 19981 40477 19993 40511
rect 20027 40508 20039 40511
rect 20438 40508 20444 40520
rect 20027 40480 20444 40508
rect 20027 40477 20039 40480
rect 19981 40471 20039 40477
rect 20438 40468 20444 40480
rect 20496 40468 20502 40520
rect 20622 40508 20628 40520
rect 20583 40480 20628 40508
rect 20622 40468 20628 40480
rect 20680 40468 20686 40520
rect 22664 40517 22692 40616
rect 23106 40604 23112 40656
rect 23164 40644 23170 40656
rect 23860 40644 23888 40684
rect 30282 40672 30288 40684
rect 30340 40672 30346 40724
rect 33870 40712 33876 40724
rect 33831 40684 33876 40712
rect 33870 40672 33876 40684
rect 33928 40672 33934 40724
rect 45922 40712 45928 40724
rect 45883 40684 45928 40712
rect 45922 40672 45928 40684
rect 45980 40672 45986 40724
rect 23164 40616 23888 40644
rect 23164 40604 23170 40616
rect 30466 40604 30472 40656
rect 30524 40644 30530 40656
rect 30929 40647 30987 40653
rect 30929 40644 30941 40647
rect 30524 40616 30941 40644
rect 30524 40604 30530 40616
rect 30929 40613 30941 40616
rect 30975 40613 30987 40647
rect 30929 40607 30987 40613
rect 33781 40647 33839 40653
rect 33781 40613 33793 40647
rect 33827 40644 33839 40647
rect 34146 40644 34152 40656
rect 33827 40616 34152 40644
rect 33827 40613 33839 40616
rect 33781 40607 33839 40613
rect 34146 40604 34152 40616
rect 34204 40604 34210 40656
rect 22738 40536 22744 40588
rect 22796 40576 22802 40588
rect 25774 40576 25780 40588
rect 22796 40548 23796 40576
rect 25735 40548 25780 40576
rect 22796 40536 22802 40548
rect 22649 40511 22707 40517
rect 22649 40477 22661 40511
rect 22695 40477 22707 40511
rect 22649 40471 22707 40477
rect 22922 40468 22928 40520
rect 22980 40517 22986 40520
rect 22980 40511 23009 40517
rect 22997 40477 23009 40511
rect 23106 40508 23112 40520
rect 23067 40480 23112 40508
rect 22980 40471 23009 40477
rect 22980 40468 22986 40471
rect 23106 40468 23112 40480
rect 23164 40468 23170 40520
rect 23569 40511 23627 40517
rect 23569 40477 23581 40511
rect 23615 40508 23627 40511
rect 23658 40508 23664 40520
rect 23615 40480 23664 40508
rect 23615 40477 23627 40480
rect 23569 40471 23627 40477
rect 23658 40468 23664 40480
rect 23716 40468 23722 40520
rect 23768 40517 23796 40548
rect 25774 40536 25780 40548
rect 25832 40536 25838 40588
rect 26970 40576 26976 40588
rect 26528 40548 26976 40576
rect 26528 40520 26556 40548
rect 26970 40536 26976 40548
rect 27028 40536 27034 40588
rect 32858 40576 32864 40588
rect 31726 40548 32864 40576
rect 23753 40511 23811 40517
rect 23753 40477 23765 40511
rect 23799 40477 23811 40511
rect 24670 40508 24676 40520
rect 24631 40480 24676 40508
rect 23753 40471 23811 40477
rect 24670 40468 24676 40480
rect 24728 40468 24734 40520
rect 25682 40508 25688 40520
rect 25643 40480 25688 40508
rect 25682 40468 25688 40480
rect 25740 40468 25746 40520
rect 26510 40508 26516 40520
rect 26471 40480 26516 40508
rect 26510 40468 26516 40480
rect 26568 40468 26574 40520
rect 26697 40511 26755 40517
rect 26697 40477 26709 40511
rect 26743 40508 26755 40511
rect 26786 40508 26792 40520
rect 26743 40480 26792 40508
rect 26743 40477 26755 40480
rect 26697 40471 26755 40477
rect 26786 40468 26792 40480
rect 26844 40468 26850 40520
rect 27062 40468 27068 40520
rect 27120 40508 27126 40520
rect 27157 40511 27215 40517
rect 27157 40508 27169 40511
rect 27120 40480 27169 40508
rect 27120 40468 27126 40480
rect 27157 40477 27169 40480
rect 27203 40508 27215 40511
rect 30926 40508 30932 40520
rect 27203 40480 27568 40508
rect 30887 40480 30932 40508
rect 27203 40477 27215 40480
rect 27157 40471 27215 40477
rect 27540 40452 27568 40480
rect 30926 40468 30932 40480
rect 30984 40468 30990 40520
rect 31205 40511 31263 40517
rect 31205 40477 31217 40511
rect 31251 40508 31263 40511
rect 31726 40508 31754 40548
rect 32858 40536 32864 40548
rect 32916 40536 32922 40588
rect 33965 40579 34023 40585
rect 33965 40545 33977 40579
rect 34011 40576 34023 40579
rect 34422 40576 34428 40588
rect 34011 40548 34428 40576
rect 34011 40545 34023 40548
rect 33965 40539 34023 40545
rect 34422 40536 34428 40548
rect 34480 40536 34486 40588
rect 46474 40576 46480 40588
rect 46435 40548 46480 40576
rect 46474 40536 46480 40548
rect 46532 40536 46538 40588
rect 31251 40480 31754 40508
rect 32217 40511 32275 40517
rect 31251 40477 31263 40480
rect 31205 40471 31263 40477
rect 32217 40477 32229 40511
rect 32263 40508 32275 40511
rect 32766 40508 32772 40520
rect 32263 40480 32772 40508
rect 32263 40477 32275 40480
rect 32217 40471 32275 40477
rect 32766 40468 32772 40480
rect 32824 40468 32830 40520
rect 33042 40468 33048 40520
rect 33100 40508 33106 40520
rect 33689 40511 33747 40517
rect 33689 40508 33701 40511
rect 33100 40480 33701 40508
rect 33100 40468 33106 40480
rect 33689 40477 33701 40480
rect 33735 40477 33747 40511
rect 33689 40471 33747 40477
rect 45833 40511 45891 40517
rect 45833 40477 45845 40511
rect 45879 40508 45891 40511
rect 45879 40480 46520 40508
rect 45879 40477 45891 40480
rect 45833 40471 45891 40477
rect 20530 40440 20536 40452
rect 17236 40412 20536 40440
rect 20530 40400 20536 40412
rect 20588 40400 20594 40452
rect 20892 40443 20950 40449
rect 20892 40409 20904 40443
rect 20938 40440 20950 40443
rect 22465 40443 22523 40449
rect 22465 40440 22477 40443
rect 20938 40412 22477 40440
rect 20938 40409 20950 40412
rect 20892 40403 20950 40409
rect 22465 40409 22477 40412
rect 22511 40409 22523 40443
rect 22465 40403 22523 40409
rect 22741 40443 22799 40449
rect 22741 40409 22753 40443
rect 22787 40409 22799 40443
rect 22741 40403 22799 40409
rect 22833 40443 22891 40449
rect 22833 40409 22845 40443
rect 22879 40440 22891 40443
rect 23198 40440 23204 40452
rect 22879 40412 23204 40440
rect 22879 40409 22891 40412
rect 22833 40403 22891 40409
rect 19426 40372 19432 40384
rect 19387 40344 19432 40372
rect 19426 40332 19432 40344
rect 19484 40332 19490 40384
rect 19613 40375 19671 40381
rect 19613 40341 19625 40375
rect 19659 40372 19671 40375
rect 19978 40372 19984 40384
rect 19659 40344 19984 40372
rect 19659 40341 19671 40344
rect 19613 40335 19671 40341
rect 19978 40332 19984 40344
rect 20036 40332 20042 40384
rect 22756 40372 22784 40403
rect 23198 40400 23204 40412
rect 23256 40440 23262 40452
rect 25041 40443 25099 40449
rect 25041 40440 25053 40443
rect 23256 40412 25053 40440
rect 23256 40400 23262 40412
rect 25041 40409 25053 40412
rect 25087 40440 25099 40443
rect 26878 40440 26884 40452
rect 25087 40412 26884 40440
rect 25087 40409 25099 40412
rect 25041 40403 25099 40409
rect 26878 40400 26884 40412
rect 26936 40400 26942 40452
rect 27424 40443 27482 40449
rect 27424 40409 27436 40443
rect 27470 40409 27482 40443
rect 27424 40403 27482 40409
rect 23474 40372 23480 40384
rect 22756 40344 23480 40372
rect 23474 40332 23480 40344
rect 23532 40332 23538 40384
rect 26053 40375 26111 40381
rect 26053 40341 26065 40375
rect 26099 40372 26111 40375
rect 26510 40372 26516 40384
rect 26099 40344 26516 40372
rect 26099 40341 26111 40344
rect 26053 40335 26111 40341
rect 26510 40332 26516 40344
rect 26568 40332 26574 40384
rect 26694 40372 26700 40384
rect 26655 40344 26700 40372
rect 26694 40332 26700 40344
rect 26752 40332 26758 40384
rect 27448 40372 27476 40403
rect 27522 40400 27528 40452
rect 27580 40400 27586 40452
rect 28442 40400 28448 40452
rect 28500 40440 28506 40452
rect 34238 40440 34244 40452
rect 28500 40412 34244 40440
rect 28500 40400 28506 40412
rect 34238 40400 34244 40412
rect 34296 40400 34302 40452
rect 27706 40372 27712 40384
rect 27448 40344 27712 40372
rect 27706 40332 27712 40344
rect 27764 40332 27770 40384
rect 28534 40372 28540 40384
rect 28495 40344 28540 40372
rect 28534 40332 28540 40344
rect 28592 40332 28598 40384
rect 31110 40372 31116 40384
rect 31071 40344 31116 40372
rect 31110 40332 31116 40344
rect 31168 40332 31174 40384
rect 32306 40372 32312 40384
rect 32267 40344 32312 40372
rect 32306 40332 32312 40344
rect 32364 40332 32370 40384
rect 46492 40372 46520 40480
rect 46661 40443 46719 40449
rect 46661 40409 46673 40443
rect 46707 40440 46719 40443
rect 47118 40440 47124 40452
rect 46707 40412 47124 40440
rect 46707 40409 46719 40412
rect 46661 40403 46719 40409
rect 47118 40400 47124 40412
rect 47176 40400 47182 40452
rect 48314 40440 48320 40452
rect 48275 40412 48320 40440
rect 48314 40400 48320 40412
rect 48372 40400 48378 40452
rect 47026 40372 47032 40384
rect 46492 40344 47032 40372
rect 47026 40332 47032 40344
rect 47084 40332 47090 40384
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 19797 40171 19855 40177
rect 19797 40137 19809 40171
rect 19843 40168 19855 40171
rect 20346 40168 20352 40180
rect 19843 40140 20352 40168
rect 19843 40137 19855 40140
rect 19797 40131 19855 40137
rect 20346 40128 20352 40140
rect 20404 40128 20410 40180
rect 25774 40128 25780 40180
rect 25832 40168 25838 40180
rect 27706 40168 27712 40180
rect 25832 40140 27476 40168
rect 27667 40140 27712 40168
rect 25832 40128 25838 40140
rect 21818 40060 21824 40112
rect 21876 40100 21882 40112
rect 23106 40100 23112 40112
rect 21876 40072 23112 40100
rect 21876 40060 21882 40072
rect 18684 40035 18742 40041
rect 18684 40001 18696 40035
rect 18730 40032 18742 40035
rect 19426 40032 19432 40044
rect 18730 40004 19432 40032
rect 18730 40001 18742 40004
rect 18684 39995 18742 40001
rect 19426 39992 19432 40004
rect 19484 39992 19490 40044
rect 22572 40041 22600 40072
rect 23106 40060 23112 40072
rect 23164 40060 23170 40112
rect 25682 40100 25688 40112
rect 23400 40072 25688 40100
rect 22557 40035 22615 40041
rect 22557 40001 22569 40035
rect 22603 40001 22615 40035
rect 22557 39995 22615 40001
rect 22741 40035 22799 40041
rect 22741 40001 22753 40035
rect 22787 40032 22799 40035
rect 22830 40032 22836 40044
rect 22787 40004 22836 40032
rect 22787 40001 22799 40004
rect 22741 39995 22799 40001
rect 22830 39992 22836 40004
rect 22888 40032 22894 40044
rect 23400 40032 23428 40072
rect 25682 40060 25688 40072
rect 25740 40060 25746 40112
rect 26694 40060 26700 40112
rect 26752 40100 26758 40112
rect 27448 40109 27476 40140
rect 27706 40128 27712 40140
rect 27764 40128 27770 40180
rect 27798 40128 27804 40180
rect 27856 40168 27862 40180
rect 32585 40171 32643 40177
rect 32585 40168 32597 40171
rect 27856 40140 32597 40168
rect 27856 40128 27862 40140
rect 32585 40137 32597 40140
rect 32631 40137 32643 40171
rect 32585 40131 32643 40137
rect 27341 40103 27399 40109
rect 27341 40100 27353 40103
rect 26752 40072 27353 40100
rect 26752 40060 26758 40072
rect 27341 40069 27353 40072
rect 27387 40069 27399 40103
rect 27341 40063 27399 40069
rect 27433 40103 27491 40109
rect 27433 40069 27445 40103
rect 27479 40100 27491 40103
rect 28534 40100 28540 40112
rect 27479 40072 28540 40100
rect 27479 40069 27491 40072
rect 27433 40063 27491 40069
rect 28534 40060 28540 40072
rect 28592 40060 28598 40112
rect 30466 40100 30472 40112
rect 28644 40072 30328 40100
rect 30427 40072 30472 40100
rect 27154 40032 27160 40044
rect 22888 40004 23428 40032
rect 27115 40004 27160 40032
rect 22888 39992 22894 40004
rect 27154 39992 27160 40004
rect 27212 39992 27218 40044
rect 27522 40032 27528 40044
rect 27483 40004 27528 40032
rect 27522 39992 27528 40004
rect 27580 39992 27586 40044
rect 28261 40035 28319 40041
rect 28261 40001 28273 40035
rect 28307 40032 28319 40035
rect 28644 40032 28672 40072
rect 28307 40004 28672 40032
rect 30300 40032 30328 40072
rect 30466 40060 30472 40072
rect 30524 40060 30530 40112
rect 32306 40060 32312 40112
rect 32364 40060 32370 40112
rect 32401 40103 32459 40109
rect 32401 40069 32413 40103
rect 32447 40100 32459 40103
rect 32858 40100 32864 40112
rect 32447 40072 32864 40100
rect 32447 40069 32459 40072
rect 32401 40063 32459 40069
rect 32858 40060 32864 40072
rect 32916 40060 32922 40112
rect 32308 40057 32366 40060
rect 30653 40035 30711 40041
rect 30300 40004 30604 40032
rect 28307 40001 28319 40004
rect 28261 39995 28319 40001
rect 18414 39964 18420 39976
rect 18375 39936 18420 39964
rect 18414 39924 18420 39936
rect 18472 39924 18478 39976
rect 22649 39967 22707 39973
rect 22649 39933 22661 39967
rect 22695 39964 22707 39967
rect 23658 39964 23664 39976
rect 22695 39936 23664 39964
rect 22695 39933 22707 39936
rect 22649 39927 22707 39933
rect 23658 39924 23664 39936
rect 23716 39924 23722 39976
rect 26234 39924 26240 39976
rect 26292 39964 26298 39976
rect 27540 39964 27568 39992
rect 30190 39964 30196 39976
rect 26292 39936 30196 39964
rect 26292 39924 26298 39936
rect 30190 39924 30196 39936
rect 30248 39924 30254 39976
rect 30576 39964 30604 40004
rect 30653 40001 30665 40035
rect 30699 40032 30711 40035
rect 30926 40032 30932 40044
rect 30699 40004 30932 40032
rect 30699 40001 30711 40004
rect 30653 39995 30711 40001
rect 30926 39992 30932 40004
rect 30984 39992 30990 40044
rect 32308 40023 32320 40057
rect 32354 40023 32366 40057
rect 32674 40032 32680 40044
rect 32308 40017 32366 40023
rect 32635 40004 32680 40032
rect 32674 39992 32680 40004
rect 32732 39992 32738 40044
rect 47026 40032 47032 40044
rect 46939 40004 47032 40032
rect 47026 39992 47032 40004
rect 47084 39992 47090 40044
rect 47118 39992 47124 40044
rect 47176 40032 47182 40044
rect 47176 40004 47221 40032
rect 47176 39992 47182 40004
rect 30742 39964 30748 39976
rect 30576 39936 30748 39964
rect 30742 39924 30748 39936
rect 30800 39964 30806 39976
rect 31018 39964 31024 39976
rect 30800 39936 31024 39964
rect 30800 39924 30806 39936
rect 31018 39924 31024 39936
rect 31076 39924 31082 39976
rect 32493 39967 32551 39973
rect 32493 39933 32505 39967
rect 32539 39964 32551 39967
rect 33042 39964 33048 39976
rect 32539 39936 33048 39964
rect 32539 39933 32551 39936
rect 32493 39927 32551 39933
rect 25590 39856 25596 39908
rect 25648 39896 25654 39908
rect 31110 39896 31116 39908
rect 25648 39868 31116 39896
rect 25648 39856 25654 39868
rect 31110 39856 31116 39868
rect 31168 39896 31174 39908
rect 32508 39896 32536 39927
rect 33042 39924 33048 39936
rect 33100 39924 33106 39976
rect 47044 39964 47072 39992
rect 47486 39964 47492 39976
rect 47044 39936 47492 39964
rect 47486 39924 47492 39936
rect 47544 39924 47550 39976
rect 31168 39868 32536 39896
rect 31168 39856 31174 39868
rect 28353 39831 28411 39837
rect 28353 39797 28365 39831
rect 28399 39828 28411 39831
rect 28442 39828 28448 39840
rect 28399 39800 28448 39828
rect 28399 39797 28411 39800
rect 28353 39791 28411 39797
rect 28442 39788 28448 39800
rect 28500 39788 28506 39840
rect 30374 39788 30380 39840
rect 30432 39828 30438 39840
rect 30837 39831 30895 39837
rect 30837 39828 30849 39831
rect 30432 39800 30849 39828
rect 30432 39788 30438 39800
rect 30837 39797 30849 39800
rect 30883 39797 30895 39831
rect 30837 39791 30895 39797
rect 46474 39788 46480 39840
rect 46532 39828 46538 39840
rect 47949 39831 48007 39837
rect 47949 39828 47961 39831
rect 46532 39800 47961 39828
rect 46532 39788 46538 39800
rect 47949 39797 47961 39800
rect 47995 39797 48007 39831
rect 47949 39791 48007 39797
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 26697 39627 26755 39633
rect 26697 39593 26709 39627
rect 26743 39624 26755 39627
rect 27154 39624 27160 39636
rect 26743 39596 27160 39624
rect 26743 39593 26755 39596
rect 26697 39587 26755 39593
rect 27154 39584 27160 39596
rect 27212 39584 27218 39636
rect 30466 39584 30472 39636
rect 30524 39624 30530 39636
rect 30837 39627 30895 39633
rect 30837 39624 30849 39627
rect 30524 39596 30849 39624
rect 30524 39584 30530 39596
rect 30837 39593 30849 39596
rect 30883 39593 30895 39627
rect 32033 39627 32091 39633
rect 32033 39624 32045 39627
rect 30837 39587 30895 39593
rect 31404 39596 32045 39624
rect 26510 39516 26516 39568
rect 26568 39556 26574 39568
rect 27065 39559 27123 39565
rect 27065 39556 27077 39559
rect 26568 39528 27077 39556
rect 26568 39516 26574 39528
rect 27065 39525 27077 39528
rect 27111 39525 27123 39559
rect 27985 39559 28043 39565
rect 27985 39556 27997 39559
rect 27065 39519 27123 39525
rect 27172 39528 27997 39556
rect 14090 39448 14096 39500
rect 14148 39488 14154 39500
rect 14274 39488 14280 39500
rect 14148 39460 14280 39488
rect 14148 39448 14154 39460
rect 14274 39448 14280 39460
rect 14332 39448 14338 39500
rect 18414 39448 18420 39500
rect 18472 39488 18478 39500
rect 20165 39491 20223 39497
rect 20165 39488 20177 39491
rect 18472 39460 20177 39488
rect 18472 39448 18478 39460
rect 20165 39457 20177 39460
rect 20211 39488 20223 39491
rect 20622 39488 20628 39500
rect 20211 39460 20628 39488
rect 20211 39457 20223 39460
rect 20165 39451 20223 39457
rect 20622 39448 20628 39460
rect 20680 39448 20686 39500
rect 26786 39448 26792 39500
rect 26844 39488 26850 39500
rect 27172 39497 27200 39528
rect 27985 39525 27997 39528
rect 28031 39525 28043 39559
rect 27985 39519 28043 39525
rect 27157 39491 27215 39497
rect 27157 39488 27169 39491
rect 26844 39460 27169 39488
rect 26844 39448 26850 39460
rect 27157 39457 27169 39460
rect 27203 39457 27215 39491
rect 27157 39451 27215 39457
rect 27617 39491 27675 39497
rect 27617 39457 27629 39491
rect 27663 39488 27675 39491
rect 29454 39488 29460 39500
rect 27663 39460 29460 39488
rect 27663 39457 27675 39460
rect 27617 39451 27675 39457
rect 29454 39448 29460 39460
rect 29512 39448 29518 39500
rect 29917 39491 29975 39497
rect 29917 39457 29929 39491
rect 29963 39488 29975 39491
rect 30852 39488 30880 39587
rect 31404 39488 31432 39596
rect 32033 39593 32045 39596
rect 32079 39593 32091 39627
rect 32033 39587 32091 39593
rect 33597 39559 33655 39565
rect 33597 39556 33609 39559
rect 29963 39460 30696 39488
rect 30852 39460 31432 39488
rect 29963 39457 29975 39460
rect 29917 39451 29975 39457
rect 30668 39432 30696 39460
rect 26878 39420 26884 39432
rect 26791 39392 26884 39420
rect 26878 39380 26884 39392
rect 26936 39420 26942 39432
rect 27798 39420 27804 39432
rect 26936 39392 27476 39420
rect 27759 39392 27804 39420
rect 26936 39380 26942 39392
rect 13906 39312 13912 39364
rect 13964 39352 13970 39364
rect 14522 39355 14580 39361
rect 14522 39352 14534 39355
rect 13964 39324 14534 39352
rect 13964 39312 13970 39324
rect 14522 39321 14534 39324
rect 14568 39321 14580 39355
rect 19426 39352 19432 39364
rect 19387 39324 19432 39352
rect 14522 39315 14580 39321
rect 19426 39312 19432 39324
rect 19484 39312 19490 39364
rect 15194 39244 15200 39296
rect 15252 39284 15258 39296
rect 15657 39287 15715 39293
rect 15657 39284 15669 39287
rect 15252 39256 15669 39284
rect 15252 39244 15258 39256
rect 15657 39253 15669 39256
rect 15703 39253 15715 39287
rect 27448 39284 27476 39392
rect 27798 39380 27804 39392
rect 27856 39380 27862 39432
rect 29825 39423 29883 39429
rect 29825 39389 29837 39423
rect 29871 39389 29883 39423
rect 29825 39383 29883 39389
rect 30009 39423 30067 39429
rect 30009 39389 30021 39423
rect 30055 39420 30067 39423
rect 30466 39420 30472 39432
rect 30055 39392 30472 39420
rect 30055 39389 30067 39392
rect 30009 39383 30067 39389
rect 29840 39352 29868 39383
rect 30466 39380 30472 39392
rect 30524 39380 30530 39432
rect 30650 39420 30656 39432
rect 30563 39392 30656 39420
rect 30650 39380 30656 39392
rect 30708 39380 30714 39432
rect 30926 39420 30932 39432
rect 30839 39392 30932 39420
rect 30926 39380 30932 39392
rect 30984 39380 30990 39432
rect 31404 39429 31432 39460
rect 32048 39528 33609 39556
rect 32048 39432 32076 39528
rect 33597 39525 33609 39528
rect 33643 39556 33655 39559
rect 34054 39556 34060 39568
rect 33643 39528 34060 39556
rect 33643 39525 33655 39528
rect 33597 39519 33655 39525
rect 34054 39516 34060 39528
rect 34112 39516 34118 39568
rect 33321 39491 33379 39497
rect 33321 39457 33333 39491
rect 33367 39488 33379 39491
rect 34146 39488 34152 39500
rect 33367 39460 34152 39488
rect 33367 39457 33379 39460
rect 33321 39451 33379 39457
rect 34146 39448 34152 39460
rect 34204 39448 34210 39500
rect 46474 39488 46480 39500
rect 46435 39460 46480 39488
rect 46474 39448 46480 39460
rect 46532 39448 46538 39500
rect 48222 39488 48228 39500
rect 48183 39460 48228 39488
rect 48222 39448 48228 39460
rect 48280 39448 48286 39500
rect 31389 39423 31447 39429
rect 31389 39389 31401 39423
rect 31435 39389 31447 39423
rect 31389 39383 31447 39389
rect 31573 39423 31631 39429
rect 31573 39389 31585 39423
rect 31619 39420 31631 39423
rect 32030 39420 32036 39432
rect 31619 39392 31708 39420
rect 31991 39392 32036 39420
rect 31619 39389 31631 39392
rect 31573 39383 31631 39389
rect 30558 39352 30564 39364
rect 29840 39324 30564 39352
rect 30558 39312 30564 39324
rect 30616 39312 30622 39364
rect 30944 39352 30972 39380
rect 31680 39364 31708 39392
rect 32030 39380 32036 39392
rect 32088 39380 32094 39432
rect 32125 39423 32183 39429
rect 32125 39389 32137 39423
rect 32171 39389 32183 39423
rect 32125 39383 32183 39389
rect 33229 39423 33287 39429
rect 33229 39389 33241 39423
rect 33275 39389 33287 39423
rect 33229 39383 33287 39389
rect 31662 39352 31668 39364
rect 30944 39324 31668 39352
rect 31662 39312 31668 39324
rect 31720 39352 31726 39364
rect 32140 39352 32168 39383
rect 33244 39352 33272 39383
rect 31720 39324 32168 39352
rect 32324 39324 33272 39352
rect 46661 39355 46719 39361
rect 31720 39312 31726 39324
rect 30098 39284 30104 39296
rect 27448 39256 30104 39284
rect 15657 39247 15715 39253
rect 30098 39244 30104 39256
rect 30156 39244 30162 39296
rect 30466 39284 30472 39296
rect 30427 39256 30472 39284
rect 30466 39244 30472 39256
rect 30524 39244 30530 39296
rect 31478 39284 31484 39296
rect 31439 39256 31484 39284
rect 31478 39244 31484 39256
rect 31536 39244 31542 39296
rect 31570 39244 31576 39296
rect 31628 39284 31634 39296
rect 32324 39284 32352 39324
rect 46661 39321 46673 39355
rect 46707 39352 46719 39355
rect 47854 39352 47860 39364
rect 46707 39324 47860 39352
rect 46707 39321 46719 39324
rect 46661 39315 46719 39321
rect 47854 39312 47860 39324
rect 47912 39312 47918 39364
rect 31628 39256 32352 39284
rect 31628 39244 31634 39256
rect 32398 39244 32404 39296
rect 32456 39284 32462 39296
rect 32456 39256 32501 39284
rect 32456 39244 32462 39256
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 13906 39080 13912 39092
rect 13867 39052 13912 39080
rect 13906 39040 13912 39052
rect 13964 39040 13970 39092
rect 19797 39083 19855 39089
rect 19797 39049 19809 39083
rect 19843 39080 19855 39083
rect 19978 39080 19984 39092
rect 19843 39052 19984 39080
rect 19843 39049 19855 39052
rect 19797 39043 19855 39049
rect 19978 39040 19984 39052
rect 20036 39040 20042 39092
rect 20441 39083 20499 39089
rect 20441 39049 20453 39083
rect 20487 39080 20499 39083
rect 21082 39080 21088 39092
rect 20487 39052 21088 39080
rect 20487 39049 20499 39052
rect 20441 39043 20499 39049
rect 21082 39040 21088 39052
rect 21140 39080 21146 39092
rect 22370 39080 22376 39092
rect 21140 39052 22376 39080
rect 21140 39040 21146 39052
rect 22370 39040 22376 39052
rect 22428 39040 22434 39092
rect 30377 39083 30435 39089
rect 30377 39049 30389 39083
rect 30423 39080 30435 39083
rect 30558 39080 30564 39092
rect 30423 39052 30564 39080
rect 30423 39049 30435 39052
rect 30377 39043 30435 39049
rect 30558 39040 30564 39052
rect 30616 39040 30622 39092
rect 31018 39080 31024 39092
rect 30979 39052 31024 39080
rect 31018 39040 31024 39052
rect 31076 39080 31082 39092
rect 32309 39083 32367 39089
rect 31076 39052 32168 39080
rect 31076 39040 31082 39052
rect 18414 39012 18420 39024
rect 14844 38984 18420 39012
rect 1578 38944 1584 38956
rect 1539 38916 1584 38944
rect 1578 38904 1584 38916
rect 1636 38904 1642 38956
rect 14090 38944 14096 38956
rect 14051 38916 14096 38944
rect 14090 38904 14096 38916
rect 14148 38904 14154 38956
rect 14274 38904 14280 38956
rect 14332 38944 14338 38956
rect 14844 38953 14872 38984
rect 14829 38947 14887 38953
rect 14829 38944 14841 38947
rect 14332 38916 14841 38944
rect 14332 38904 14338 38916
rect 14829 38913 14841 38916
rect 14875 38913 14887 38947
rect 14829 38907 14887 38913
rect 15096 38947 15154 38953
rect 15096 38913 15108 38947
rect 15142 38944 15154 38947
rect 15470 38944 15476 38956
rect 15142 38916 15476 38944
rect 15142 38913 15154 38916
rect 15096 38907 15154 38913
rect 15470 38904 15476 38916
rect 15528 38904 15534 38956
rect 17236 38953 17264 38984
rect 18414 38972 18420 38984
rect 18472 38972 18478 39024
rect 25406 39012 25412 39024
rect 19628 38984 25412 39012
rect 19628 38956 19656 38984
rect 25406 38972 25412 38984
rect 25464 38972 25470 39024
rect 17494 38953 17500 38956
rect 17221 38947 17279 38953
rect 17221 38913 17233 38947
rect 17267 38913 17279 38947
rect 17221 38907 17279 38913
rect 17488 38907 17500 38953
rect 17552 38944 17558 38956
rect 19610 38944 19616 38956
rect 17552 38916 17588 38944
rect 19571 38916 19616 38944
rect 17494 38904 17500 38907
rect 17552 38904 17558 38916
rect 19610 38904 19616 38916
rect 19668 38904 19674 38956
rect 19978 38904 19984 38956
rect 20036 38944 20042 38956
rect 20257 38947 20315 38953
rect 20257 38944 20269 38947
rect 20036 38916 20269 38944
rect 20036 38904 20042 38916
rect 20257 38913 20269 38916
rect 20303 38913 20315 38947
rect 20257 38907 20315 38913
rect 20530 38904 20536 38956
rect 20588 38944 20594 38956
rect 22373 38947 22431 38953
rect 20588 38916 22094 38944
rect 20588 38904 20594 38916
rect 14366 38876 14372 38888
rect 14327 38848 14372 38876
rect 14366 38836 14372 38848
rect 14424 38836 14430 38888
rect 19429 38879 19487 38885
rect 19429 38845 19441 38879
rect 19475 38876 19487 38879
rect 20438 38876 20444 38888
rect 19475 38848 20444 38876
rect 19475 38845 19487 38848
rect 19429 38839 19487 38845
rect 20438 38836 20444 38848
rect 20496 38836 20502 38888
rect 22066 38876 22094 38916
rect 22373 38913 22385 38947
rect 22419 38944 22431 38947
rect 22646 38944 22652 38956
rect 22419 38916 22652 38944
rect 22419 38913 22431 38916
rect 22373 38907 22431 38913
rect 22646 38904 22652 38916
rect 22704 38904 22710 38956
rect 24210 38944 24216 38956
rect 24171 38916 24216 38944
rect 24210 38904 24216 38916
rect 24268 38904 24274 38956
rect 24673 38947 24731 38953
rect 24673 38913 24685 38947
rect 24719 38944 24731 38947
rect 25038 38944 25044 38956
rect 24719 38916 25044 38944
rect 24719 38913 24731 38916
rect 24673 38907 24731 38913
rect 25038 38904 25044 38916
rect 25096 38904 25102 38956
rect 25314 38944 25320 38956
rect 25275 38916 25320 38944
rect 25314 38904 25320 38916
rect 25372 38904 25378 38956
rect 26053 38947 26111 38953
rect 26053 38944 26065 38947
rect 25700 38916 26065 38944
rect 22465 38879 22523 38885
rect 22465 38876 22477 38879
rect 22066 38848 22477 38876
rect 22465 38845 22477 38848
rect 22511 38845 22523 38879
rect 22465 38839 22523 38845
rect 23201 38879 23259 38885
rect 23201 38845 23213 38879
rect 23247 38876 23259 38879
rect 23382 38876 23388 38888
rect 23247 38848 23388 38876
rect 23247 38845 23259 38848
rect 23201 38839 23259 38845
rect 23382 38836 23388 38848
rect 23440 38836 23446 38888
rect 24946 38876 24952 38888
rect 24907 38848 24952 38876
rect 24946 38836 24952 38848
rect 25004 38836 25010 38888
rect 25130 38836 25136 38888
rect 25188 38876 25194 38888
rect 25700 38876 25728 38916
rect 26053 38913 26065 38916
rect 26099 38913 26111 38947
rect 26053 38907 26111 38913
rect 29264 38947 29322 38953
rect 29264 38913 29276 38947
rect 29310 38944 29322 38947
rect 29730 38944 29736 38956
rect 29310 38916 29736 38944
rect 29310 38913 29322 38916
rect 29264 38907 29322 38913
rect 29730 38904 29736 38916
rect 29788 38904 29794 38956
rect 30926 38944 30932 38956
rect 30887 38916 30932 38944
rect 30926 38904 30932 38916
rect 30984 38944 30990 38956
rect 31570 38944 31576 38956
rect 30984 38916 31576 38944
rect 30984 38904 30990 38916
rect 31570 38904 31576 38916
rect 31628 38904 31634 38956
rect 32140 38944 32168 39052
rect 32309 39049 32321 39083
rect 32355 39080 32367 39083
rect 32674 39080 32680 39092
rect 32355 39052 32680 39080
rect 32355 39049 32367 39052
rect 32309 39043 32367 39049
rect 32674 39040 32680 39052
rect 32732 39040 32738 39092
rect 33134 39080 33140 39092
rect 32784 39052 33140 39080
rect 32784 38953 32812 39052
rect 33134 39040 33140 39052
rect 33192 39040 33198 39092
rect 47854 39080 47860 39092
rect 47815 39052 47860 39080
rect 47854 39040 47860 39052
rect 47912 39040 47918 39092
rect 32858 38972 32864 39024
rect 32916 39012 32922 39024
rect 32916 38984 33088 39012
rect 32916 38972 32922 38984
rect 33060 38953 33088 38984
rect 34716 38984 45554 39012
rect 32585 38947 32643 38953
rect 32585 38944 32597 38947
rect 32140 38916 32597 38944
rect 32585 38913 32597 38916
rect 32631 38913 32643 38947
rect 32585 38907 32643 38913
rect 32769 38947 32827 38953
rect 32769 38913 32781 38947
rect 32815 38913 32827 38947
rect 32769 38907 32827 38913
rect 33045 38947 33103 38953
rect 33045 38913 33057 38947
rect 33091 38913 33103 38947
rect 34054 38944 34060 38956
rect 34015 38916 34060 38944
rect 33045 38907 33103 38913
rect 34054 38904 34060 38916
rect 34112 38904 34118 38956
rect 26142 38876 26148 38888
rect 25188 38848 25728 38876
rect 26103 38848 26148 38876
rect 25188 38836 25194 38848
rect 26142 38836 26148 38848
rect 26200 38836 26206 38888
rect 27062 38836 27068 38888
rect 27120 38876 27126 38888
rect 28997 38879 29055 38885
rect 28997 38876 29009 38879
rect 27120 38848 29009 38876
rect 27120 38836 27126 38848
rect 28997 38845 29009 38848
rect 29043 38845 29055 38879
rect 28997 38839 29055 38845
rect 30466 38836 30472 38888
rect 30524 38876 30530 38888
rect 33965 38879 34023 38885
rect 33965 38876 33977 38879
rect 30524 38848 33977 38876
rect 30524 38836 30530 38848
rect 33965 38845 33977 38848
rect 34011 38845 34023 38879
rect 33965 38839 34023 38845
rect 23474 38808 23480 38820
rect 23435 38780 23480 38808
rect 23474 38768 23480 38780
rect 23532 38768 23538 38820
rect 25590 38808 25596 38820
rect 25551 38780 25596 38808
rect 25590 38768 25596 38780
rect 25648 38768 25654 38820
rect 26421 38811 26479 38817
rect 26421 38808 26433 38811
rect 25700 38780 26433 38808
rect 1765 38743 1823 38749
rect 1765 38709 1777 38743
rect 1811 38740 1823 38743
rect 1854 38740 1860 38752
rect 1811 38712 1860 38740
rect 1811 38709 1823 38712
rect 1765 38703 1823 38709
rect 1854 38700 1860 38712
rect 1912 38700 1918 38752
rect 14277 38743 14335 38749
rect 14277 38709 14289 38743
rect 14323 38740 14335 38743
rect 15562 38740 15568 38752
rect 14323 38712 15568 38740
rect 14323 38709 14335 38712
rect 14277 38703 14335 38709
rect 15562 38700 15568 38712
rect 15620 38700 15626 38752
rect 16114 38700 16120 38752
rect 16172 38740 16178 38752
rect 16209 38743 16267 38749
rect 16209 38740 16221 38743
rect 16172 38712 16221 38740
rect 16172 38700 16178 38712
rect 16209 38709 16221 38712
rect 16255 38709 16267 38743
rect 16209 38703 16267 38709
rect 18414 38700 18420 38752
rect 18472 38740 18478 38752
rect 18601 38743 18659 38749
rect 18601 38740 18613 38743
rect 18472 38712 18613 38740
rect 18472 38700 18478 38712
rect 18601 38709 18613 38712
rect 18647 38709 18659 38743
rect 22554 38740 22560 38752
rect 22515 38712 22560 38740
rect 18601 38703 18659 38709
rect 22554 38700 22560 38712
rect 22612 38700 22618 38752
rect 22738 38740 22744 38752
rect 22699 38712 22744 38740
rect 22738 38700 22744 38712
rect 22796 38700 22802 38752
rect 23566 38700 23572 38752
rect 23624 38740 23630 38752
rect 23661 38743 23719 38749
rect 23661 38740 23673 38743
rect 23624 38712 23673 38740
rect 23624 38700 23630 38712
rect 23661 38709 23673 38712
rect 23707 38709 23719 38743
rect 23661 38703 23719 38709
rect 24854 38700 24860 38752
rect 24912 38740 24918 38752
rect 25700 38740 25728 38780
rect 26421 38777 26433 38780
rect 26467 38777 26479 38811
rect 34716 38808 34744 38984
rect 35342 38953 35348 38956
rect 35336 38907 35348 38953
rect 35400 38944 35406 38956
rect 45526 38944 45554 38984
rect 47302 38944 47308 38956
rect 35400 38916 35436 38944
rect 45526 38916 47308 38944
rect 35342 38904 35348 38907
rect 35400 38904 35406 38916
rect 47302 38904 47308 38916
rect 47360 38944 47366 38956
rect 47765 38947 47823 38953
rect 47765 38944 47777 38947
rect 47360 38916 47777 38944
rect 47360 38904 47366 38916
rect 47765 38913 47777 38916
rect 47811 38913 47823 38947
rect 47765 38907 47823 38913
rect 34790 38836 34796 38888
rect 34848 38876 34854 38888
rect 35069 38879 35127 38885
rect 35069 38876 35081 38879
rect 34848 38848 35081 38876
rect 34848 38836 34854 38848
rect 35069 38845 35081 38848
rect 35115 38845 35127 38879
rect 35069 38839 35127 38845
rect 26421 38771 26479 38777
rect 29932 38780 34744 38808
rect 26142 38740 26148 38752
rect 24912 38712 25728 38740
rect 26103 38712 26148 38740
rect 24912 38700 24918 38712
rect 26142 38700 26148 38712
rect 26200 38700 26206 38752
rect 29178 38700 29184 38752
rect 29236 38740 29242 38752
rect 29932 38740 29960 38780
rect 32674 38740 32680 38752
rect 29236 38712 29960 38740
rect 32635 38712 32680 38740
rect 29236 38700 29242 38712
rect 32674 38700 32680 38712
rect 32732 38700 32738 38752
rect 32861 38743 32919 38749
rect 32861 38709 32873 38743
rect 32907 38740 32919 38743
rect 34146 38740 34152 38752
rect 32907 38712 34152 38740
rect 32907 38709 32919 38712
rect 32861 38703 32919 38709
rect 34146 38700 34152 38712
rect 34204 38700 34210 38752
rect 34425 38743 34483 38749
rect 34425 38709 34437 38743
rect 34471 38740 34483 38743
rect 34698 38740 34704 38752
rect 34471 38712 34704 38740
rect 34471 38709 34483 38712
rect 34425 38703 34483 38709
rect 34698 38700 34704 38712
rect 34756 38700 34762 38752
rect 35434 38700 35440 38752
rect 35492 38740 35498 38752
rect 36449 38743 36507 38749
rect 36449 38740 36461 38743
rect 35492 38712 36461 38740
rect 35492 38700 35498 38712
rect 36449 38709 36461 38712
rect 36495 38709 36507 38743
rect 36449 38703 36507 38709
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 14090 38496 14096 38548
rect 14148 38536 14154 38548
rect 14369 38539 14427 38545
rect 14369 38536 14381 38539
rect 14148 38508 14381 38536
rect 14148 38496 14154 38508
rect 14369 38505 14381 38508
rect 14415 38505 14427 38539
rect 14369 38499 14427 38505
rect 17126 38496 17132 38548
rect 17184 38536 17190 38548
rect 19610 38536 19616 38548
rect 17184 38508 19616 38536
rect 17184 38496 17190 38508
rect 19610 38496 19616 38508
rect 19668 38496 19674 38548
rect 22833 38539 22891 38545
rect 22833 38505 22845 38539
rect 22879 38536 22891 38539
rect 23106 38536 23112 38548
rect 22879 38508 23112 38536
rect 22879 38505 22891 38508
rect 22833 38499 22891 38505
rect 23106 38496 23112 38508
rect 23164 38536 23170 38548
rect 24210 38536 24216 38548
rect 23164 38508 24216 38536
rect 23164 38496 23170 38508
rect 24210 38496 24216 38508
rect 24268 38496 24274 38548
rect 24854 38536 24860 38548
rect 24815 38508 24860 38536
rect 24854 38496 24860 38508
rect 24912 38496 24918 38548
rect 25038 38536 25044 38548
rect 24999 38508 25044 38536
rect 25038 38496 25044 38508
rect 25096 38496 25102 38548
rect 29730 38536 29736 38548
rect 29691 38508 29736 38536
rect 29730 38496 29736 38508
rect 29788 38496 29794 38548
rect 32030 38496 32036 38548
rect 32088 38536 32094 38548
rect 32309 38539 32367 38545
rect 32309 38536 32321 38539
rect 32088 38508 32321 38536
rect 32088 38496 32094 38508
rect 32309 38505 32321 38508
rect 32355 38505 32367 38539
rect 32766 38536 32772 38548
rect 32727 38508 32772 38536
rect 32309 38499 32367 38505
rect 32766 38496 32772 38508
rect 32824 38496 32830 38548
rect 32858 38496 32864 38548
rect 32916 38496 32922 38548
rect 35342 38496 35348 38548
rect 35400 38536 35406 38548
rect 35437 38539 35495 38545
rect 35437 38536 35449 38539
rect 35400 38508 35449 38536
rect 35400 38496 35406 38508
rect 35437 38505 35449 38508
rect 35483 38505 35495 38539
rect 35437 38499 35495 38505
rect 22554 38428 22560 38480
rect 22612 38468 22618 38480
rect 23017 38471 23075 38477
rect 23017 38468 23029 38471
rect 22612 38440 23029 38468
rect 22612 38428 22618 38440
rect 23017 38437 23029 38440
rect 23063 38437 23075 38471
rect 23017 38431 23075 38437
rect 23842 38428 23848 38480
rect 23900 38428 23906 38480
rect 23934 38428 23940 38480
rect 23992 38428 23998 38480
rect 24872 38468 24900 38496
rect 24044 38440 24900 38468
rect 14568 38372 20208 38400
rect 14568 38341 14596 38372
rect 14553 38335 14611 38341
rect 14553 38301 14565 38335
rect 14599 38301 14611 38335
rect 14553 38295 14611 38301
rect 14829 38335 14887 38341
rect 14829 38301 14841 38335
rect 14875 38301 14887 38335
rect 14829 38295 14887 38301
rect 15013 38335 15071 38341
rect 15013 38301 15025 38335
rect 15059 38332 15071 38335
rect 15194 38332 15200 38344
rect 15059 38304 15200 38332
rect 15059 38301 15071 38304
rect 15013 38295 15071 38301
rect 14844 38264 14872 38295
rect 15194 38292 15200 38304
rect 15252 38292 15258 38344
rect 15672 38341 15700 38372
rect 15657 38335 15715 38341
rect 15657 38301 15669 38335
rect 15703 38301 15715 38335
rect 15657 38295 15715 38301
rect 15933 38335 15991 38341
rect 15933 38301 15945 38335
rect 15979 38301 15991 38335
rect 16114 38332 16120 38344
rect 16075 38304 16120 38332
rect 15933 38295 15991 38301
rect 15948 38264 15976 38295
rect 16114 38292 16120 38304
rect 16172 38292 16178 38344
rect 16850 38332 16856 38344
rect 16811 38304 16856 38332
rect 16850 38292 16856 38304
rect 16908 38292 16914 38344
rect 17972 38341 18000 38372
rect 17957 38335 18015 38341
rect 17957 38301 17969 38335
rect 18003 38301 18015 38335
rect 17957 38295 18015 38301
rect 18233 38335 18291 38341
rect 18233 38301 18245 38335
rect 18279 38301 18291 38335
rect 18414 38332 18420 38344
rect 18375 38304 18420 38332
rect 18233 38295 18291 38301
rect 17126 38264 17132 38276
rect 14844 38236 15976 38264
rect 17087 38236 17132 38264
rect 15378 38156 15384 38208
rect 15436 38196 15442 38208
rect 15473 38199 15531 38205
rect 15473 38196 15485 38199
rect 15436 38168 15485 38196
rect 15436 38156 15442 38168
rect 15473 38165 15485 38168
rect 15519 38165 15531 38199
rect 15948 38196 15976 38236
rect 17126 38224 17132 38236
rect 17184 38224 17190 38276
rect 17586 38224 17592 38276
rect 17644 38264 17650 38276
rect 18248 38264 18276 38295
rect 18414 38292 18420 38304
rect 18472 38292 18478 38344
rect 19978 38264 19984 38276
rect 17644 38236 18276 38264
rect 19939 38236 19984 38264
rect 17644 38224 17650 38236
rect 19978 38224 19984 38236
rect 20036 38224 20042 38276
rect 17604 38196 17632 38224
rect 15948 38168 17632 38196
rect 15473 38159 15531 38165
rect 17678 38156 17684 38208
rect 17736 38196 17742 38208
rect 17773 38199 17831 38205
rect 17773 38196 17785 38199
rect 17736 38168 17785 38196
rect 17736 38156 17742 38168
rect 17773 38165 17785 38168
rect 17819 38165 17831 38199
rect 17773 38159 17831 38165
rect 19242 38156 19248 38208
rect 19300 38196 19306 38208
rect 20073 38199 20131 38205
rect 20073 38196 20085 38199
rect 19300 38168 20085 38196
rect 19300 38156 19306 38168
rect 20073 38165 20085 38168
rect 20119 38165 20131 38199
rect 20180 38196 20208 38372
rect 20622 38360 20628 38412
rect 20680 38400 20686 38412
rect 20809 38403 20867 38409
rect 20809 38400 20821 38403
rect 20680 38372 20821 38400
rect 20680 38360 20686 38372
rect 20809 38369 20821 38372
rect 20855 38369 20867 38403
rect 20809 38363 20867 38369
rect 23664 38345 23722 38351
rect 22922 38332 22928 38344
rect 22664 38304 22928 38332
rect 21076 38267 21134 38273
rect 21076 38233 21088 38267
rect 21122 38264 21134 38267
rect 22554 38264 22560 38276
rect 21122 38236 22560 38264
rect 21122 38233 21134 38236
rect 21076 38227 21134 38233
rect 22554 38224 22560 38236
rect 22612 38224 22618 38276
rect 22664 38273 22692 38304
rect 22922 38292 22928 38304
rect 22980 38292 22986 38344
rect 23474 38292 23480 38344
rect 23532 38332 23538 38344
rect 23664 38334 23676 38345
rect 23584 38332 23676 38334
rect 23532 38311 23676 38332
rect 23710 38311 23722 38345
rect 23860 38341 23888 38428
rect 23952 38341 23980 38428
rect 24044 38351 24072 38440
rect 26142 38428 26148 38480
rect 26200 38468 26206 38480
rect 28077 38471 28135 38477
rect 28077 38468 28089 38471
rect 26200 38440 28089 38468
rect 26200 38428 26206 38440
rect 28077 38437 28089 38440
rect 28123 38437 28135 38471
rect 28077 38431 28135 38437
rect 30558 38428 30564 38480
rect 30616 38468 30622 38480
rect 32876 38468 32904 38496
rect 30616 38440 34100 38468
rect 30616 38428 30622 38440
rect 24854 38360 24860 38412
rect 24912 38400 24918 38412
rect 27522 38400 27528 38412
rect 24912 38372 27528 38400
rect 24912 38360 24918 38372
rect 24039 38345 24097 38351
rect 23532 38306 23722 38311
rect 23532 38304 23612 38306
rect 23664 38305 23722 38306
rect 23826 38335 23888 38341
rect 23532 38292 23538 38304
rect 23826 38301 23838 38335
rect 23872 38304 23888 38335
rect 23949 38335 24007 38341
rect 23872 38301 23884 38304
rect 23826 38295 23884 38301
rect 23949 38301 23961 38335
rect 23995 38301 24007 38335
rect 24039 38311 24051 38345
rect 24085 38311 24097 38345
rect 24039 38305 24097 38311
rect 24581 38335 24639 38341
rect 23949 38295 24007 38301
rect 24581 38301 24593 38335
rect 24627 38301 24639 38335
rect 24581 38295 24639 38301
rect 22649 38267 22707 38273
rect 22649 38233 22661 38267
rect 22695 38233 22707 38267
rect 23566 38264 23572 38276
rect 22649 38227 22707 38233
rect 23400 38236 23572 38264
rect 21266 38196 21272 38208
rect 20180 38168 21272 38196
rect 20073 38159 20131 38165
rect 21266 38156 21272 38168
rect 21324 38156 21330 38208
rect 22189 38199 22247 38205
rect 22189 38165 22201 38199
rect 22235 38196 22247 38199
rect 22462 38196 22468 38208
rect 22235 38168 22468 38196
rect 22235 38165 22247 38168
rect 22189 38159 22247 38165
rect 22462 38156 22468 38168
rect 22520 38156 22526 38208
rect 22830 38156 22836 38208
rect 22888 38205 22894 38208
rect 22888 38199 22907 38205
rect 22895 38196 22907 38199
rect 23400 38196 23428 38236
rect 23566 38224 23572 38236
rect 23624 38264 23630 38276
rect 24596 38264 24624 38295
rect 25958 38292 25964 38344
rect 26016 38332 26022 38344
rect 27448 38341 27476 38372
rect 27522 38360 27528 38372
rect 27580 38360 27586 38412
rect 31478 38400 31484 38412
rect 29932 38372 31484 38400
rect 27065 38335 27123 38341
rect 27065 38332 27077 38335
rect 26016 38304 27077 38332
rect 26016 38292 26022 38304
rect 27065 38301 27077 38304
rect 27111 38301 27123 38335
rect 27065 38295 27123 38301
rect 27433 38335 27491 38341
rect 27433 38301 27445 38335
rect 27479 38301 27491 38335
rect 27433 38295 27491 38301
rect 28077 38335 28135 38341
rect 28077 38301 28089 38335
rect 28123 38301 28135 38335
rect 28258 38332 28264 38344
rect 28219 38304 28264 38332
rect 28077 38295 28135 38301
rect 23624 38236 24624 38264
rect 23624 38224 23630 38236
rect 25498 38224 25504 38276
rect 25556 38264 25562 38276
rect 25685 38267 25743 38273
rect 25685 38264 25697 38267
rect 25556 38236 25697 38264
rect 25556 38224 25562 38236
rect 25685 38233 25697 38236
rect 25731 38233 25743 38267
rect 25685 38227 25743 38233
rect 26513 38267 26571 38273
rect 26513 38233 26525 38267
rect 26559 38233 26571 38267
rect 27246 38264 27252 38276
rect 27207 38236 27252 38264
rect 26513 38227 26571 38233
rect 22895 38168 23428 38196
rect 23477 38199 23535 38205
rect 22895 38165 22907 38168
rect 22888 38159 22907 38165
rect 23477 38165 23489 38199
rect 23523 38196 23535 38199
rect 24946 38196 24952 38208
rect 23523 38168 24952 38196
rect 23523 38165 23535 38168
rect 23477 38159 23535 38165
rect 22888 38156 22894 38159
rect 24946 38156 24952 38168
rect 25004 38156 25010 38208
rect 26528 38196 26556 38227
rect 27246 38224 27252 38236
rect 27304 38224 27310 38276
rect 27341 38267 27399 38273
rect 27341 38233 27353 38267
rect 27387 38264 27399 38267
rect 27706 38264 27712 38276
rect 27387 38236 27712 38264
rect 27387 38233 27399 38236
rect 27341 38227 27399 38233
rect 27706 38224 27712 38236
rect 27764 38264 27770 38276
rect 28092 38264 28120 38295
rect 28258 38292 28264 38304
rect 28316 38292 28322 38344
rect 29932 38341 29960 38372
rect 31478 38360 31484 38372
rect 31536 38360 31542 38412
rect 32493 38403 32551 38409
rect 32493 38369 32505 38403
rect 32539 38400 32551 38403
rect 33410 38400 33416 38412
rect 32539 38372 33416 38400
rect 32539 38369 32551 38372
rect 32493 38363 32551 38369
rect 33410 38360 33416 38372
rect 33468 38360 33474 38412
rect 29917 38335 29975 38341
rect 29917 38301 29929 38335
rect 29963 38301 29975 38335
rect 29917 38295 29975 38301
rect 30377 38335 30435 38341
rect 30377 38301 30389 38335
rect 30423 38332 30435 38335
rect 30558 38332 30564 38344
rect 30423 38304 30564 38332
rect 30423 38301 30435 38304
rect 30377 38295 30435 38301
rect 30558 38292 30564 38304
rect 30616 38332 30622 38344
rect 30837 38335 30895 38341
rect 30837 38332 30849 38335
rect 30616 38304 30849 38332
rect 30616 38292 30622 38304
rect 30837 38301 30849 38304
rect 30883 38301 30895 38335
rect 30837 38295 30895 38301
rect 31202 38292 31208 38344
rect 31260 38332 31266 38344
rect 31662 38332 31668 38344
rect 31260 38304 31668 38332
rect 31260 38292 31266 38304
rect 31662 38292 31668 38304
rect 31720 38332 31726 38344
rect 32585 38335 32643 38341
rect 32585 38332 32597 38335
rect 31720 38304 32597 38332
rect 31720 38292 31726 38304
rect 32585 38301 32597 38304
rect 32631 38301 32643 38335
rect 32585 38295 32643 38301
rect 33229 38335 33287 38341
rect 33229 38301 33241 38335
rect 33275 38301 33287 38335
rect 33229 38295 33287 38301
rect 28534 38264 28540 38276
rect 27764 38236 28540 38264
rect 27764 38224 27770 38236
rect 28534 38224 28540 38236
rect 28592 38224 28598 38276
rect 30009 38267 30067 38273
rect 30009 38233 30021 38267
rect 30055 38233 30067 38267
rect 30009 38227 30067 38233
rect 27062 38196 27068 38208
rect 26528 38168 27068 38196
rect 27062 38156 27068 38168
rect 27120 38156 27126 38208
rect 27614 38196 27620 38208
rect 27575 38168 27620 38196
rect 27614 38156 27620 38168
rect 27672 38156 27678 38208
rect 30024 38196 30052 38227
rect 30098 38224 30104 38276
rect 30156 38264 30162 38276
rect 30239 38267 30297 38273
rect 30156 38236 30201 38264
rect 30156 38224 30162 38236
rect 30239 38233 30251 38267
rect 30285 38264 30297 38267
rect 30466 38264 30472 38276
rect 30285 38236 30472 38264
rect 30285 38233 30297 38236
rect 30239 38227 30297 38233
rect 30466 38224 30472 38236
rect 30524 38224 30530 38276
rect 30926 38224 30932 38276
rect 30984 38264 30990 38276
rect 31021 38267 31079 38273
rect 31021 38264 31033 38267
rect 30984 38236 31033 38264
rect 30984 38224 30990 38236
rect 31021 38233 31033 38236
rect 31067 38264 31079 38267
rect 32306 38264 32312 38276
rect 31067 38236 31708 38264
rect 32267 38236 32312 38264
rect 31067 38233 31079 38236
rect 31021 38227 31079 38233
rect 31680 38208 31708 38236
rect 32306 38224 32312 38236
rect 32364 38224 32370 38276
rect 32950 38224 32956 38276
rect 33008 38264 33014 38276
rect 33244 38264 33272 38295
rect 33502 38292 33508 38344
rect 33560 38332 33566 38344
rect 34072 38341 34100 38440
rect 34146 38428 34152 38480
rect 34204 38468 34210 38480
rect 34204 38440 35204 38468
rect 34204 38428 34210 38440
rect 34238 38360 34244 38412
rect 34296 38400 34302 38412
rect 34333 38403 34391 38409
rect 34333 38400 34345 38403
rect 34296 38372 34345 38400
rect 34296 38360 34302 38372
rect 34333 38369 34345 38372
rect 34379 38369 34391 38403
rect 34333 38363 34391 38369
rect 35176 38400 35204 38440
rect 35434 38400 35440 38412
rect 35176 38372 35440 38400
rect 33597 38335 33655 38341
rect 33597 38332 33609 38335
rect 33560 38304 33609 38332
rect 33560 38292 33566 38304
rect 33597 38301 33609 38304
rect 33643 38301 33655 38335
rect 33597 38295 33655 38301
rect 34057 38335 34115 38341
rect 34057 38301 34069 38335
rect 34103 38301 34115 38335
rect 34057 38295 34115 38301
rect 34698 38292 34704 38344
rect 34756 38332 34762 38344
rect 35176 38341 35204 38372
rect 35434 38360 35440 38372
rect 35492 38360 35498 38412
rect 34885 38335 34943 38341
rect 34885 38332 34897 38335
rect 34756 38304 34897 38332
rect 34756 38292 34762 38304
rect 34885 38301 34897 38304
rect 34931 38301 34943 38335
rect 34885 38295 34943 38301
rect 35161 38335 35219 38341
rect 35161 38301 35173 38335
rect 35207 38301 35219 38335
rect 35161 38295 35219 38301
rect 35253 38335 35311 38341
rect 35253 38301 35265 38335
rect 35299 38301 35311 38335
rect 47670 38332 47676 38344
rect 47631 38304 47676 38332
rect 35253 38295 35311 38301
rect 34333 38267 34391 38273
rect 34333 38264 34345 38267
rect 33008 38236 34345 38264
rect 33008 38224 33014 38236
rect 34333 38233 34345 38236
rect 34379 38233 34391 38267
rect 34333 38227 34391 38233
rect 34422 38224 34428 38276
rect 34480 38264 34486 38276
rect 35069 38267 35127 38273
rect 35069 38264 35081 38267
rect 34480 38236 35081 38264
rect 34480 38224 34486 38236
rect 35069 38233 35081 38236
rect 35115 38233 35127 38267
rect 35268 38264 35296 38295
rect 47670 38292 47676 38304
rect 47728 38292 47734 38344
rect 35069 38227 35127 38233
rect 35176 38236 35296 38264
rect 30374 38196 30380 38208
rect 30024 38168 30380 38196
rect 30374 38156 30380 38168
rect 30432 38156 30438 38208
rect 30558 38156 30564 38208
rect 30616 38196 30622 38208
rect 31205 38199 31263 38205
rect 31205 38196 31217 38199
rect 30616 38168 31217 38196
rect 30616 38156 30622 38168
rect 31205 38165 31217 38168
rect 31251 38165 31263 38199
rect 31205 38159 31263 38165
rect 31662 38156 31668 38208
rect 31720 38156 31726 38208
rect 33042 38156 33048 38208
rect 33100 38196 33106 38208
rect 33321 38199 33379 38205
rect 33321 38196 33333 38199
rect 33100 38168 33333 38196
rect 33100 38156 33106 38168
rect 33321 38165 33333 38168
rect 33367 38165 33379 38199
rect 33321 38159 33379 38165
rect 33505 38199 33563 38205
rect 33505 38165 33517 38199
rect 33551 38196 33563 38199
rect 33870 38196 33876 38208
rect 33551 38168 33876 38196
rect 33551 38165 33563 38168
rect 33505 38159 33563 38165
rect 33870 38156 33876 38168
rect 33928 38156 33934 38208
rect 34238 38156 34244 38208
rect 34296 38196 34302 38208
rect 35176 38196 35204 38236
rect 34296 38168 35204 38196
rect 34296 38156 34302 38168
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 15197 37995 15255 38001
rect 15197 37961 15209 37995
rect 15243 37992 15255 37995
rect 15470 37992 15476 38004
rect 15243 37964 15476 37992
rect 15243 37961 15255 37964
rect 15197 37955 15255 37961
rect 15470 37952 15476 37964
rect 15528 37952 15534 38004
rect 17494 37992 17500 38004
rect 17455 37964 17500 37992
rect 17494 37952 17500 37964
rect 17552 37952 17558 38004
rect 19521 37995 19579 38001
rect 19521 37961 19533 37995
rect 19567 37992 19579 37995
rect 20254 37992 20260 38004
rect 19567 37964 20260 37992
rect 19567 37961 19579 37964
rect 19521 37955 19579 37961
rect 20254 37952 20260 37964
rect 20312 37952 20318 38004
rect 24854 37992 24860 38004
rect 23769 37964 24860 37992
rect 20272 37924 20300 37952
rect 22373 37927 22431 37933
rect 20272 37896 22140 37924
rect 12894 37856 12900 37868
rect 12855 37828 12900 37856
rect 12894 37816 12900 37828
rect 12952 37816 12958 37868
rect 15378 37856 15384 37868
rect 15339 37828 15384 37856
rect 15378 37816 15384 37828
rect 15436 37816 15442 37868
rect 15562 37856 15568 37868
rect 15523 37828 15568 37856
rect 15562 37816 15568 37828
rect 15620 37856 15626 37868
rect 17678 37856 17684 37868
rect 15620 37828 16436 37856
rect 17639 37828 17684 37856
rect 15620 37816 15626 37828
rect 15654 37788 15660 37800
rect 15615 37760 15660 37788
rect 15654 37748 15660 37760
rect 15712 37748 15718 37800
rect 16408 37788 16436 37828
rect 17678 37816 17684 37828
rect 17736 37816 17742 37868
rect 17954 37856 17960 37868
rect 17915 37828 17960 37856
rect 17954 37816 17960 37828
rect 18012 37816 18018 37868
rect 18690 37816 18696 37868
rect 18748 37856 18754 37868
rect 19245 37859 19303 37865
rect 19245 37856 19257 37859
rect 18748 37828 19257 37856
rect 18748 37816 18754 37828
rect 19245 37825 19257 37828
rect 19291 37825 19303 37859
rect 19245 37819 19303 37825
rect 20162 37816 20168 37868
rect 20220 37856 20226 37868
rect 20329 37859 20387 37865
rect 20329 37856 20341 37859
rect 20220 37828 20341 37856
rect 20220 37816 20226 37828
rect 20329 37825 20341 37828
rect 20375 37825 20387 37859
rect 20329 37819 20387 37825
rect 17218 37788 17224 37800
rect 16408 37760 17224 37788
rect 17218 37748 17224 37760
rect 17276 37788 17282 37800
rect 17865 37791 17923 37797
rect 17865 37788 17877 37791
rect 17276 37760 17877 37788
rect 17276 37748 17282 37760
rect 17865 37757 17877 37760
rect 17911 37757 17923 37791
rect 20070 37788 20076 37800
rect 20031 37760 20076 37788
rect 17865 37751 17923 37757
rect 20070 37748 20076 37760
rect 20128 37748 20134 37800
rect 22112 37788 22140 37896
rect 22373 37893 22385 37927
rect 22419 37924 22431 37927
rect 22738 37924 22744 37936
rect 22419 37896 22744 37924
rect 22419 37893 22431 37896
rect 22373 37887 22431 37893
rect 22738 37884 22744 37896
rect 22796 37884 22802 37936
rect 22189 37859 22247 37865
rect 22189 37825 22201 37859
rect 22235 37856 22247 37859
rect 22278 37856 22284 37868
rect 22235 37828 22284 37856
rect 22235 37825 22247 37828
rect 22189 37819 22247 37825
rect 22278 37816 22284 37828
rect 22336 37816 22342 37868
rect 22462 37856 22468 37868
rect 22423 37828 22468 37856
rect 22462 37816 22468 37828
rect 22520 37816 22526 37868
rect 22557 37859 22615 37865
rect 22557 37825 22569 37859
rect 22603 37856 22615 37859
rect 23769 37856 23797 37964
rect 24854 37952 24860 37964
rect 24912 37952 24918 38004
rect 25314 37992 25320 38004
rect 25275 37964 25320 37992
rect 25314 37952 25320 37964
rect 25372 37952 25378 38004
rect 28534 37992 28540 38004
rect 28495 37964 28540 37992
rect 28534 37952 28540 37964
rect 28592 37952 28598 38004
rect 30561 37995 30619 38001
rect 30561 37961 30573 37995
rect 30607 37992 30619 37995
rect 31202 37992 31208 38004
rect 30607 37964 31208 37992
rect 30607 37961 30619 37964
rect 30561 37955 30619 37961
rect 31202 37952 31208 37964
rect 31260 37952 31266 38004
rect 32398 37952 32404 38004
rect 32456 37992 32462 38004
rect 32861 37995 32919 38001
rect 32861 37992 32873 37995
rect 32456 37964 32873 37992
rect 32456 37952 32462 37964
rect 32861 37961 32873 37964
rect 32907 37992 32919 37995
rect 33042 37992 33048 38004
rect 32907 37964 33048 37992
rect 32907 37961 32919 37964
rect 32861 37955 32919 37961
rect 33042 37952 33048 37964
rect 33100 37952 33106 38004
rect 26050 37924 26056 37936
rect 25516 37896 26056 37924
rect 22603 37828 23797 37856
rect 22603 37825 22615 37828
rect 22557 37819 22615 37825
rect 22572 37788 22600 37819
rect 23842 37816 23848 37868
rect 23900 37856 23906 37868
rect 25516 37865 25544 37896
rect 26050 37884 26056 37896
rect 26108 37924 26114 37936
rect 27424 37927 27482 37933
rect 26108 37896 26648 37924
rect 26108 37884 26114 37896
rect 25501 37859 25559 37865
rect 23900 37828 23945 37856
rect 23900 37816 23906 37828
rect 25501 37825 25513 37859
rect 25547 37825 25559 37859
rect 25774 37856 25780 37868
rect 25735 37828 25780 37856
rect 25501 37819 25559 37825
rect 25774 37816 25780 37828
rect 25832 37816 25838 37868
rect 25961 37859 26019 37865
rect 25961 37825 25973 37859
rect 26007 37856 26019 37859
rect 26142 37856 26148 37868
rect 26007 37828 26148 37856
rect 26007 37825 26019 37828
rect 25961 37819 26019 37825
rect 26142 37816 26148 37828
rect 26200 37856 26206 37868
rect 26620 37865 26648 37896
rect 27424 37893 27436 37927
rect 27470 37924 27482 37927
rect 27614 37924 27620 37936
rect 27470 37896 27620 37924
rect 27470 37893 27482 37896
rect 27424 37887 27482 37893
rect 27614 37884 27620 37896
rect 27672 37884 27678 37936
rect 30650 37924 30656 37936
rect 30392 37896 30656 37924
rect 26421 37859 26479 37865
rect 26421 37856 26433 37859
rect 26200 37828 26433 37856
rect 26200 37816 26206 37828
rect 26421 37825 26433 37828
rect 26467 37825 26479 37859
rect 26421 37819 26479 37825
rect 26605 37859 26663 37865
rect 26605 37825 26617 37859
rect 26651 37856 26663 37859
rect 27890 37856 27896 37868
rect 26651 37828 27896 37856
rect 26651 37825 26663 37828
rect 26605 37819 26663 37825
rect 27890 37816 27896 37828
rect 27948 37816 27954 37868
rect 30392 37865 30420 37896
rect 30650 37884 30656 37896
rect 30708 37884 30714 37936
rect 33410 37924 33416 37936
rect 32692 37896 33416 37924
rect 30377 37859 30435 37865
rect 30377 37825 30389 37859
rect 30423 37825 30435 37859
rect 30558 37856 30564 37868
rect 30519 37828 30564 37856
rect 30377 37819 30435 37825
rect 30558 37816 30564 37828
rect 30616 37816 30622 37868
rect 32692 37865 32720 37896
rect 33410 37884 33416 37896
rect 33468 37884 33474 37936
rect 34146 37924 34152 37936
rect 34107 37896 34152 37924
rect 34146 37884 34152 37896
rect 34204 37884 34210 37936
rect 32677 37859 32735 37865
rect 32677 37825 32689 37859
rect 32723 37825 32735 37859
rect 32677 37819 32735 37825
rect 32950 37816 32956 37868
rect 33008 37856 33014 37868
rect 33870 37856 33876 37868
rect 33008 37828 33053 37856
rect 33831 37828 33876 37856
rect 33008 37816 33014 37828
rect 33870 37816 33876 37828
rect 33928 37816 33934 37868
rect 34057 37859 34115 37865
rect 34057 37825 34069 37859
rect 34103 37825 34115 37859
rect 34057 37819 34115 37825
rect 34241 37859 34299 37865
rect 34241 37825 34253 37859
rect 34287 37856 34299 37859
rect 34330 37856 34336 37868
rect 34287 37828 34336 37856
rect 34287 37825 34299 37828
rect 34241 37819 34299 37825
rect 22112 37760 22600 37788
rect 23474 37748 23480 37800
rect 23532 37788 23538 37800
rect 23661 37791 23719 37797
rect 23661 37788 23673 37791
rect 23532 37760 23673 37788
rect 23532 37748 23538 37760
rect 23661 37757 23673 37760
rect 23707 37757 23719 37791
rect 23661 37751 23719 37757
rect 23753 37791 23811 37797
rect 23753 37757 23765 37791
rect 23799 37757 23811 37791
rect 23753 37751 23811 37757
rect 22554 37680 22560 37732
rect 22612 37720 22618 37732
rect 22741 37723 22799 37729
rect 22741 37720 22753 37723
rect 22612 37692 22753 37720
rect 22612 37680 22618 37692
rect 22741 37689 22753 37692
rect 22787 37689 22799 37723
rect 22741 37683 22799 37689
rect 23106 37680 23112 37732
rect 23164 37720 23170 37732
rect 23768 37720 23796 37751
rect 23934 37748 23940 37800
rect 23992 37788 23998 37800
rect 23992 37760 24037 37788
rect 23992 37748 23998 37760
rect 27062 37748 27068 37800
rect 27120 37788 27126 37800
rect 27157 37791 27215 37797
rect 27157 37788 27169 37791
rect 27120 37760 27169 37788
rect 27120 37748 27126 37760
rect 27157 37757 27169 37760
rect 27203 37757 27215 37791
rect 34072 37788 34100 37819
rect 34330 37816 34336 37828
rect 34388 37816 34394 37868
rect 47762 37856 47768 37868
rect 47723 37828 47768 37856
rect 47762 37816 47768 37828
rect 47820 37816 47826 37868
rect 27157 37751 27215 37757
rect 32968 37760 34100 37788
rect 23164 37692 23796 37720
rect 23164 37680 23170 37692
rect 32968 37664 32996 37760
rect 12618 37612 12624 37664
rect 12676 37652 12682 37664
rect 12713 37655 12771 37661
rect 12713 37652 12725 37655
rect 12676 37624 12725 37652
rect 12676 37612 12682 37624
rect 12713 37621 12725 37624
rect 12759 37621 12771 37655
rect 12713 37615 12771 37621
rect 21453 37655 21511 37661
rect 21453 37621 21465 37655
rect 21499 37652 21511 37655
rect 21726 37652 21732 37664
rect 21499 37624 21732 37652
rect 21499 37621 21511 37624
rect 21453 37615 21511 37621
rect 21726 37612 21732 37624
rect 21784 37612 21790 37664
rect 23477 37655 23535 37661
rect 23477 37621 23489 37655
rect 23523 37652 23535 37655
rect 24762 37652 24768 37664
rect 23523 37624 24768 37652
rect 23523 37621 23535 37624
rect 23477 37615 23535 37621
rect 24762 37612 24768 37624
rect 24820 37612 24826 37664
rect 26418 37652 26424 37664
rect 26379 37624 26424 37652
rect 26418 37612 26424 37624
rect 26476 37612 26482 37664
rect 32493 37655 32551 37661
rect 32493 37621 32505 37655
rect 32539 37652 32551 37655
rect 32950 37652 32956 37664
rect 32539 37624 32956 37652
rect 32539 37621 32551 37624
rect 32493 37615 32551 37621
rect 32950 37612 32956 37624
rect 33008 37612 33014 37664
rect 34425 37655 34483 37661
rect 34425 37621 34437 37655
rect 34471 37652 34483 37655
rect 34698 37652 34704 37664
rect 34471 37624 34704 37652
rect 34471 37621 34483 37624
rect 34425 37615 34483 37621
rect 34698 37612 34704 37624
rect 34756 37612 34762 37664
rect 47854 37652 47860 37664
rect 47815 37624 47860 37652
rect 47854 37612 47860 37624
rect 47912 37612 47918 37664
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 16850 37408 16856 37460
rect 16908 37448 16914 37460
rect 17313 37451 17371 37457
rect 17313 37448 17325 37451
rect 16908 37420 17325 37448
rect 16908 37408 16914 37420
rect 17313 37417 17325 37420
rect 17359 37417 17371 37451
rect 17313 37411 17371 37417
rect 18693 37451 18751 37457
rect 18693 37417 18705 37451
rect 18739 37448 18751 37451
rect 19978 37448 19984 37460
rect 18739 37420 19984 37448
rect 18739 37417 18751 37420
rect 18693 37411 18751 37417
rect 19978 37408 19984 37420
rect 20036 37408 20042 37460
rect 22646 37448 22652 37460
rect 22607 37420 22652 37448
rect 22646 37408 22652 37420
rect 22704 37408 22710 37460
rect 23474 37448 23480 37460
rect 22756 37420 23244 37448
rect 23435 37420 23480 37448
rect 22462 37340 22468 37392
rect 22520 37380 22526 37392
rect 22756 37380 22784 37420
rect 22520 37352 22784 37380
rect 22520 37340 22526 37352
rect 15654 37312 15660 37324
rect 13832 37284 15660 37312
rect 1578 37244 1584 37256
rect 1539 37216 1584 37244
rect 1578 37204 1584 37216
rect 1636 37204 1642 37256
rect 12342 37244 12348 37256
rect 12303 37216 12348 37244
rect 12342 37204 12348 37216
rect 12400 37204 12406 37256
rect 12618 37253 12624 37256
rect 12612 37244 12624 37253
rect 12579 37216 12624 37244
rect 12612 37207 12624 37216
rect 12618 37204 12624 37207
rect 12676 37204 12682 37256
rect 13832 37244 13860 37284
rect 15654 37272 15660 37284
rect 15712 37272 15718 37324
rect 13372 37216 13860 37244
rect 16945 37247 17003 37253
rect 12434 37176 12440 37188
rect 6886 37148 12440 37176
rect 1765 37111 1823 37117
rect 1765 37077 1777 37111
rect 1811 37108 1823 37111
rect 6886 37108 6914 37148
rect 12434 37136 12440 37148
rect 12492 37176 12498 37188
rect 13372 37176 13400 37216
rect 16945 37213 16957 37247
rect 16991 37244 17003 37247
rect 16991 37216 17816 37244
rect 16991 37213 17003 37216
rect 16945 37207 17003 37213
rect 12492 37148 13400 37176
rect 17129 37179 17187 37185
rect 12492 37136 12498 37148
rect 17129 37145 17141 37179
rect 17175 37145 17187 37179
rect 17788 37176 17816 37216
rect 17862 37204 17868 37256
rect 17920 37244 17926 37256
rect 18141 37247 18199 37253
rect 17920 37216 17965 37244
rect 17920 37204 17926 37216
rect 18141 37213 18153 37247
rect 18187 37213 18199 37247
rect 18141 37207 18199 37213
rect 18233 37247 18291 37253
rect 18233 37213 18245 37247
rect 18279 37244 18291 37247
rect 18690 37244 18696 37256
rect 18279 37216 18696 37244
rect 18279 37213 18291 37216
rect 18233 37207 18291 37213
rect 18156 37176 18184 37207
rect 18690 37204 18696 37216
rect 18748 37204 18754 37256
rect 18877 37247 18935 37253
rect 18877 37213 18889 37247
rect 18923 37213 18935 37247
rect 18877 37207 18935 37213
rect 18892 37176 18920 37207
rect 19334 37204 19340 37256
rect 19392 37244 19398 37256
rect 20070 37244 20076 37256
rect 19392 37216 20076 37244
rect 19392 37204 19398 37216
rect 20070 37204 20076 37216
rect 20128 37244 20134 37256
rect 20165 37247 20223 37253
rect 20165 37244 20177 37247
rect 20128 37216 20177 37244
rect 20128 37204 20134 37216
rect 20165 37213 20177 37216
rect 20211 37213 20223 37247
rect 21266 37244 21272 37256
rect 21227 37216 21272 37244
rect 20165 37207 20223 37213
rect 21266 37204 21272 37216
rect 21324 37204 21330 37256
rect 21542 37244 21548 37256
rect 21503 37216 21548 37244
rect 21542 37204 21548 37216
rect 21600 37204 21606 37256
rect 21726 37244 21732 37256
rect 21687 37216 21732 37244
rect 21726 37204 21732 37216
rect 21784 37204 21790 37256
rect 22925 37247 22983 37253
rect 22925 37213 22937 37247
rect 22971 37238 22983 37247
rect 23106 37244 23112 37256
rect 23032 37238 23112 37244
rect 22971 37216 23112 37238
rect 22971 37213 23060 37216
rect 22925 37210 23060 37213
rect 22925 37207 22983 37210
rect 23106 37204 23112 37216
rect 23164 37204 23170 37256
rect 23216 37244 23244 37420
rect 23474 37408 23480 37420
rect 23532 37408 23538 37460
rect 27065 37451 27123 37457
rect 27065 37417 27077 37451
rect 27111 37448 27123 37451
rect 27246 37448 27252 37460
rect 27111 37420 27252 37448
rect 27111 37417 27123 37420
rect 27065 37411 27123 37417
rect 27246 37408 27252 37420
rect 27304 37408 27310 37460
rect 27890 37448 27896 37460
rect 27851 37420 27896 37448
rect 27890 37408 27896 37420
rect 27948 37408 27954 37460
rect 33410 37408 33416 37460
rect 33468 37448 33474 37460
rect 33781 37451 33839 37457
rect 33781 37448 33793 37451
rect 33468 37420 33793 37448
rect 33468 37408 33474 37420
rect 33781 37417 33793 37420
rect 33827 37417 33839 37451
rect 33781 37411 33839 37417
rect 25774 37272 25780 37324
rect 25832 37312 25838 37324
rect 25961 37315 26019 37321
rect 25961 37312 25973 37315
rect 25832 37284 25973 37312
rect 25832 37272 25838 37284
rect 25961 37281 25973 37284
rect 26007 37281 26019 37315
rect 25961 37275 26019 37281
rect 26053 37315 26111 37321
rect 26053 37281 26065 37315
rect 26099 37312 26111 37315
rect 26418 37312 26424 37324
rect 26099 37284 26424 37312
rect 26099 37281 26111 37284
rect 26053 37275 26111 37281
rect 26418 37272 26424 37284
rect 26476 37272 26482 37324
rect 27525 37315 27583 37321
rect 27525 37281 27537 37315
rect 27571 37312 27583 37315
rect 28258 37312 28264 37324
rect 27571 37284 28264 37312
rect 27571 37281 27583 37284
rect 27525 37275 27583 37281
rect 28258 37272 28264 37284
rect 28316 37272 28322 37324
rect 48222 37312 48228 37324
rect 48183 37284 48228 37312
rect 48222 37272 48228 37284
rect 48280 37272 48286 37324
rect 23385 37247 23443 37253
rect 23385 37244 23397 37247
rect 23216 37216 23397 37244
rect 23385 37213 23397 37216
rect 23431 37213 23443 37247
rect 23566 37244 23572 37256
rect 23527 37216 23572 37244
rect 23385 37207 23443 37213
rect 23566 37204 23572 37216
rect 23624 37204 23630 37256
rect 24762 37204 24768 37256
rect 24820 37244 24826 37256
rect 24857 37247 24915 37253
rect 24857 37244 24869 37247
rect 24820 37216 24869 37244
rect 24820 37204 24826 37216
rect 24857 37213 24869 37216
rect 24903 37213 24915 37247
rect 24857 37207 24915 37213
rect 25225 37247 25283 37253
rect 25225 37213 25237 37247
rect 25271 37244 25283 37247
rect 25866 37244 25872 37256
rect 25271 37216 25872 37244
rect 25271 37213 25283 37216
rect 25225 37207 25283 37213
rect 25866 37204 25872 37216
rect 25924 37204 25930 37256
rect 26145 37247 26203 37253
rect 26145 37213 26157 37247
rect 26191 37213 26203 37247
rect 27706 37244 27712 37256
rect 27667 37216 27712 37244
rect 26145 37207 26203 37213
rect 19426 37176 19432 37188
rect 17788 37148 18920 37176
rect 19387 37148 19432 37176
rect 17129 37139 17187 37145
rect 1811 37080 6914 37108
rect 1811 37077 1823 37080
rect 1765 37071 1823 37077
rect 13630 37068 13636 37120
rect 13688 37108 13694 37120
rect 13725 37111 13783 37117
rect 13725 37108 13737 37111
rect 13688 37080 13737 37108
rect 13688 37068 13694 37080
rect 13725 37077 13737 37080
rect 13771 37077 13783 37111
rect 13725 37071 13783 37077
rect 16942 37068 16948 37120
rect 17000 37108 17006 37120
rect 17144 37108 17172 37139
rect 17770 37108 17776 37120
rect 17000 37080 17776 37108
rect 17000 37068 17006 37080
rect 17770 37068 17776 37080
rect 17828 37068 17834 37120
rect 18892 37108 18920 37148
rect 19426 37136 19432 37148
rect 19484 37136 19490 37188
rect 22646 37176 22652 37188
rect 19536 37148 22094 37176
rect 22607 37148 22652 37176
rect 19536 37108 19564 37148
rect 18892 37080 19564 37108
rect 20346 37068 20352 37120
rect 20404 37108 20410 37120
rect 21085 37111 21143 37117
rect 21085 37108 21097 37111
rect 20404 37080 21097 37108
rect 20404 37068 20410 37080
rect 21085 37077 21097 37080
rect 21131 37077 21143 37111
rect 22066 37108 22094 37148
rect 22646 37136 22652 37148
rect 22704 37136 22710 37188
rect 22830 37136 22836 37188
rect 22888 37176 22894 37188
rect 25038 37176 25044 37188
rect 22888 37148 22933 37176
rect 24999 37148 25044 37176
rect 22888 37136 22894 37148
rect 25038 37136 25044 37148
rect 25096 37136 25102 37188
rect 26160 37176 26188 37207
rect 27706 37204 27712 37216
rect 27764 37204 27770 37256
rect 31662 37204 31668 37256
rect 31720 37244 31726 37256
rect 33045 37247 33103 37253
rect 33045 37244 33057 37247
rect 31720 37216 33057 37244
rect 31720 37204 31726 37216
rect 33045 37213 33057 37216
rect 33091 37213 33103 37247
rect 33045 37207 33103 37213
rect 33229 37247 33287 37253
rect 33229 37213 33241 37247
rect 33275 37244 33287 37247
rect 33689 37247 33747 37253
rect 33689 37244 33701 37247
rect 33275 37216 33701 37244
rect 33275 37213 33287 37216
rect 33229 37207 33287 37213
rect 33689 37213 33701 37216
rect 33735 37213 33747 37247
rect 33870 37244 33876 37256
rect 33831 37216 33876 37244
rect 33689 37207 33747 37213
rect 25608 37148 26188 37176
rect 26697 37179 26755 37185
rect 25130 37108 25136 37120
rect 22066 37080 25136 37108
rect 21085 37071 21143 37077
rect 25130 37068 25136 37080
rect 25188 37108 25194 37120
rect 25608 37108 25636 37148
rect 26697 37145 26709 37179
rect 26743 37145 26755 37179
rect 26878 37176 26884 37188
rect 26839 37148 26884 37176
rect 26697 37139 26755 37145
rect 25188 37080 25636 37108
rect 25685 37111 25743 37117
rect 25188 37068 25194 37080
rect 25685 37077 25697 37111
rect 25731 37108 25743 37111
rect 26712 37108 26740 37139
rect 26878 37136 26884 37148
rect 26936 37136 26942 37188
rect 32861 37179 32919 37185
rect 32861 37145 32873 37179
rect 32907 37145 32919 37179
rect 33060 37176 33088 37207
rect 33870 37204 33876 37216
rect 33928 37204 33934 37256
rect 34790 37204 34796 37256
rect 34848 37244 34854 37256
rect 34885 37247 34943 37253
rect 34885 37244 34897 37247
rect 34848 37216 34897 37244
rect 34848 37204 34854 37216
rect 34885 37213 34897 37216
rect 34931 37244 34943 37247
rect 36630 37244 36636 37256
rect 34931 37216 36636 37244
rect 34931 37213 34943 37216
rect 34885 37207 34943 37213
rect 36630 37204 36636 37216
rect 36688 37204 36694 37256
rect 46477 37247 46535 37253
rect 46477 37213 46489 37247
rect 46523 37213 46535 37247
rect 46477 37207 46535 37213
rect 33594 37176 33600 37188
rect 33060 37148 33600 37176
rect 32861 37139 32919 37145
rect 25731 37080 26740 37108
rect 32876 37108 32904 37139
rect 33594 37136 33600 37148
rect 33652 37136 33658 37188
rect 34698 37136 34704 37188
rect 34756 37176 34762 37188
rect 35130 37179 35188 37185
rect 35130 37176 35142 37179
rect 34756 37148 35142 37176
rect 34756 37136 34762 37148
rect 35130 37145 35142 37148
rect 35176 37145 35188 37179
rect 35130 37139 35188 37145
rect 33134 37108 33140 37120
rect 32876 37080 33140 37108
rect 25731 37077 25743 37080
rect 25685 37071 25743 37077
rect 33134 37068 33140 37080
rect 33192 37108 33198 37120
rect 33410 37108 33416 37120
rect 33192 37080 33416 37108
rect 33192 37068 33198 37080
rect 33410 37068 33416 37080
rect 33468 37108 33474 37120
rect 34146 37108 34152 37120
rect 33468 37080 34152 37108
rect 33468 37068 33474 37080
rect 34146 37068 34152 37080
rect 34204 37108 34210 37120
rect 36265 37111 36323 37117
rect 36265 37108 36277 37111
rect 34204 37080 36277 37108
rect 34204 37068 34210 37080
rect 36265 37077 36277 37080
rect 36311 37077 36323 37111
rect 46492 37108 46520 37207
rect 46661 37179 46719 37185
rect 46661 37145 46673 37179
rect 46707 37176 46719 37179
rect 47854 37176 47860 37188
rect 46707 37148 47860 37176
rect 46707 37145 46719 37148
rect 46661 37139 46719 37145
rect 47854 37136 47860 37148
rect 47912 37136 47918 37188
rect 47670 37108 47676 37120
rect 46492 37080 47676 37108
rect 36265 37071 36323 37077
rect 47670 37068 47676 37080
rect 47728 37068 47734 37120
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 1762 36864 1768 36916
rect 1820 36904 1826 36916
rect 1820 36876 6914 36904
rect 1820 36864 1826 36876
rect 6886 36836 6914 36876
rect 12894 36864 12900 36916
rect 12952 36904 12958 36916
rect 13265 36907 13323 36913
rect 13265 36904 13277 36907
rect 12952 36876 13277 36904
rect 12952 36864 12958 36876
rect 13265 36873 13277 36876
rect 13311 36873 13323 36907
rect 13630 36904 13636 36916
rect 13591 36876 13636 36904
rect 13265 36867 13323 36873
rect 13630 36864 13636 36876
rect 13688 36864 13694 36916
rect 13725 36907 13783 36913
rect 13725 36873 13737 36907
rect 13771 36904 13783 36907
rect 15565 36907 15623 36913
rect 15565 36904 15577 36907
rect 13771 36876 15577 36904
rect 13771 36873 13783 36876
rect 13725 36867 13783 36873
rect 15565 36873 15577 36876
rect 15611 36873 15623 36907
rect 15565 36867 15623 36873
rect 15933 36907 15991 36913
rect 15933 36873 15945 36907
rect 15979 36904 15991 36907
rect 16114 36904 16120 36916
rect 15979 36876 16120 36904
rect 15979 36873 15991 36876
rect 15933 36867 15991 36873
rect 16114 36864 16120 36876
rect 16172 36864 16178 36916
rect 20809 36907 20867 36913
rect 20809 36904 20821 36907
rect 19352 36876 20821 36904
rect 18322 36836 18328 36848
rect 6886 36808 18328 36836
rect 18322 36796 18328 36808
rect 18380 36796 18386 36848
rect 18592 36839 18650 36845
rect 18592 36805 18604 36839
rect 18638 36836 18650 36839
rect 19352 36836 19380 36876
rect 20809 36873 20821 36876
rect 20855 36873 20867 36907
rect 20809 36867 20867 36873
rect 21726 36864 21732 36916
rect 21784 36864 21790 36916
rect 22649 36907 22707 36913
rect 22649 36873 22661 36907
rect 22695 36904 22707 36907
rect 23382 36904 23388 36916
rect 22695 36876 23388 36904
rect 22695 36873 22707 36876
rect 22649 36867 22707 36873
rect 23382 36864 23388 36876
rect 23440 36864 23446 36916
rect 26059 36907 26117 36913
rect 26059 36873 26071 36907
rect 26105 36904 26117 36907
rect 26878 36904 26884 36916
rect 26105 36876 26884 36904
rect 26105 36873 26117 36876
rect 26059 36867 26117 36873
rect 26878 36864 26884 36876
rect 26936 36864 26942 36916
rect 29917 36907 29975 36913
rect 29917 36873 29929 36907
rect 29963 36904 29975 36907
rect 31662 36904 31668 36916
rect 29963 36876 31668 36904
rect 29963 36873 29975 36876
rect 29917 36867 29975 36873
rect 31662 36864 31668 36876
rect 31720 36864 31726 36916
rect 32861 36907 32919 36913
rect 32861 36873 32873 36907
rect 32907 36904 32919 36907
rect 33597 36907 33655 36913
rect 33597 36904 33609 36907
rect 32907 36876 33609 36904
rect 32907 36873 32919 36876
rect 32861 36867 32919 36873
rect 33597 36873 33609 36876
rect 33643 36904 33655 36907
rect 33686 36904 33692 36916
rect 33643 36876 33692 36904
rect 33643 36873 33655 36876
rect 33597 36867 33655 36873
rect 33686 36864 33692 36876
rect 33744 36904 33750 36916
rect 33870 36904 33876 36916
rect 33744 36876 33876 36904
rect 33744 36864 33750 36876
rect 33870 36864 33876 36876
rect 33928 36864 33934 36916
rect 18638 36808 19380 36836
rect 18638 36805 18650 36808
rect 18592 36799 18650 36805
rect 20070 36796 20076 36848
rect 20128 36836 20134 36848
rect 20441 36839 20499 36845
rect 20441 36836 20453 36839
rect 20128 36808 20453 36836
rect 20128 36796 20134 36808
rect 20441 36805 20453 36808
rect 20487 36805 20499 36839
rect 21744 36836 21772 36864
rect 23566 36836 23572 36848
rect 21744 36808 23572 36836
rect 20441 36799 20499 36805
rect 17126 36768 17132 36780
rect 14108 36740 17132 36768
rect 14108 36712 14136 36740
rect 17126 36728 17132 36740
rect 17184 36728 17190 36780
rect 18414 36728 18420 36780
rect 18472 36768 18478 36780
rect 19886 36768 19892 36780
rect 18472 36740 19892 36768
rect 18472 36728 18478 36740
rect 19886 36728 19892 36740
rect 19944 36728 19950 36780
rect 19978 36728 19984 36780
rect 20036 36768 20042 36780
rect 20165 36771 20223 36777
rect 20165 36768 20177 36771
rect 20036 36740 20177 36768
rect 20036 36728 20042 36740
rect 20165 36737 20177 36740
rect 20211 36737 20223 36771
rect 20165 36731 20223 36737
rect 20258 36774 20316 36777
rect 20258 36771 20372 36774
rect 20258 36737 20270 36771
rect 20304 36746 20372 36771
rect 20304 36737 20316 36746
rect 20258 36731 20316 36737
rect 13909 36703 13967 36709
rect 13909 36669 13921 36703
rect 13955 36700 13967 36703
rect 14090 36700 14096 36712
rect 13955 36672 14096 36700
rect 13955 36669 13967 36672
rect 13909 36663 13967 36669
rect 14090 36660 14096 36672
rect 14148 36660 14154 36712
rect 16022 36700 16028 36712
rect 15983 36672 16028 36700
rect 16022 36660 16028 36672
rect 16080 36660 16086 36712
rect 16114 36660 16120 36712
rect 16172 36700 16178 36712
rect 18325 36703 18383 36709
rect 16172 36672 16217 36700
rect 16172 36660 16178 36672
rect 18325 36669 18337 36703
rect 18371 36669 18383 36703
rect 18325 36663 18383 36669
rect 18340 36564 18368 36663
rect 19426 36564 19432 36576
rect 18340 36536 19432 36564
rect 19426 36524 19432 36536
rect 19484 36524 19490 36576
rect 19702 36564 19708 36576
rect 19663 36536 19708 36564
rect 19702 36524 19708 36536
rect 19760 36564 19766 36576
rect 20344 36564 20372 36746
rect 20533 36771 20591 36777
rect 20533 36737 20545 36771
rect 20579 36737 20591 36771
rect 20533 36731 20591 36737
rect 20548 36644 20576 36731
rect 20622 36728 20628 36780
rect 20680 36777 20686 36780
rect 20680 36768 20688 36777
rect 21726 36768 21732 36780
rect 20680 36740 21732 36768
rect 20680 36731 20688 36740
rect 20680 36728 20686 36731
rect 21726 36728 21732 36740
rect 21784 36728 21790 36780
rect 22462 36728 22468 36780
rect 22520 36768 22526 36780
rect 22756 36777 22784 36808
rect 23566 36796 23572 36808
rect 23624 36796 23630 36848
rect 25961 36839 26019 36845
rect 25961 36805 25973 36839
rect 26007 36836 26019 36839
rect 26418 36836 26424 36848
rect 26007 36808 26424 36836
rect 26007 36805 26019 36808
rect 25961 36799 26019 36805
rect 26418 36796 26424 36808
rect 26476 36796 26482 36848
rect 22557 36771 22615 36777
rect 22557 36768 22569 36771
rect 22520 36740 22569 36768
rect 22520 36728 22526 36740
rect 22557 36737 22569 36740
rect 22603 36737 22615 36771
rect 22557 36731 22615 36737
rect 22741 36771 22799 36777
rect 22741 36737 22753 36771
rect 22787 36737 22799 36771
rect 24578 36768 24584 36780
rect 24491 36740 24584 36768
rect 22741 36731 22799 36737
rect 24578 36728 24584 36740
rect 24636 36768 24642 36780
rect 25498 36768 25504 36780
rect 24636 36740 25504 36768
rect 24636 36728 24642 36740
rect 25498 36728 25504 36740
rect 25556 36728 25562 36780
rect 25774 36728 25780 36780
rect 25832 36768 25838 36780
rect 26145 36771 26203 36777
rect 26145 36768 26157 36771
rect 25832 36740 26157 36768
rect 25832 36728 25838 36740
rect 26145 36737 26157 36740
rect 26191 36737 26203 36771
rect 26145 36731 26203 36737
rect 26237 36771 26295 36777
rect 26237 36737 26249 36771
rect 26283 36737 26295 36771
rect 26237 36731 26295 36737
rect 22002 36660 22008 36712
rect 22060 36700 22066 36712
rect 25317 36703 25375 36709
rect 25317 36700 25329 36703
rect 22060 36672 25329 36700
rect 22060 36660 22066 36672
rect 25317 36669 25329 36672
rect 25363 36669 25375 36703
rect 25317 36663 25375 36669
rect 25866 36660 25872 36712
rect 25924 36700 25930 36712
rect 26252 36700 26280 36731
rect 27062 36728 27068 36780
rect 27120 36768 27126 36780
rect 28537 36771 28595 36777
rect 28537 36768 28549 36771
rect 27120 36740 28549 36768
rect 27120 36728 27126 36740
rect 28537 36737 28549 36740
rect 28583 36737 28595 36771
rect 28537 36731 28595 36737
rect 28626 36728 28632 36780
rect 28684 36768 28690 36780
rect 28793 36771 28851 36777
rect 28793 36768 28805 36771
rect 28684 36740 28805 36768
rect 28684 36728 28690 36740
rect 28793 36737 28805 36740
rect 28839 36737 28851 36771
rect 28793 36731 28851 36737
rect 32306 36728 32312 36780
rect 32364 36768 32370 36780
rect 32677 36771 32735 36777
rect 32677 36768 32689 36771
rect 32364 36740 32689 36768
rect 32364 36728 32370 36740
rect 32677 36737 32689 36740
rect 32723 36737 32735 36771
rect 32950 36768 32956 36780
rect 32911 36740 32956 36768
rect 32677 36731 32735 36737
rect 25924 36672 26280 36700
rect 32692 36700 32720 36731
rect 32950 36728 32956 36740
rect 33008 36728 33014 36780
rect 33410 36768 33416 36780
rect 33371 36740 33416 36768
rect 33410 36728 33416 36740
rect 33468 36728 33474 36780
rect 33594 36768 33600 36780
rect 33555 36740 33600 36768
rect 33594 36728 33600 36740
rect 33652 36728 33658 36780
rect 33318 36700 33324 36712
rect 32692 36672 33324 36700
rect 25924 36660 25930 36672
rect 33318 36660 33324 36672
rect 33376 36660 33382 36712
rect 20530 36592 20536 36644
rect 20588 36592 20594 36644
rect 19760 36536 20372 36564
rect 19760 36524 19766 36536
rect 21266 36524 21272 36576
rect 21324 36564 21330 36576
rect 28718 36564 28724 36576
rect 21324 36536 28724 36564
rect 21324 36524 21330 36536
rect 28718 36524 28724 36536
rect 28776 36524 28782 36576
rect 32493 36567 32551 36573
rect 32493 36533 32505 36567
rect 32539 36564 32551 36567
rect 33042 36564 33048 36576
rect 32539 36536 33048 36564
rect 32539 36533 32551 36536
rect 32493 36527 32551 36533
rect 33042 36524 33048 36536
rect 33100 36524 33106 36576
rect 46474 36524 46480 36576
rect 46532 36564 46538 36576
rect 47949 36567 48007 36573
rect 47949 36564 47961 36567
rect 46532 36536 47961 36564
rect 46532 36524 46538 36536
rect 47949 36533 47961 36536
rect 47995 36533 48007 36567
rect 47949 36527 48007 36533
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 16022 36320 16028 36372
rect 16080 36360 16086 36372
rect 16577 36363 16635 36369
rect 16577 36360 16589 36363
rect 16080 36332 16589 36360
rect 16080 36320 16086 36332
rect 16577 36329 16589 36332
rect 16623 36329 16635 36363
rect 20162 36360 20168 36372
rect 20123 36332 20168 36360
rect 16577 36323 16635 36329
rect 20162 36320 20168 36332
rect 20220 36320 20226 36372
rect 25774 36320 25780 36372
rect 25832 36360 25838 36372
rect 26329 36363 26387 36369
rect 26329 36360 26341 36363
rect 25832 36332 26341 36360
rect 25832 36320 25838 36332
rect 26329 36329 26341 36332
rect 26375 36329 26387 36363
rect 26329 36323 26387 36329
rect 28261 36363 28319 36369
rect 28261 36329 28273 36363
rect 28307 36360 28319 36363
rect 28626 36360 28632 36372
rect 28307 36332 28632 36360
rect 28307 36329 28319 36332
rect 28261 36323 28319 36329
rect 24762 36292 24768 36304
rect 24596 36264 24768 36292
rect 15473 36227 15531 36233
rect 15473 36193 15485 36227
rect 15519 36224 15531 36227
rect 16114 36224 16120 36236
rect 15519 36196 16120 36224
rect 15519 36193 15531 36196
rect 15473 36187 15531 36193
rect 16114 36184 16120 36196
rect 16172 36184 16178 36236
rect 16393 36227 16451 36233
rect 16393 36193 16405 36227
rect 16439 36224 16451 36227
rect 16942 36224 16948 36236
rect 16439 36196 16948 36224
rect 16439 36193 16451 36196
rect 16393 36187 16451 36193
rect 16942 36184 16948 36196
rect 17000 36184 17006 36236
rect 18322 36184 18328 36236
rect 18380 36224 18386 36236
rect 20622 36224 20628 36236
rect 18380 36196 20628 36224
rect 18380 36184 18386 36196
rect 20622 36184 20628 36196
rect 20680 36184 20686 36236
rect 11790 36116 11796 36168
rect 11848 36156 11854 36168
rect 12342 36156 12348 36168
rect 11848 36128 12348 36156
rect 11848 36116 11854 36128
rect 12342 36116 12348 36128
rect 12400 36116 12406 36168
rect 15194 36156 15200 36168
rect 15155 36128 15200 36156
rect 15194 36116 15200 36128
rect 15252 36116 15258 36168
rect 16298 36156 16304 36168
rect 16259 36128 16304 36156
rect 16298 36116 16304 36128
rect 16356 36116 16362 36168
rect 19429 36159 19487 36165
rect 19429 36125 19441 36159
rect 19475 36125 19487 36159
rect 19429 36119 19487 36125
rect 19613 36159 19671 36165
rect 19613 36125 19625 36159
rect 19659 36156 19671 36159
rect 20162 36156 20168 36168
rect 19659 36128 20168 36156
rect 19659 36125 19671 36128
rect 19613 36119 19671 36125
rect 12612 36091 12670 36097
rect 12612 36057 12624 36091
rect 12658 36088 12670 36091
rect 12802 36088 12808 36100
rect 12658 36060 12808 36088
rect 12658 36057 12670 36060
rect 12612 36051 12670 36057
rect 12802 36048 12808 36060
rect 12860 36048 12866 36100
rect 19444 36088 19472 36119
rect 20162 36116 20168 36128
rect 20220 36116 20226 36168
rect 20346 36156 20352 36168
rect 20307 36128 20352 36156
rect 20346 36116 20352 36128
rect 20404 36116 20410 36168
rect 20530 36156 20536 36168
rect 20491 36128 20536 36156
rect 20530 36116 20536 36128
rect 20588 36116 20594 36168
rect 22186 36156 22192 36168
rect 22147 36128 22192 36156
rect 22186 36116 22192 36128
rect 22244 36116 22250 36168
rect 22373 36159 22431 36165
rect 22373 36125 22385 36159
rect 22419 36156 22431 36159
rect 22646 36156 22652 36168
rect 22419 36128 22652 36156
rect 22419 36125 22431 36128
rect 22373 36119 22431 36125
rect 22646 36116 22652 36128
rect 22704 36116 22710 36168
rect 24596 36165 24624 36264
rect 24762 36252 24768 36264
rect 24820 36252 24826 36304
rect 24673 36227 24731 36233
rect 24673 36193 24685 36227
rect 24719 36224 24731 36227
rect 25409 36227 25467 36233
rect 25409 36224 25421 36227
rect 24719 36196 25421 36224
rect 24719 36193 24731 36196
rect 24673 36187 24731 36193
rect 25409 36193 25421 36196
rect 25455 36193 25467 36227
rect 25409 36187 25467 36193
rect 25501 36227 25559 36233
rect 25501 36193 25513 36227
rect 25547 36224 25559 36227
rect 25866 36224 25872 36236
rect 25547 36196 25872 36224
rect 25547 36193 25559 36196
rect 25501 36187 25559 36193
rect 25866 36184 25872 36196
rect 25924 36184 25930 36236
rect 26344 36224 26372 36323
rect 28626 36320 28632 36332
rect 28684 36320 28690 36372
rect 32309 36363 32367 36369
rect 32309 36329 32321 36363
rect 32355 36360 32367 36363
rect 32674 36360 32680 36372
rect 32355 36332 32680 36360
rect 32355 36329 32367 36332
rect 32309 36323 32367 36329
rect 32674 36320 32680 36332
rect 32732 36320 32738 36372
rect 33318 36320 33324 36372
rect 33376 36360 33382 36372
rect 33965 36363 34023 36369
rect 33965 36360 33977 36363
rect 33376 36332 33977 36360
rect 33376 36320 33382 36332
rect 33965 36329 33977 36332
rect 34011 36329 34023 36363
rect 33965 36323 34023 36329
rect 33134 36252 33140 36304
rect 33192 36292 33198 36304
rect 34422 36292 34428 36304
rect 33192 36264 34428 36292
rect 33192 36252 33198 36264
rect 34422 36252 34428 36264
rect 34480 36252 34486 36304
rect 26344 36196 27108 36224
rect 24581 36159 24639 36165
rect 24581 36125 24593 36159
rect 24627 36125 24639 36159
rect 24581 36119 24639 36125
rect 24765 36159 24823 36165
rect 24765 36125 24777 36159
rect 24811 36156 24823 36159
rect 25038 36156 25044 36168
rect 24811 36128 25044 36156
rect 24811 36125 24823 36128
rect 24765 36119 24823 36125
rect 25038 36116 25044 36128
rect 25096 36156 25102 36168
rect 25593 36159 25651 36165
rect 25096 36128 25544 36156
rect 25096 36116 25102 36128
rect 19702 36088 19708 36100
rect 19444 36060 19708 36088
rect 19702 36048 19708 36060
rect 19760 36088 19766 36100
rect 20070 36088 20076 36100
rect 19760 36060 20076 36088
rect 19760 36048 19766 36060
rect 20070 36048 20076 36060
rect 20128 36048 20134 36100
rect 22278 36048 22284 36100
rect 22336 36088 22342 36100
rect 22830 36088 22836 36100
rect 22336 36060 22836 36088
rect 22336 36048 22342 36060
rect 22830 36048 22836 36060
rect 22888 36048 22894 36100
rect 13725 36023 13783 36029
rect 13725 35989 13737 36023
rect 13771 36020 13783 36023
rect 13814 36020 13820 36032
rect 13771 35992 13820 36020
rect 13771 35989 13783 35992
rect 13725 35983 13783 35989
rect 13814 35980 13820 35992
rect 13872 35980 13878 36032
rect 14826 36020 14832 36032
rect 14787 35992 14832 36020
rect 14826 35980 14832 35992
rect 14884 35980 14890 36032
rect 15286 35980 15292 36032
rect 15344 36020 15350 36032
rect 15344 35992 15389 36020
rect 15344 35980 15350 35992
rect 19334 35980 19340 36032
rect 19392 36020 19398 36032
rect 19521 36023 19579 36029
rect 19521 36020 19533 36023
rect 19392 35992 19533 36020
rect 19392 35980 19398 35992
rect 19521 35989 19533 35992
rect 19567 35989 19579 36023
rect 19521 35983 19579 35989
rect 22373 36023 22431 36029
rect 22373 35989 22385 36023
rect 22419 36020 22431 36023
rect 22738 36020 22744 36032
rect 22419 35992 22744 36020
rect 22419 35989 22431 35992
rect 22373 35983 22431 35989
rect 22738 35980 22744 35992
rect 22796 35980 22802 36032
rect 25222 36020 25228 36032
rect 25183 35992 25228 36020
rect 25222 35980 25228 35992
rect 25280 35980 25286 36032
rect 25516 36020 25544 36128
rect 25593 36125 25605 36159
rect 25639 36125 25651 36159
rect 25593 36119 25651 36125
rect 25608 36088 25636 36119
rect 25682 36116 25688 36168
rect 25740 36156 25746 36168
rect 26237 36159 26295 36165
rect 25740 36128 25785 36156
rect 25740 36116 25746 36128
rect 26237 36125 26249 36159
rect 26283 36156 26295 36159
rect 26326 36156 26332 36168
rect 26283 36128 26332 36156
rect 26283 36125 26295 36128
rect 26237 36119 26295 36125
rect 26326 36116 26332 36128
rect 26384 36116 26390 36168
rect 26418 36116 26424 36168
rect 26476 36156 26482 36168
rect 26878 36156 26884 36168
rect 26476 36128 26521 36156
rect 26839 36128 26884 36156
rect 26476 36116 26482 36128
rect 26878 36116 26884 36128
rect 26936 36116 26942 36168
rect 27080 36165 27108 36196
rect 32674 36184 32680 36236
rect 32732 36224 32738 36236
rect 33413 36227 33471 36233
rect 33413 36224 33425 36227
rect 32732 36196 33425 36224
rect 32732 36184 32738 36196
rect 33413 36193 33425 36196
rect 33459 36193 33471 36227
rect 46474 36224 46480 36236
rect 46435 36196 46480 36224
rect 33413 36187 33471 36193
rect 46474 36184 46480 36196
rect 46532 36184 46538 36236
rect 48222 36224 48228 36236
rect 48183 36196 48228 36224
rect 48222 36184 48228 36196
rect 48280 36184 48286 36236
rect 27065 36159 27123 36165
rect 27065 36125 27077 36159
rect 27111 36125 27123 36159
rect 27065 36119 27123 36125
rect 28258 36116 28264 36168
rect 28316 36156 28322 36168
rect 28445 36159 28503 36165
rect 28445 36156 28457 36159
rect 28316 36128 28457 36156
rect 28316 36116 28322 36128
rect 28445 36125 28457 36128
rect 28491 36125 28503 36159
rect 28445 36119 28503 36125
rect 28721 36159 28779 36165
rect 28721 36125 28733 36159
rect 28767 36125 28779 36159
rect 28721 36119 28779 36125
rect 26694 36088 26700 36100
rect 25608 36060 26700 36088
rect 26694 36048 26700 36060
rect 26752 36048 26758 36100
rect 27614 36048 27620 36100
rect 27672 36088 27678 36100
rect 28736 36088 28764 36119
rect 30282 36116 30288 36168
rect 30340 36156 30346 36168
rect 30929 36159 30987 36165
rect 30929 36156 30941 36159
rect 30340 36128 30941 36156
rect 30340 36116 30346 36128
rect 30929 36125 30941 36128
rect 30975 36125 30987 36159
rect 30929 36119 30987 36125
rect 32953 36159 33011 36165
rect 32953 36125 32965 36159
rect 32999 36125 33011 36159
rect 32953 36119 33011 36125
rect 27672 36060 28764 36088
rect 31196 36091 31254 36097
rect 27672 36048 27678 36060
rect 31196 36057 31208 36091
rect 31242 36088 31254 36091
rect 32769 36091 32827 36097
rect 32769 36088 32781 36091
rect 31242 36060 32781 36088
rect 31242 36057 31254 36060
rect 31196 36051 31254 36057
rect 32769 36057 32781 36060
rect 32815 36057 32827 36091
rect 32769 36051 32827 36057
rect 26973 36023 27031 36029
rect 26973 36020 26985 36023
rect 25516 35992 26985 36020
rect 26973 35989 26985 35992
rect 27019 35989 27031 36023
rect 26973 35983 27031 35989
rect 28442 35980 28448 36032
rect 28500 36020 28506 36032
rect 28629 36023 28687 36029
rect 28629 36020 28641 36023
rect 28500 35992 28641 36020
rect 28500 35980 28506 35992
rect 28629 35989 28641 35992
rect 28675 35989 28687 36023
rect 32968 36020 32996 36119
rect 33042 36116 33048 36168
rect 33100 36156 33106 36168
rect 33870 36156 33876 36168
rect 33100 36128 33145 36156
rect 33831 36128 33876 36156
rect 33100 36116 33106 36128
rect 33870 36116 33876 36128
rect 33928 36116 33934 36168
rect 33134 36088 33140 36100
rect 33095 36060 33140 36088
rect 33134 36048 33140 36060
rect 33192 36048 33198 36100
rect 33226 36048 33232 36100
rect 33284 36097 33290 36100
rect 33284 36091 33313 36097
rect 33301 36057 33313 36091
rect 33284 36051 33313 36057
rect 46661 36091 46719 36097
rect 46661 36057 46673 36091
rect 46707 36088 46719 36091
rect 47854 36088 47860 36100
rect 46707 36060 47860 36088
rect 46707 36057 46719 36060
rect 46661 36051 46719 36057
rect 33284 36048 33290 36051
rect 47854 36048 47860 36060
rect 47912 36048 47918 36100
rect 33410 36020 33416 36032
rect 32968 35992 33416 36020
rect 28629 35983 28687 35989
rect 33410 35980 33416 35992
rect 33468 35980 33474 36032
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 12802 35816 12808 35828
rect 12763 35788 12808 35816
rect 12802 35776 12808 35788
rect 12860 35776 12866 35828
rect 13814 35816 13820 35828
rect 13775 35788 13820 35816
rect 13814 35776 13820 35788
rect 13872 35776 13878 35828
rect 13909 35819 13967 35825
rect 13909 35785 13921 35819
rect 13955 35816 13967 35819
rect 14826 35816 14832 35828
rect 13955 35788 14832 35816
rect 13955 35785 13967 35788
rect 13909 35779 13967 35785
rect 14826 35776 14832 35788
rect 14884 35776 14890 35828
rect 16942 35816 16948 35828
rect 16903 35788 16948 35816
rect 16942 35776 16948 35788
rect 17000 35776 17006 35828
rect 18785 35819 18843 35825
rect 18785 35785 18797 35819
rect 18831 35816 18843 35819
rect 19978 35816 19984 35828
rect 18831 35788 19984 35816
rect 18831 35785 18843 35788
rect 18785 35779 18843 35785
rect 19978 35776 19984 35788
rect 20036 35776 20042 35828
rect 22186 35776 22192 35828
rect 22244 35816 22250 35828
rect 23290 35816 23296 35828
rect 22244 35788 23296 35816
rect 22244 35776 22250 35788
rect 23290 35776 23296 35788
rect 23348 35816 23354 35828
rect 23385 35819 23443 35825
rect 23385 35816 23397 35819
rect 23348 35788 23397 35816
rect 23348 35776 23354 35788
rect 23385 35785 23397 35788
rect 23431 35785 23443 35819
rect 23385 35779 23443 35785
rect 25133 35819 25191 35825
rect 25133 35785 25145 35819
rect 25179 35816 25191 35819
rect 25222 35816 25228 35828
rect 25179 35788 25228 35816
rect 25179 35785 25191 35788
rect 25133 35779 25191 35785
rect 25222 35776 25228 35788
rect 25280 35776 25286 35828
rect 26237 35819 26295 35825
rect 26237 35785 26249 35819
rect 26283 35816 26295 35819
rect 26878 35816 26884 35828
rect 26283 35788 26884 35816
rect 26283 35785 26295 35788
rect 26237 35779 26295 35785
rect 26878 35776 26884 35788
rect 26936 35776 26942 35828
rect 30098 35776 30104 35828
rect 30156 35816 30162 35828
rect 30926 35816 30932 35828
rect 30156 35788 30932 35816
rect 30156 35776 30162 35788
rect 30926 35776 30932 35788
rect 30984 35816 30990 35828
rect 33134 35816 33140 35828
rect 30984 35788 33140 35816
rect 30984 35776 30990 35788
rect 33134 35776 33140 35788
rect 33192 35776 33198 35828
rect 33410 35816 33416 35828
rect 33371 35788 33416 35816
rect 33410 35776 33416 35788
rect 33468 35776 33474 35828
rect 47854 35816 47860 35828
rect 47815 35788 47860 35816
rect 47854 35776 47860 35788
rect 47912 35776 47918 35828
rect 13630 35708 13636 35760
rect 13688 35748 13694 35760
rect 14645 35751 14703 35757
rect 14645 35748 14657 35751
rect 13688 35720 14657 35748
rect 13688 35708 13694 35720
rect 14645 35717 14657 35720
rect 14691 35717 14703 35751
rect 14645 35711 14703 35717
rect 15378 35708 15384 35760
rect 15436 35748 15442 35760
rect 15657 35751 15715 35757
rect 15657 35748 15669 35751
rect 15436 35720 15669 35748
rect 15436 35708 15442 35720
rect 15657 35717 15669 35720
rect 15703 35748 15715 35751
rect 19334 35748 19340 35760
rect 15703 35720 17080 35748
rect 15703 35717 15715 35720
rect 15657 35711 15715 35717
rect 12989 35683 13047 35689
rect 12989 35649 13001 35683
rect 13035 35680 13047 35683
rect 13035 35652 13492 35680
rect 13035 35649 13047 35652
rect 12989 35643 13047 35649
rect 13464 35553 13492 35652
rect 13722 35640 13728 35692
rect 13780 35680 13786 35692
rect 17052 35689 17080 35720
rect 17696 35720 19340 35748
rect 17696 35692 17724 35720
rect 14829 35683 14887 35689
rect 14829 35680 14841 35683
rect 13780 35652 14841 35680
rect 13780 35640 13786 35652
rect 14829 35649 14841 35652
rect 14875 35649 14887 35683
rect 14829 35643 14887 35649
rect 15013 35683 15071 35689
rect 15013 35649 15025 35683
rect 15059 35680 15071 35683
rect 16117 35683 16175 35689
rect 16117 35680 16129 35683
rect 15059 35652 16129 35680
rect 15059 35649 15071 35652
rect 15013 35643 15071 35649
rect 16117 35649 16129 35652
rect 16163 35680 16175 35683
rect 16853 35683 16911 35689
rect 16853 35680 16865 35683
rect 16163 35652 16865 35680
rect 16163 35649 16175 35652
rect 16117 35643 16175 35649
rect 16853 35649 16865 35652
rect 16899 35649 16911 35683
rect 16853 35643 16911 35649
rect 17037 35683 17095 35689
rect 17037 35649 17049 35683
rect 17083 35649 17095 35683
rect 17678 35680 17684 35692
rect 17639 35652 17684 35680
rect 17037 35643 17095 35649
rect 17678 35640 17684 35652
rect 17736 35640 17742 35692
rect 17862 35680 17868 35692
rect 17823 35652 17868 35680
rect 17862 35640 17868 35652
rect 17920 35640 17926 35692
rect 18984 35689 19012 35720
rect 19334 35708 19340 35720
rect 19392 35708 19398 35760
rect 25041 35751 25099 35757
rect 25041 35717 25053 35751
rect 25087 35748 25099 35751
rect 25869 35751 25927 35757
rect 25869 35748 25881 35751
rect 25087 35720 25881 35748
rect 25087 35717 25099 35720
rect 25041 35711 25099 35717
rect 25869 35717 25881 35720
rect 25915 35748 25927 35751
rect 26326 35748 26332 35760
rect 25915 35720 26332 35748
rect 25915 35717 25927 35720
rect 25869 35711 25927 35717
rect 26326 35708 26332 35720
rect 26384 35708 26390 35760
rect 30282 35748 30288 35760
rect 28368 35720 30288 35748
rect 17957 35683 18015 35689
rect 17957 35649 17969 35683
rect 18003 35649 18015 35683
rect 17957 35643 18015 35649
rect 18969 35683 19027 35689
rect 18969 35649 18981 35683
rect 19015 35649 19027 35683
rect 18969 35643 19027 35649
rect 14090 35612 14096 35624
rect 14051 35584 14096 35612
rect 14090 35572 14096 35584
rect 14148 35572 14154 35624
rect 16025 35615 16083 35621
rect 16025 35581 16037 35615
rect 16071 35612 16083 35615
rect 16298 35612 16304 35624
rect 16071 35584 16304 35612
rect 16071 35581 16083 35584
rect 16025 35575 16083 35581
rect 16298 35572 16304 35584
rect 16356 35612 16362 35624
rect 16356 35584 17724 35612
rect 16356 35572 16362 35584
rect 17696 35553 17724 35584
rect 13449 35547 13507 35553
rect 13449 35513 13461 35547
rect 13495 35513 13507 35547
rect 13449 35507 13507 35513
rect 17681 35547 17739 35553
rect 17681 35513 17693 35547
rect 17727 35513 17739 35547
rect 17972 35544 18000 35643
rect 19058 35640 19064 35692
rect 19116 35680 19122 35692
rect 19242 35680 19248 35692
rect 19116 35652 19161 35680
rect 19203 35652 19248 35680
rect 19116 35640 19122 35652
rect 19242 35640 19248 35652
rect 19300 35640 19306 35692
rect 19429 35683 19487 35689
rect 19429 35649 19441 35683
rect 19475 35680 19487 35683
rect 19610 35680 19616 35692
rect 19475 35652 19616 35680
rect 19475 35649 19487 35652
rect 19429 35643 19487 35649
rect 19610 35640 19616 35652
rect 19668 35640 19674 35692
rect 20070 35680 20076 35692
rect 20031 35652 20076 35680
rect 20070 35640 20076 35652
rect 20128 35640 20134 35692
rect 22094 35640 22100 35692
rect 22152 35680 22158 35692
rect 22261 35683 22319 35689
rect 22261 35680 22273 35683
rect 22152 35652 22273 35680
rect 22152 35640 22158 35652
rect 22261 35649 22273 35652
rect 22307 35649 22319 35683
rect 22261 35643 22319 35649
rect 26053 35683 26111 35689
rect 26053 35649 26065 35683
rect 26099 35680 26111 35683
rect 26418 35680 26424 35692
rect 26099 35652 26424 35680
rect 26099 35649 26111 35652
rect 26053 35643 26111 35649
rect 26418 35640 26424 35652
rect 26476 35680 26482 35692
rect 27430 35680 27436 35692
rect 26476 35652 27436 35680
rect 26476 35640 26482 35652
rect 27430 35640 27436 35652
rect 27488 35640 27494 35692
rect 28368 35689 28396 35720
rect 30282 35708 30288 35720
rect 30340 35708 30346 35760
rect 30466 35748 30472 35760
rect 30427 35720 30472 35748
rect 30466 35708 30472 35720
rect 30524 35708 30530 35760
rect 32950 35708 32956 35760
rect 33008 35748 33014 35760
rect 33505 35751 33563 35757
rect 33505 35748 33517 35751
rect 33008 35720 33517 35748
rect 33008 35708 33014 35720
rect 33505 35717 33517 35720
rect 33551 35717 33563 35751
rect 33505 35711 33563 35717
rect 28353 35683 28411 35689
rect 28353 35649 28365 35683
rect 28399 35649 28411 35683
rect 28353 35643 28411 35649
rect 28620 35683 28678 35689
rect 28620 35649 28632 35683
rect 28666 35680 28678 35683
rect 28994 35680 29000 35692
rect 28666 35652 29000 35680
rect 28666 35649 28678 35652
rect 28620 35643 28678 35649
rect 28994 35640 29000 35652
rect 29052 35640 29058 35692
rect 30098 35640 30104 35692
rect 30156 35680 30162 35692
rect 30193 35683 30251 35689
rect 30193 35680 30205 35683
rect 30156 35652 30205 35680
rect 30156 35640 30162 35652
rect 30193 35649 30205 35652
rect 30239 35649 30251 35683
rect 30193 35643 30251 35649
rect 31662 35640 31668 35692
rect 31720 35680 31726 35692
rect 32493 35683 32551 35689
rect 32493 35680 32505 35683
rect 31720 35652 32505 35680
rect 31720 35640 31726 35652
rect 32493 35649 32505 35652
rect 32539 35649 32551 35683
rect 33318 35680 33324 35692
rect 33279 35652 33324 35680
rect 32493 35643 32551 35649
rect 33318 35640 33324 35652
rect 33376 35640 33382 35692
rect 33597 35683 33655 35689
rect 33597 35649 33609 35683
rect 33643 35680 33655 35683
rect 33686 35680 33692 35692
rect 33643 35652 33692 35680
rect 33643 35649 33655 35652
rect 33597 35643 33655 35649
rect 33686 35640 33692 35652
rect 33744 35640 33750 35692
rect 47394 35640 47400 35692
rect 47452 35680 47458 35692
rect 47765 35683 47823 35689
rect 47765 35680 47777 35683
rect 47452 35652 47777 35680
rect 47452 35640 47458 35652
rect 47765 35649 47777 35652
rect 47811 35649 47823 35683
rect 47765 35643 47823 35649
rect 18874 35572 18880 35624
rect 18932 35612 18938 35624
rect 19889 35615 19947 35621
rect 19889 35612 19901 35615
rect 18932 35584 19901 35612
rect 18932 35572 18938 35584
rect 19889 35581 19901 35584
rect 19935 35612 19947 35615
rect 20162 35612 20168 35624
rect 19935 35584 20168 35612
rect 19935 35581 19947 35584
rect 19889 35575 19947 35581
rect 20162 35572 20168 35584
rect 20220 35572 20226 35624
rect 22002 35612 22008 35624
rect 21963 35584 22008 35612
rect 22002 35572 22008 35584
rect 22060 35572 22066 35624
rect 25317 35615 25375 35621
rect 25317 35581 25329 35615
rect 25363 35612 25375 35615
rect 25406 35612 25412 35624
rect 25363 35584 25412 35612
rect 25363 35581 25375 35584
rect 25317 35575 25375 35581
rect 25406 35572 25412 35584
rect 25464 35572 25470 35624
rect 32585 35615 32643 35621
rect 32585 35581 32597 35615
rect 32631 35612 32643 35615
rect 32674 35612 32680 35624
rect 32631 35584 32680 35612
rect 32631 35581 32643 35584
rect 32585 35575 32643 35581
rect 32674 35572 32680 35584
rect 32732 35572 32738 35624
rect 32861 35615 32919 35621
rect 32861 35581 32873 35615
rect 32907 35612 32919 35615
rect 33870 35612 33876 35624
rect 32907 35584 33876 35612
rect 32907 35581 32919 35584
rect 32861 35575 32919 35581
rect 33870 35572 33876 35584
rect 33928 35572 33934 35624
rect 19153 35547 19211 35553
rect 19153 35544 19165 35547
rect 17972 35516 19165 35544
rect 17681 35507 17739 35513
rect 19153 35513 19165 35516
rect 19199 35544 19211 35547
rect 19794 35544 19800 35556
rect 19199 35516 19800 35544
rect 19199 35513 19211 35516
rect 19153 35507 19211 35513
rect 19794 35504 19800 35516
rect 19852 35504 19858 35556
rect 30466 35504 30472 35556
rect 30524 35544 30530 35556
rect 31662 35544 31668 35556
rect 30524 35516 31668 35544
rect 30524 35504 30530 35516
rect 31662 35504 31668 35516
rect 31720 35544 31726 35556
rect 33226 35544 33232 35556
rect 31720 35516 33232 35544
rect 31720 35504 31726 35516
rect 33226 35504 33232 35516
rect 33284 35504 33290 35556
rect 15654 35436 15660 35488
rect 15712 35476 15718 35488
rect 16301 35479 16359 35485
rect 16301 35476 16313 35479
rect 15712 35448 16313 35476
rect 15712 35436 15718 35448
rect 16301 35445 16313 35448
rect 16347 35445 16359 35479
rect 16301 35439 16359 35445
rect 19518 35436 19524 35488
rect 19576 35476 19582 35488
rect 20257 35479 20315 35485
rect 20257 35476 20269 35479
rect 19576 35448 20269 35476
rect 19576 35436 19582 35448
rect 20257 35445 20269 35448
rect 20303 35445 20315 35479
rect 20257 35439 20315 35445
rect 20898 35436 20904 35488
rect 20956 35476 20962 35488
rect 22646 35476 22652 35488
rect 20956 35448 22652 35476
rect 20956 35436 20962 35448
rect 22646 35436 22652 35448
rect 22704 35436 22710 35488
rect 24578 35436 24584 35488
rect 24636 35476 24642 35488
rect 24673 35479 24731 35485
rect 24673 35476 24685 35479
rect 24636 35448 24685 35476
rect 24636 35436 24642 35448
rect 24673 35445 24685 35448
rect 24719 35445 24731 35479
rect 24673 35439 24731 35445
rect 29733 35479 29791 35485
rect 29733 35445 29745 35479
rect 29779 35476 29791 35479
rect 30190 35476 30196 35488
rect 29779 35448 30196 35476
rect 29779 35445 29791 35448
rect 29733 35439 29791 35445
rect 30190 35436 30196 35448
rect 30248 35436 30254 35488
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 15286 35232 15292 35284
rect 15344 35272 15350 35284
rect 15841 35275 15899 35281
rect 15841 35272 15853 35275
rect 15344 35244 15853 35272
rect 15344 35232 15350 35244
rect 15841 35241 15853 35244
rect 15887 35241 15899 35275
rect 15841 35235 15899 35241
rect 16942 35232 16948 35284
rect 17000 35272 17006 35284
rect 17405 35275 17463 35281
rect 17405 35272 17417 35275
rect 17000 35244 17417 35272
rect 17000 35232 17006 35244
rect 17405 35241 17417 35244
rect 17451 35241 17463 35275
rect 19610 35272 19616 35284
rect 19571 35244 19616 35272
rect 17405 35235 17463 35241
rect 19610 35232 19616 35244
rect 19668 35232 19674 35284
rect 22649 35275 22707 35281
rect 22649 35241 22661 35275
rect 22695 35272 22707 35275
rect 23382 35272 23388 35284
rect 22695 35244 23388 35272
rect 22695 35241 22707 35244
rect 22649 35235 22707 35241
rect 23382 35232 23388 35244
rect 23440 35232 23446 35284
rect 25961 35275 26019 35281
rect 24596 35244 25544 35272
rect 13633 35207 13691 35213
rect 13633 35173 13645 35207
rect 13679 35204 13691 35207
rect 15378 35204 15384 35216
rect 13679 35176 15384 35204
rect 13679 35173 13691 35176
rect 13633 35167 13691 35173
rect 15378 35164 15384 35176
rect 15436 35164 15442 35216
rect 17313 35207 17371 35213
rect 17313 35173 17325 35207
rect 17359 35204 17371 35207
rect 17678 35204 17684 35216
rect 17359 35176 17684 35204
rect 17359 35173 17371 35176
rect 17313 35167 17371 35173
rect 17678 35164 17684 35176
rect 17736 35164 17742 35216
rect 19058 35164 19064 35216
rect 19116 35204 19122 35216
rect 19518 35204 19524 35216
rect 19116 35176 19524 35204
rect 19116 35164 19122 35176
rect 19518 35164 19524 35176
rect 19576 35164 19582 35216
rect 19794 35164 19800 35216
rect 19852 35204 19858 35216
rect 24596 35204 24624 35244
rect 19852 35176 24624 35204
rect 25516 35204 25544 35244
rect 25961 35241 25973 35275
rect 26007 35272 26019 35275
rect 26326 35272 26332 35284
rect 26007 35244 26332 35272
rect 26007 35241 26019 35244
rect 25961 35235 26019 35241
rect 26326 35232 26332 35244
rect 26384 35232 26390 35284
rect 27890 35204 27896 35216
rect 25516 35176 27896 35204
rect 19852 35164 19858 35176
rect 27890 35164 27896 35176
rect 27948 35164 27954 35216
rect 13814 35096 13820 35148
rect 13872 35136 13878 35148
rect 15654 35136 15660 35148
rect 13872 35108 14596 35136
rect 15615 35108 15660 35136
rect 13872 35096 13878 35108
rect 14568 35080 14596 35108
rect 15654 35096 15660 35108
rect 15712 35096 15718 35148
rect 19705 35139 19763 35145
rect 19705 35136 19717 35139
rect 17696 35108 19717 35136
rect 13541 35071 13599 35077
rect 13541 35037 13553 35071
rect 13587 35068 13599 35071
rect 13630 35068 13636 35080
rect 13587 35040 13636 35068
rect 13587 35037 13599 35040
rect 13541 35031 13599 35037
rect 13630 35028 13636 35040
rect 13688 35028 13694 35080
rect 13722 35028 13728 35080
rect 13780 35068 13786 35080
rect 14550 35068 14556 35080
rect 13780 35040 13825 35068
rect 14463 35040 14556 35068
rect 13780 35028 13786 35040
rect 14550 35028 14556 35040
rect 14608 35028 14614 35080
rect 14734 35068 14740 35080
rect 14695 35040 14740 35068
rect 14734 35028 14740 35040
rect 14792 35028 14798 35080
rect 15565 35071 15623 35077
rect 15565 35037 15577 35071
rect 15611 35068 15623 35071
rect 15838 35068 15844 35080
rect 15611 35040 15844 35068
rect 15611 35037 15623 35040
rect 15565 35031 15623 35037
rect 15838 35028 15844 35040
rect 15896 35068 15902 35080
rect 17696 35077 17724 35108
rect 19705 35105 19717 35108
rect 19751 35136 19763 35139
rect 19812 35136 19840 35164
rect 21634 35136 21640 35148
rect 19751 35108 19840 35136
rect 21595 35108 21640 35136
rect 19751 35105 19763 35108
rect 19705 35099 19763 35105
rect 21634 35096 21640 35108
rect 21692 35096 21698 35148
rect 22370 35096 22376 35148
rect 22428 35096 22434 35148
rect 27341 35139 27399 35145
rect 27341 35105 27353 35139
rect 27387 35136 27399 35139
rect 27522 35136 27528 35148
rect 27387 35108 27528 35136
rect 27387 35105 27399 35108
rect 27341 35099 27399 35105
rect 27522 35096 27528 35108
rect 27580 35096 27586 35148
rect 17221 35071 17279 35077
rect 17221 35068 17233 35071
rect 15896 35040 17233 35068
rect 15896 35028 15902 35040
rect 17221 35037 17233 35040
rect 17267 35037 17279 35071
rect 17221 35031 17279 35037
rect 17681 35071 17739 35077
rect 17681 35037 17693 35071
rect 17727 35037 17739 35071
rect 17681 35031 17739 35037
rect 18509 35071 18567 35077
rect 18509 35037 18521 35071
rect 18555 35037 18567 35071
rect 18509 35031 18567 35037
rect 18693 35071 18751 35077
rect 18693 35037 18705 35071
rect 18739 35068 18751 35071
rect 18874 35068 18880 35080
rect 18739 35040 18880 35068
rect 18739 35037 18751 35040
rect 18693 35031 18751 35037
rect 18524 35000 18552 35031
rect 18874 35028 18880 35040
rect 18932 35028 18938 35080
rect 19334 35028 19340 35080
rect 19392 35068 19398 35080
rect 19429 35071 19487 35077
rect 19429 35068 19441 35071
rect 19392 35040 19441 35068
rect 19392 35028 19398 35040
rect 19429 35037 19441 35040
rect 19475 35037 19487 35071
rect 19429 35031 19487 35037
rect 21726 35028 21732 35080
rect 21784 35077 21790 35080
rect 21784 35068 21792 35077
rect 22278 35068 22284 35080
rect 21784 35040 21829 35068
rect 22239 35040 22284 35068
rect 21784 35031 21792 35040
rect 21784 35028 21790 35031
rect 22278 35028 22284 35040
rect 22336 35028 22342 35080
rect 22388 35068 22416 35096
rect 22557 35071 22615 35077
rect 22557 35068 22569 35071
rect 22388 35040 22569 35068
rect 22557 35037 22569 35040
rect 22603 35037 22615 35071
rect 22557 35031 22615 35037
rect 22646 35028 22652 35080
rect 22704 35068 22710 35080
rect 23477 35071 23535 35077
rect 23477 35068 23489 35071
rect 22704 35040 23489 35068
rect 22704 35028 22710 35040
rect 23477 35037 23489 35040
rect 23523 35037 23535 35071
rect 23477 35031 23535 35037
rect 24581 35071 24639 35077
rect 24581 35037 24593 35071
rect 24627 35068 24639 35071
rect 27062 35068 27068 35080
rect 24627 35040 27068 35068
rect 24627 35037 24639 35040
rect 24581 35031 24639 35037
rect 27062 35028 27068 35040
rect 27120 35028 27126 35080
rect 27154 35028 27160 35080
rect 27212 35068 27218 35080
rect 27433 35071 27491 35077
rect 27212 35040 27257 35068
rect 27212 35028 27218 35040
rect 27433 35037 27445 35071
rect 27479 35037 27491 35071
rect 28718 35068 28724 35080
rect 28679 35040 28724 35068
rect 27433 35031 27491 35037
rect 20070 35000 20076 35012
rect 18524 34972 20076 35000
rect 20070 34960 20076 34972
rect 20128 34960 20134 35012
rect 21361 35003 21419 35009
rect 21361 34969 21373 35003
rect 21407 34969 21419 35003
rect 21361 34963 21419 34969
rect 14645 34935 14703 34941
rect 14645 34901 14657 34935
rect 14691 34932 14703 34935
rect 15010 34932 15016 34944
rect 14691 34904 15016 34932
rect 14691 34901 14703 34904
rect 14645 34895 14703 34901
rect 15010 34892 15016 34904
rect 15068 34892 15074 34944
rect 16666 34892 16672 34944
rect 16724 34932 16730 34944
rect 16945 34935 17003 34941
rect 16945 34932 16957 34935
rect 16724 34904 16957 34932
rect 16724 34892 16730 34904
rect 16945 34901 16957 34904
rect 16991 34901 17003 34935
rect 16945 34895 17003 34901
rect 17589 34935 17647 34941
rect 17589 34901 17601 34935
rect 17635 34932 17647 34935
rect 17862 34932 17868 34944
rect 17635 34904 17868 34932
rect 17635 34901 17647 34904
rect 17589 34895 17647 34901
rect 17862 34892 17868 34904
rect 17920 34932 17926 34944
rect 18601 34935 18659 34941
rect 18601 34932 18613 34935
rect 17920 34904 18613 34932
rect 17920 34892 17926 34904
rect 18601 34901 18613 34904
rect 18647 34901 18659 34935
rect 21376 34932 21404 34963
rect 21450 34960 21456 35012
rect 21508 35000 21514 35012
rect 21545 35003 21603 35009
rect 21545 35000 21557 35003
rect 21508 34972 21557 35000
rect 21508 34960 21514 34972
rect 21545 34969 21557 34972
rect 21591 34969 21603 35003
rect 21545 34963 21603 34969
rect 21637 35003 21695 35009
rect 21637 34969 21649 35003
rect 21683 35000 21695 35003
rect 21910 35000 21916 35012
rect 21683 34972 21916 35000
rect 21683 34969 21695 34972
rect 21637 34963 21695 34969
rect 21910 34960 21916 34972
rect 21968 34960 21974 35012
rect 22296 35000 22324 35028
rect 23106 35000 23112 35012
rect 22296 34972 23112 35000
rect 23106 34960 23112 34972
rect 23164 34960 23170 35012
rect 23290 35000 23296 35012
rect 23251 34972 23296 35000
rect 23290 34960 23296 34972
rect 23348 34960 23354 35012
rect 24394 34960 24400 35012
rect 24452 35000 24458 35012
rect 24826 35003 24884 35009
rect 24826 35000 24838 35003
rect 24452 34972 24838 35000
rect 24452 34960 24458 34972
rect 24826 34969 24838 34972
rect 24872 34969 24884 35003
rect 24826 34963 24884 34969
rect 26418 34960 26424 35012
rect 26476 35000 26482 35012
rect 27448 35000 27476 35031
rect 28718 35028 28724 35040
rect 28776 35028 28782 35080
rect 28997 35071 29055 35077
rect 28997 35037 29009 35071
rect 29043 35068 29055 35071
rect 29086 35068 29092 35080
rect 29043 35040 29092 35068
rect 29043 35037 29055 35040
rect 28997 35031 29055 35037
rect 29086 35028 29092 35040
rect 29144 35028 29150 35080
rect 29181 35071 29239 35077
rect 29181 35037 29193 35071
rect 29227 35068 29239 35071
rect 30190 35068 30196 35080
rect 29227 35040 30196 35068
rect 29227 35037 29239 35040
rect 29181 35031 29239 35037
rect 30190 35028 30196 35040
rect 30248 35028 30254 35080
rect 30742 35068 30748 35080
rect 30703 35040 30748 35068
rect 30742 35028 30748 35040
rect 30800 35028 30806 35080
rect 31018 35068 31024 35080
rect 30979 35040 31024 35068
rect 31018 35028 31024 35040
rect 31076 35028 31082 35080
rect 30926 35000 30932 35012
rect 26476 34972 27476 35000
rect 30887 34972 30932 35000
rect 26476 34960 26482 34972
rect 30926 34960 30932 34972
rect 30984 34960 30990 35012
rect 22186 34932 22192 34944
rect 21376 34904 22192 34932
rect 18601 34895 18659 34901
rect 22186 34892 22192 34904
rect 22244 34892 22250 34944
rect 22462 34892 22468 34944
rect 22520 34932 22526 34944
rect 22833 34935 22891 34941
rect 22833 34932 22845 34935
rect 22520 34904 22845 34932
rect 22520 34892 22526 34904
rect 22833 34901 22845 34904
rect 22879 34901 22891 34935
rect 23658 34932 23664 34944
rect 23619 34904 23664 34932
rect 22833 34895 22891 34901
rect 23658 34892 23664 34904
rect 23716 34892 23722 34944
rect 26970 34932 26976 34944
rect 26931 34904 26976 34932
rect 26970 34892 26976 34904
rect 27028 34892 27034 34944
rect 28537 34935 28595 34941
rect 28537 34901 28549 34935
rect 28583 34932 28595 34935
rect 29178 34932 29184 34944
rect 28583 34904 29184 34932
rect 28583 34901 28595 34904
rect 28537 34895 28595 34901
rect 29178 34892 29184 34904
rect 29236 34892 29242 34944
rect 30558 34932 30564 34944
rect 30519 34904 30564 34932
rect 30558 34892 30564 34904
rect 30616 34892 30622 34944
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 15838 34728 15844 34740
rect 15799 34700 15844 34728
rect 15838 34688 15844 34700
rect 15896 34688 15902 34740
rect 22097 34731 22155 34737
rect 22097 34697 22109 34731
rect 22143 34728 22155 34731
rect 22278 34728 22284 34740
rect 22143 34700 22284 34728
rect 22143 34697 22155 34700
rect 22097 34691 22155 34697
rect 22278 34688 22284 34700
rect 22336 34688 22342 34740
rect 22646 34728 22652 34740
rect 22388 34700 22652 34728
rect 1578 34592 1584 34604
rect 1539 34564 1584 34592
rect 1578 34552 1584 34564
rect 1636 34552 1642 34604
rect 14550 34592 14556 34604
rect 14511 34564 14556 34592
rect 14550 34552 14556 34564
rect 14608 34552 14614 34604
rect 14734 34592 14740 34604
rect 14695 34564 14740 34592
rect 14734 34552 14740 34564
rect 14792 34552 14798 34604
rect 15381 34595 15439 34601
rect 15381 34561 15393 34595
rect 15427 34561 15439 34595
rect 15381 34555 15439 34561
rect 22281 34595 22339 34601
rect 22281 34561 22293 34595
rect 22327 34592 22339 34595
rect 22388 34592 22416 34700
rect 22646 34688 22652 34700
rect 22704 34728 22710 34740
rect 23217 34731 23275 34737
rect 23217 34728 23229 34731
rect 22704 34700 23229 34728
rect 22704 34688 22710 34700
rect 23217 34697 23229 34700
rect 23263 34697 23275 34731
rect 23382 34728 23388 34740
rect 23343 34700 23388 34728
rect 23217 34691 23275 34697
rect 23382 34688 23388 34700
rect 23440 34688 23446 34740
rect 24394 34728 24400 34740
rect 24355 34700 24400 34728
rect 24394 34688 24400 34700
rect 24452 34688 24458 34740
rect 25409 34731 25467 34737
rect 25409 34697 25421 34731
rect 25455 34728 25467 34731
rect 25682 34728 25688 34740
rect 25455 34700 25688 34728
rect 25455 34697 25467 34700
rect 25409 34691 25467 34697
rect 25682 34688 25688 34700
rect 25740 34688 25746 34740
rect 26896 34700 28304 34728
rect 23017 34663 23075 34669
rect 23017 34660 23029 34663
rect 22480 34632 23029 34660
rect 22480 34601 22508 34632
rect 23017 34629 23029 34632
rect 23063 34629 23075 34663
rect 26896 34660 26924 34700
rect 23017 34623 23075 34629
rect 24964 34632 26924 34660
rect 22327 34564 22416 34592
rect 22465 34595 22523 34601
rect 22327 34561 22339 34564
rect 22281 34555 22339 34561
rect 22465 34561 22477 34595
rect 22511 34561 22523 34595
rect 22465 34555 22523 34561
rect 14645 34527 14703 34533
rect 14645 34493 14657 34527
rect 14691 34524 14703 34527
rect 15194 34524 15200 34536
rect 14691 34496 15200 34524
rect 14691 34493 14703 34496
rect 14645 34487 14703 34493
rect 15194 34484 15200 34496
rect 15252 34524 15258 34536
rect 15396 34524 15424 34555
rect 15252 34496 15424 34524
rect 15252 34484 15258 34496
rect 18690 34484 18696 34536
rect 18748 34524 18754 34536
rect 21450 34524 21456 34536
rect 18748 34496 21456 34524
rect 18748 34484 18754 34496
rect 21450 34484 21456 34496
rect 21508 34524 21514 34536
rect 21508 34496 22140 34524
rect 21508 34484 21514 34496
rect 22112 34456 22140 34496
rect 22186 34484 22192 34536
rect 22244 34524 22250 34536
rect 22480 34524 22508 34555
rect 22554 34552 22560 34604
rect 22612 34592 22618 34604
rect 24578 34592 24584 34604
rect 22612 34564 22657 34592
rect 24539 34564 24584 34592
rect 22612 34552 22618 34564
rect 24578 34552 24584 34564
rect 24636 34552 24642 34604
rect 24964 34524 24992 34632
rect 26970 34620 26976 34672
rect 27028 34660 27034 34672
rect 27402 34663 27460 34669
rect 27402 34660 27414 34663
rect 27028 34632 27414 34660
rect 27028 34620 27034 34632
rect 27402 34629 27414 34632
rect 27448 34629 27460 34663
rect 28276 34660 28304 34700
rect 28350 34688 28356 34740
rect 28408 34728 28414 34740
rect 28537 34731 28595 34737
rect 28537 34728 28549 34731
rect 28408 34700 28549 34728
rect 28408 34688 28414 34700
rect 28537 34697 28549 34700
rect 28583 34697 28595 34731
rect 28994 34728 29000 34740
rect 28955 34700 29000 34728
rect 28537 34691 28595 34697
rect 28994 34688 29000 34700
rect 29052 34688 29058 34740
rect 30098 34660 30104 34672
rect 28276 34632 30104 34660
rect 27402 34623 27460 34629
rect 30098 34620 30104 34632
rect 30156 34620 30162 34672
rect 30558 34669 30564 34672
rect 30552 34660 30564 34669
rect 30519 34632 30564 34660
rect 30552 34623 30564 34632
rect 30558 34620 30564 34623
rect 30616 34620 30622 34672
rect 25130 34552 25136 34604
rect 25188 34592 25194 34604
rect 25225 34595 25283 34601
rect 25225 34592 25237 34595
rect 25188 34564 25237 34592
rect 25188 34552 25194 34564
rect 25225 34561 25237 34564
rect 25271 34561 25283 34595
rect 25225 34555 25283 34561
rect 25406 34552 25412 34604
rect 25464 34592 25470 34604
rect 26053 34595 26111 34601
rect 26053 34592 26065 34595
rect 25464 34564 26065 34592
rect 25464 34552 25470 34564
rect 26053 34561 26065 34564
rect 26099 34561 26111 34595
rect 26053 34555 26111 34561
rect 26237 34595 26295 34601
rect 26237 34561 26249 34595
rect 26283 34592 26295 34595
rect 26694 34592 26700 34604
rect 26283 34564 26700 34592
rect 26283 34561 26295 34564
rect 26237 34555 26295 34561
rect 22244 34496 22508 34524
rect 22572 34496 24992 34524
rect 25041 34527 25099 34533
rect 22244 34484 22250 34496
rect 22572 34456 22600 34496
rect 25041 34493 25053 34527
rect 25087 34524 25099 34527
rect 25958 34524 25964 34536
rect 25087 34496 25964 34524
rect 25087 34493 25099 34496
rect 25041 34487 25099 34493
rect 25958 34484 25964 34496
rect 26016 34484 26022 34536
rect 26068 34524 26096 34555
rect 26694 34552 26700 34564
rect 26752 34552 26758 34604
rect 27062 34552 27068 34604
rect 27120 34592 27126 34604
rect 27157 34595 27215 34601
rect 27157 34592 27169 34595
rect 27120 34564 27169 34592
rect 27120 34552 27126 34564
rect 27157 34561 27169 34564
rect 27203 34561 27215 34595
rect 28166 34592 28172 34604
rect 27157 34555 27215 34561
rect 27264 34564 28172 34592
rect 26326 34524 26332 34536
rect 26068 34496 26188 34524
rect 26287 34496 26332 34524
rect 25866 34456 25872 34468
rect 22112 34428 22600 34456
rect 25827 34428 25872 34456
rect 25866 34416 25872 34428
rect 25924 34416 25930 34468
rect 26160 34456 26188 34496
rect 26326 34484 26332 34496
rect 26384 34484 26390 34536
rect 27264 34524 27292 34564
rect 28166 34552 28172 34564
rect 28224 34552 28230 34604
rect 29178 34592 29184 34604
rect 29139 34564 29184 34592
rect 29178 34552 29184 34564
rect 29236 34552 29242 34604
rect 30282 34592 30288 34604
rect 30243 34564 30288 34592
rect 30282 34552 30288 34564
rect 30340 34552 30346 34604
rect 30834 34592 30840 34604
rect 30392 34564 30840 34592
rect 29362 34524 29368 34536
rect 26436 34496 27292 34524
rect 29323 34496 29368 34524
rect 26436 34456 26464 34496
rect 29362 34484 29368 34496
rect 29420 34484 29426 34536
rect 29457 34527 29515 34533
rect 29457 34493 29469 34527
rect 29503 34524 29515 34527
rect 30392 34524 30420 34564
rect 30834 34552 30840 34564
rect 30892 34592 30898 34604
rect 32214 34592 32220 34604
rect 30892 34564 32220 34592
rect 30892 34552 30898 34564
rect 32214 34552 32220 34564
rect 32272 34552 32278 34604
rect 29503 34496 30420 34524
rect 29503 34493 29515 34496
rect 29457 34487 29515 34493
rect 26160 34428 26464 34456
rect 1762 34388 1768 34400
rect 1723 34360 1768 34388
rect 1762 34348 1768 34360
rect 1820 34348 1826 34400
rect 15010 34348 15016 34400
rect 15068 34388 15074 34400
rect 15473 34391 15531 34397
rect 15473 34388 15485 34391
rect 15068 34360 15485 34388
rect 15068 34348 15074 34360
rect 15473 34357 15485 34360
rect 15519 34357 15531 34391
rect 15473 34351 15531 34357
rect 22554 34348 22560 34400
rect 22612 34388 22618 34400
rect 23201 34391 23259 34397
rect 23201 34388 23213 34391
rect 22612 34360 23213 34388
rect 22612 34348 22618 34360
rect 23201 34357 23213 34360
rect 23247 34357 23259 34391
rect 23201 34351 23259 34357
rect 31386 34348 31392 34400
rect 31444 34388 31450 34400
rect 31665 34391 31723 34397
rect 31665 34388 31677 34391
rect 31444 34360 31677 34388
rect 31444 34348 31450 34360
rect 31665 34357 31677 34360
rect 31711 34357 31723 34391
rect 31665 34351 31723 34357
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 1762 34144 1768 34196
rect 1820 34184 1826 34196
rect 1820 34156 12940 34184
rect 1820 34144 1826 34156
rect 12912 34116 12940 34156
rect 12986 34144 12992 34196
rect 13044 34184 13050 34196
rect 13173 34187 13231 34193
rect 13173 34184 13185 34187
rect 13044 34156 13185 34184
rect 13044 34144 13050 34156
rect 13173 34153 13185 34156
rect 13219 34184 13231 34187
rect 13722 34184 13728 34196
rect 13219 34156 13728 34184
rect 13219 34153 13231 34156
rect 13173 34147 13231 34153
rect 13722 34144 13728 34156
rect 13780 34144 13786 34196
rect 21913 34187 21971 34193
rect 15764 34156 18184 34184
rect 15764 34116 15792 34156
rect 12912 34088 15792 34116
rect 11790 34048 11796 34060
rect 11751 34020 11796 34048
rect 11790 34008 11796 34020
rect 11848 34008 11854 34060
rect 15749 34051 15807 34057
rect 15749 34048 15761 34051
rect 14936 34020 15761 34048
rect 11808 33980 11836 34008
rect 14936 33980 14964 34020
rect 15749 34017 15761 34020
rect 15795 34017 15807 34051
rect 18156 34048 18184 34156
rect 21913 34153 21925 34187
rect 21959 34184 21971 34187
rect 22094 34184 22100 34196
rect 21959 34156 22100 34184
rect 21959 34153 21971 34156
rect 21913 34147 21971 34153
rect 22094 34144 22100 34156
rect 22152 34144 22158 34196
rect 22646 34184 22652 34196
rect 22607 34156 22652 34184
rect 22646 34144 22652 34156
rect 22704 34144 22710 34196
rect 26973 34187 27031 34193
rect 26973 34153 26985 34187
rect 27019 34184 27031 34187
rect 27154 34184 27160 34196
rect 27019 34156 27160 34184
rect 27019 34153 27031 34156
rect 26973 34147 27031 34153
rect 27154 34144 27160 34156
rect 27212 34144 27218 34196
rect 30469 34187 30527 34193
rect 30469 34153 30481 34187
rect 30515 34184 30527 34187
rect 30742 34184 30748 34196
rect 30515 34156 30748 34184
rect 30515 34153 30527 34156
rect 30469 34147 30527 34153
rect 30742 34144 30748 34156
rect 30800 34144 30806 34196
rect 31018 34144 31024 34196
rect 31076 34184 31082 34196
rect 31297 34187 31355 34193
rect 31297 34184 31309 34187
rect 31076 34156 31309 34184
rect 31076 34144 31082 34156
rect 31297 34153 31309 34156
rect 31343 34153 31355 34187
rect 31297 34147 31355 34153
rect 20349 34051 20407 34057
rect 18156 34020 20300 34048
rect 15749 34011 15807 34017
rect 11808 33952 14964 33980
rect 15010 33940 15016 33992
rect 15068 33980 15074 33992
rect 15194 33980 15200 33992
rect 15068 33952 15113 33980
rect 15155 33952 15200 33980
rect 15068 33940 15074 33952
rect 15194 33940 15200 33952
rect 15252 33940 15258 33992
rect 15289 33983 15347 33989
rect 15289 33949 15301 33983
rect 15335 33980 15347 33983
rect 15378 33980 15384 33992
rect 15335 33952 15384 33980
rect 15335 33949 15347 33952
rect 15289 33943 15347 33949
rect 15378 33940 15384 33952
rect 15436 33940 15442 33992
rect 15764 33980 15792 34011
rect 17494 33980 17500 33992
rect 15764 33952 17500 33980
rect 17494 33940 17500 33952
rect 17552 33940 17558 33992
rect 20162 33980 20168 33992
rect 20123 33952 20168 33980
rect 20162 33940 20168 33952
rect 20220 33940 20226 33992
rect 20272 33980 20300 34020
rect 20349 34017 20361 34051
rect 20395 34048 20407 34051
rect 20530 34048 20536 34060
rect 20395 34020 20536 34048
rect 20395 34017 20407 34020
rect 20349 34011 20407 34017
rect 20530 34008 20536 34020
rect 20588 34048 20594 34060
rect 20806 34048 20812 34060
rect 20588 34020 20812 34048
rect 20588 34008 20594 34020
rect 20806 34008 20812 34020
rect 20864 34008 20870 34060
rect 23658 34048 23664 34060
rect 22572 34020 23664 34048
rect 20441 33983 20499 33989
rect 20441 33980 20453 33983
rect 20272 33952 20453 33980
rect 20441 33949 20453 33952
rect 20487 33980 20499 33983
rect 21450 33980 21456 33992
rect 20487 33952 21456 33980
rect 20487 33949 20499 33952
rect 20441 33943 20499 33949
rect 21450 33940 21456 33952
rect 21508 33940 21514 33992
rect 21634 33940 21640 33992
rect 21692 33980 21698 33992
rect 21821 33983 21879 33989
rect 21821 33980 21833 33983
rect 21692 33952 21833 33980
rect 21692 33940 21698 33952
rect 21821 33949 21833 33952
rect 21867 33949 21879 33983
rect 21821 33943 21879 33949
rect 22005 33983 22063 33989
rect 22005 33949 22017 33983
rect 22051 33980 22063 33983
rect 22462 33980 22468 33992
rect 22051 33952 22468 33980
rect 22051 33949 22063 33952
rect 22005 33943 22063 33949
rect 22462 33940 22468 33952
rect 22520 33940 22526 33992
rect 22572 33989 22600 34020
rect 23658 34008 23664 34020
rect 23716 34008 23722 34060
rect 31386 34048 31392 34060
rect 29932 34020 31392 34048
rect 22557 33983 22615 33989
rect 22557 33949 22569 33983
rect 22603 33949 22615 33983
rect 22738 33980 22744 33992
rect 22699 33952 22744 33980
rect 22557 33943 22615 33949
rect 22738 33940 22744 33952
rect 22796 33940 22802 33992
rect 26878 33940 26884 33992
rect 26936 33980 26942 33992
rect 27157 33983 27215 33989
rect 27157 33980 27169 33983
rect 26936 33952 27169 33980
rect 26936 33940 26942 33952
rect 27157 33949 27169 33952
rect 27203 33949 27215 33983
rect 27157 33943 27215 33949
rect 27433 33983 27491 33989
rect 27433 33949 27445 33983
rect 27479 33949 27491 33983
rect 27433 33943 27491 33949
rect 27617 33983 27675 33989
rect 27617 33949 27629 33983
rect 27663 33980 27675 33983
rect 28350 33980 28356 33992
rect 27663 33952 28356 33980
rect 27663 33949 27675 33952
rect 27617 33943 27675 33949
rect 12066 33921 12072 33924
rect 12060 33875 12072 33921
rect 12124 33912 12130 33924
rect 16016 33915 16074 33921
rect 12124 33884 12160 33912
rect 12066 33872 12072 33875
rect 12124 33872 12130 33884
rect 16016 33881 16028 33915
rect 16062 33912 16074 33915
rect 16850 33912 16856 33924
rect 16062 33884 16856 33912
rect 16062 33881 16074 33884
rect 16016 33875 16074 33881
rect 16850 33872 16856 33884
rect 16908 33872 16914 33924
rect 27062 33872 27068 33924
rect 27120 33912 27126 33924
rect 27448 33912 27476 33943
rect 28350 33940 28356 33952
rect 28408 33940 28414 33992
rect 29932 33989 29960 34020
rect 31386 34008 31392 34020
rect 31444 34008 31450 34060
rect 29917 33983 29975 33989
rect 29917 33949 29929 33983
rect 29963 33949 29975 33983
rect 30190 33980 30196 33992
rect 30151 33952 30196 33980
rect 29917 33943 29975 33949
rect 30190 33940 30196 33952
rect 30248 33940 30254 33992
rect 30285 33983 30343 33989
rect 30285 33949 30297 33983
rect 30331 33949 30343 33983
rect 31294 33980 31300 33992
rect 31255 33952 31300 33980
rect 30285 33943 30343 33949
rect 30098 33912 30104 33924
rect 27120 33884 27476 33912
rect 30059 33884 30104 33912
rect 27120 33872 27126 33884
rect 30098 33872 30104 33884
rect 30156 33872 30162 33924
rect 30300 33912 30328 33943
rect 31294 33940 31300 33952
rect 31352 33940 31358 33992
rect 31481 33983 31539 33989
rect 31481 33949 31493 33983
rect 31527 33980 31539 33983
rect 31754 33980 31760 33992
rect 31527 33952 31760 33980
rect 31527 33949 31539 33952
rect 31481 33943 31539 33949
rect 31754 33940 31760 33952
rect 31812 33940 31818 33992
rect 31570 33912 31576 33924
rect 30300 33884 31576 33912
rect 31570 33872 31576 33884
rect 31628 33872 31634 33924
rect 14829 33847 14887 33853
rect 14829 33813 14841 33847
rect 14875 33844 14887 33847
rect 15746 33844 15752 33856
rect 14875 33816 15752 33844
rect 14875 33813 14887 33816
rect 14829 33807 14887 33813
rect 15746 33804 15752 33816
rect 15804 33804 15810 33856
rect 17126 33844 17132 33856
rect 17087 33816 17132 33844
rect 17126 33804 17132 33816
rect 17184 33804 17190 33856
rect 19978 33844 19984 33856
rect 19939 33816 19984 33844
rect 19978 33804 19984 33816
rect 20036 33804 20042 33856
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 11977 33643 12035 33649
rect 11977 33609 11989 33643
rect 12023 33640 12035 33643
rect 12066 33640 12072 33652
rect 12023 33612 12072 33640
rect 12023 33609 12035 33612
rect 11977 33603 12035 33609
rect 12066 33600 12072 33612
rect 12124 33600 12130 33652
rect 14277 33643 14335 33649
rect 14277 33609 14289 33643
rect 14323 33609 14335 33643
rect 16850 33640 16856 33652
rect 16811 33612 16856 33640
rect 14277 33603 14335 33609
rect 11790 33532 11796 33584
rect 11848 33572 11854 33584
rect 14292 33572 14320 33603
rect 16850 33600 16856 33612
rect 16908 33600 16914 33652
rect 20898 33640 20904 33652
rect 20859 33612 20904 33640
rect 20898 33600 20904 33612
rect 20956 33600 20962 33652
rect 14734 33572 14740 33584
rect 11848 33544 12434 33572
rect 14292 33544 14740 33572
rect 11848 33532 11854 33544
rect 12158 33504 12164 33516
rect 12119 33476 12164 33504
rect 12158 33464 12164 33476
rect 12216 33464 12222 33516
rect 12406 33504 12434 33544
rect 14734 33532 14740 33544
rect 14792 33572 14798 33584
rect 14792 33544 15424 33572
rect 14792 33532 14798 33544
rect 12897 33507 12955 33513
rect 12897 33504 12909 33507
rect 12406 33476 12909 33504
rect 12897 33473 12909 33476
rect 12943 33473 12955 33507
rect 12897 33467 12955 33473
rect 13164 33507 13222 33513
rect 13164 33473 13176 33507
rect 13210 33504 13222 33507
rect 14274 33504 14280 33516
rect 13210 33476 14280 33504
rect 13210 33473 13222 33476
rect 13164 33467 13222 33473
rect 14274 33464 14280 33476
rect 14332 33464 14338 33516
rect 14918 33504 14924 33516
rect 14879 33476 14924 33504
rect 14918 33464 14924 33476
rect 14976 33464 14982 33516
rect 15396 33513 15424 33544
rect 17494 33532 17500 33584
rect 17552 33572 17558 33584
rect 19426 33572 19432 33584
rect 17552 33544 19432 33572
rect 17552 33532 17558 33544
rect 19426 33532 19432 33544
rect 19484 33572 19490 33584
rect 19788 33575 19846 33581
rect 19484 33544 19564 33572
rect 19484 33532 19490 33544
rect 15197 33507 15255 33513
rect 15197 33473 15209 33507
rect 15243 33473 15255 33507
rect 15197 33467 15255 33473
rect 15381 33507 15439 33513
rect 15381 33473 15393 33507
rect 15427 33473 15439 33507
rect 17034 33504 17040 33516
rect 16995 33476 17040 33504
rect 15381 33467 15439 33473
rect 12434 33396 12440 33448
rect 12492 33436 12498 33448
rect 12802 33436 12808 33448
rect 12492 33408 12808 33436
rect 12492 33396 12498 33408
rect 12802 33396 12808 33408
rect 12860 33396 12866 33448
rect 15212 33380 15240 33467
rect 17034 33464 17040 33476
rect 17092 33464 17098 33516
rect 17218 33504 17224 33516
rect 17179 33476 17224 33504
rect 17218 33464 17224 33476
rect 17276 33464 17282 33516
rect 18230 33504 18236 33516
rect 18191 33476 18236 33504
rect 18230 33464 18236 33476
rect 18288 33464 18294 33516
rect 19536 33513 19564 33544
rect 19788 33541 19800 33575
rect 19834 33572 19846 33575
rect 19978 33572 19984 33584
rect 19834 33544 19984 33572
rect 19834 33541 19846 33544
rect 19788 33535 19846 33541
rect 19978 33532 19984 33544
rect 20036 33532 20042 33584
rect 19521 33507 19579 33513
rect 19521 33473 19533 33507
rect 19567 33473 19579 33507
rect 31386 33504 31392 33516
rect 31347 33476 31392 33504
rect 19521 33467 19579 33473
rect 31386 33464 31392 33476
rect 31444 33464 31450 33516
rect 35894 33504 35900 33516
rect 35855 33476 35900 33504
rect 35894 33464 35900 33476
rect 35952 33464 35958 33516
rect 17310 33436 17316 33448
rect 17271 33408 17316 33436
rect 17310 33396 17316 33408
rect 17368 33396 17374 33448
rect 17954 33396 17960 33448
rect 18012 33436 18018 33448
rect 18509 33439 18567 33445
rect 18509 33436 18521 33439
rect 18012 33408 18521 33436
rect 18012 33396 18018 33408
rect 18509 33405 18521 33408
rect 18555 33436 18567 33439
rect 19058 33436 19064 33448
rect 18555 33408 19064 33436
rect 18555 33405 18567 33408
rect 18509 33399 18567 33405
rect 19058 33396 19064 33408
rect 19116 33396 19122 33448
rect 31205 33439 31263 33445
rect 31205 33405 31217 33439
rect 31251 33436 31263 33439
rect 36630 33436 36636 33448
rect 31251 33408 31432 33436
rect 36591 33408 36636 33436
rect 31251 33405 31263 33408
rect 31205 33399 31263 33405
rect 31404 33380 31432 33408
rect 36630 33396 36636 33408
rect 36688 33396 36694 33448
rect 15194 33368 15200 33380
rect 15107 33340 15200 33368
rect 15194 33328 15200 33340
rect 15252 33368 15258 33380
rect 18598 33368 18604 33380
rect 15252 33340 18604 33368
rect 15252 33328 15258 33340
rect 18598 33328 18604 33340
rect 18656 33328 18662 33380
rect 31386 33328 31392 33380
rect 31444 33328 31450 33380
rect 12345 33303 12403 33309
rect 12345 33269 12357 33303
rect 12391 33300 12403 33303
rect 12526 33300 12532 33312
rect 12391 33272 12532 33300
rect 12391 33269 12403 33272
rect 12345 33263 12403 33269
rect 12526 33260 12532 33272
rect 12584 33300 12590 33312
rect 13814 33300 13820 33312
rect 12584 33272 13820 33300
rect 12584 33260 12590 33272
rect 13814 33260 13820 33272
rect 13872 33260 13878 33312
rect 14458 33260 14464 33312
rect 14516 33300 14522 33312
rect 14737 33303 14795 33309
rect 14737 33300 14749 33303
rect 14516 33272 14749 33300
rect 14516 33260 14522 33272
rect 14737 33269 14749 33272
rect 14783 33269 14795 33303
rect 18046 33300 18052 33312
rect 18007 33272 18052 33300
rect 14737 33263 14795 33269
rect 18046 33260 18052 33272
rect 18104 33260 18110 33312
rect 18322 33260 18328 33312
rect 18380 33300 18386 33312
rect 18417 33303 18475 33309
rect 18417 33300 18429 33303
rect 18380 33272 18429 33300
rect 18380 33260 18386 33272
rect 18417 33269 18429 33272
rect 18463 33269 18475 33303
rect 18417 33263 18475 33269
rect 21726 33260 21732 33312
rect 21784 33300 21790 33312
rect 23198 33300 23204 33312
rect 21784 33272 23204 33300
rect 21784 33260 21790 33272
rect 23198 33260 23204 33272
rect 23256 33260 23262 33312
rect 31573 33303 31631 33309
rect 31573 33269 31585 33303
rect 31619 33300 31631 33303
rect 31754 33300 31760 33312
rect 31619 33272 31760 33300
rect 31619 33269 31631 33272
rect 31573 33263 31631 33269
rect 31754 33260 31760 33272
rect 31812 33300 31818 33312
rect 32214 33300 32220 33312
rect 31812 33272 32220 33300
rect 31812 33260 31818 33272
rect 32214 33260 32220 33272
rect 32272 33260 32278 33312
rect 47946 33300 47952 33312
rect 47907 33272 47952 33300
rect 47946 33260 47952 33272
rect 48004 33260 48010 33312
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 12158 33056 12164 33108
rect 12216 33096 12222 33108
rect 12345 33099 12403 33105
rect 12345 33096 12357 33099
rect 12216 33068 12357 33096
rect 12216 33056 12222 33068
rect 12345 33065 12357 33068
rect 12391 33065 12403 33099
rect 14274 33096 14280 33108
rect 14235 33068 14280 33096
rect 12345 33059 12403 33065
rect 14274 33056 14280 33068
rect 14332 33056 14338 33108
rect 16393 33099 16451 33105
rect 16393 33065 16405 33099
rect 16439 33096 16451 33099
rect 17034 33096 17040 33108
rect 16439 33068 17040 33096
rect 16439 33065 16451 33068
rect 16393 33059 16451 33065
rect 17034 33056 17040 33068
rect 17092 33056 17098 33108
rect 20162 33056 20168 33108
rect 20220 33096 20226 33108
rect 20441 33099 20499 33105
rect 20441 33096 20453 33099
rect 20220 33068 20453 33096
rect 20220 33056 20226 33068
rect 20441 33065 20453 33068
rect 20487 33065 20499 33099
rect 20441 33059 20499 33065
rect 21910 33056 21916 33108
rect 21968 33096 21974 33108
rect 22278 33096 22284 33108
rect 21968 33068 22284 33096
rect 21968 33056 21974 33068
rect 22278 33056 22284 33068
rect 22336 33056 22342 33108
rect 22741 33099 22799 33105
rect 22741 33065 22753 33099
rect 22787 33096 22799 33099
rect 22830 33096 22836 33108
rect 22787 33068 22836 33096
rect 22787 33065 22799 33068
rect 22741 33059 22799 33065
rect 22830 33056 22836 33068
rect 22888 33056 22894 33108
rect 25961 33099 26019 33105
rect 24596 33068 25912 33096
rect 14918 33028 14924 33040
rect 12544 33000 14924 33028
rect 2041 32895 2099 32901
rect 2041 32861 2053 32895
rect 2087 32892 2099 32895
rect 2130 32892 2136 32904
rect 2087 32864 2136 32892
rect 2087 32861 2099 32864
rect 2041 32855 2099 32861
rect 2130 32852 2136 32864
rect 2188 32852 2194 32904
rect 2498 32892 2504 32904
rect 2459 32864 2504 32892
rect 2498 32852 2504 32864
rect 2556 32892 2562 32904
rect 5258 32892 5264 32904
rect 2556 32864 5264 32892
rect 2556 32852 2562 32864
rect 5258 32852 5264 32864
rect 5316 32852 5322 32904
rect 12544 32901 12572 33000
rect 14918 32988 14924 33000
rect 14976 32988 14982 33040
rect 22002 32988 22008 33040
rect 22060 32988 22066 33040
rect 22094 32988 22100 33040
rect 22152 33028 22158 33040
rect 24596 33028 24624 33068
rect 22152 33000 24624 33028
rect 25884 33028 25912 33068
rect 25961 33065 25973 33099
rect 26007 33096 26019 33099
rect 26326 33096 26332 33108
rect 26007 33068 26332 33096
rect 26007 33065 26019 33068
rect 25961 33059 26019 33065
rect 26326 33056 26332 33068
rect 26384 33056 26390 33108
rect 28813 33099 28871 33105
rect 28813 33065 28825 33099
rect 28859 33096 28871 33099
rect 29362 33096 29368 33108
rect 28859 33068 29368 33096
rect 28859 33065 28871 33068
rect 28813 33059 28871 33065
rect 29362 33056 29368 33068
rect 29420 33056 29426 33108
rect 31205 33099 31263 33105
rect 31205 33065 31217 33099
rect 31251 33096 31263 33099
rect 31294 33096 31300 33108
rect 31251 33068 31300 33096
rect 31251 33065 31263 33068
rect 31205 33059 31263 33065
rect 31294 33056 31300 33068
rect 31352 33056 31358 33108
rect 27062 33028 27068 33040
rect 25884 33000 27068 33028
rect 22152 32988 22158 33000
rect 27062 32988 27068 33000
rect 27120 32988 27126 33040
rect 31846 33028 31852 33040
rect 31807 33000 31852 33028
rect 31846 32988 31852 33000
rect 31904 32988 31910 33040
rect 14366 32920 14372 32972
rect 14424 32960 14430 32972
rect 14737 32963 14795 32969
rect 14737 32960 14749 32963
rect 14424 32932 14749 32960
rect 14424 32920 14430 32932
rect 14737 32929 14749 32932
rect 14783 32960 14795 32963
rect 15010 32960 15016 32972
rect 14783 32932 15016 32960
rect 14783 32929 14795 32932
rect 14737 32923 14795 32929
rect 15010 32920 15016 32932
rect 15068 32920 15074 32972
rect 17494 32960 17500 32972
rect 17455 32932 17500 32960
rect 17494 32920 17500 32932
rect 17552 32920 17558 32972
rect 21542 32960 21548 32972
rect 20916 32932 21548 32960
rect 12529 32895 12587 32901
rect 12529 32861 12541 32895
rect 12575 32892 12587 32895
rect 12618 32892 12624 32904
rect 12575 32864 12624 32892
rect 12575 32861 12587 32864
rect 12529 32855 12587 32861
rect 12618 32852 12624 32864
rect 12676 32852 12682 32904
rect 12805 32895 12863 32901
rect 12805 32861 12817 32895
rect 12851 32861 12863 32895
rect 12986 32892 12992 32904
rect 12947 32864 12992 32892
rect 12805 32855 12863 32861
rect 12820 32824 12848 32855
rect 12986 32852 12992 32864
rect 13044 32852 13050 32904
rect 14458 32892 14464 32904
rect 14419 32864 14464 32892
rect 14458 32852 14464 32864
rect 14516 32852 14522 32904
rect 14645 32895 14703 32901
rect 14645 32861 14657 32895
rect 14691 32861 14703 32895
rect 14645 32855 14703 32861
rect 16577 32895 16635 32901
rect 16577 32861 16589 32895
rect 16623 32861 16635 32895
rect 16850 32892 16856 32904
rect 16811 32864 16856 32892
rect 16577 32855 16635 32861
rect 12894 32824 12900 32836
rect 12820 32796 12900 32824
rect 12894 32784 12900 32796
rect 12952 32784 12958 32836
rect 13814 32784 13820 32836
rect 13872 32824 13878 32836
rect 14660 32824 14688 32855
rect 13872 32796 14688 32824
rect 16592 32824 16620 32855
rect 16850 32852 16856 32864
rect 16908 32852 16914 32904
rect 17037 32895 17095 32901
rect 17037 32861 17049 32895
rect 17083 32892 17095 32895
rect 17126 32892 17132 32904
rect 17083 32864 17132 32892
rect 17083 32861 17095 32864
rect 17037 32855 17095 32861
rect 17126 32852 17132 32864
rect 17184 32852 17190 32904
rect 17764 32895 17822 32901
rect 17764 32861 17776 32895
rect 17810 32892 17822 32895
rect 18046 32892 18052 32904
rect 17810 32864 18052 32892
rect 17810 32861 17822 32864
rect 17764 32855 17822 32861
rect 18046 32852 18052 32864
rect 18104 32852 18110 32904
rect 18506 32852 18512 32904
rect 18564 32892 18570 32904
rect 20916 32901 20944 32932
rect 21542 32920 21548 32932
rect 21600 32920 21606 32972
rect 22020 32960 22048 32988
rect 24578 32960 24584 32972
rect 22020 32932 24584 32960
rect 24578 32920 24584 32932
rect 24636 32920 24642 32972
rect 25590 32920 25596 32972
rect 25648 32960 25654 32972
rect 28905 32963 28963 32969
rect 28905 32960 28917 32963
rect 25648 32932 28917 32960
rect 25648 32920 25654 32932
rect 28905 32929 28917 32932
rect 28951 32960 28963 32963
rect 30650 32960 30656 32972
rect 28951 32932 30656 32960
rect 28951 32929 28963 32932
rect 28905 32923 28963 32929
rect 30650 32920 30656 32932
rect 30708 32920 30714 32972
rect 31478 32960 31484 32972
rect 31220 32932 31484 32960
rect 20625 32895 20683 32901
rect 20625 32892 20637 32895
rect 18564 32864 20637 32892
rect 18564 32852 18570 32864
rect 20625 32861 20637 32864
rect 20671 32861 20683 32895
rect 20625 32855 20683 32861
rect 20901 32895 20959 32901
rect 20901 32861 20913 32895
rect 20947 32861 20959 32895
rect 20901 32855 20959 32861
rect 20990 32852 20996 32904
rect 21048 32892 21054 32904
rect 21085 32895 21143 32901
rect 21085 32892 21097 32895
rect 21048 32864 21097 32892
rect 21048 32852 21054 32864
rect 21085 32861 21097 32864
rect 21131 32861 21143 32895
rect 21818 32892 21824 32904
rect 21085 32855 21143 32861
rect 21192 32864 21824 32892
rect 21192 32824 21220 32864
rect 21818 32852 21824 32864
rect 21876 32852 21882 32904
rect 22097 32895 22155 32901
rect 22097 32861 22109 32895
rect 22143 32861 22155 32895
rect 22097 32855 22155 32861
rect 16592 32796 21220 32824
rect 22112 32824 22140 32855
rect 22278 32852 22284 32904
rect 22336 32892 22342 32904
rect 22925 32895 22983 32901
rect 22336 32864 22381 32892
rect 22336 32852 22342 32864
rect 22925 32861 22937 32895
rect 22971 32892 22983 32895
rect 23014 32892 23020 32904
rect 22971 32864 23020 32892
rect 22971 32861 22983 32864
rect 22925 32855 22983 32861
rect 23014 32852 23020 32864
rect 23072 32852 23078 32904
rect 23198 32892 23204 32904
rect 23159 32864 23204 32892
rect 23198 32852 23204 32864
rect 23256 32892 23262 32904
rect 23256 32864 24992 32892
rect 23256 32852 23262 32864
rect 22370 32824 22376 32836
rect 22112 32796 22376 32824
rect 13872 32784 13878 32796
rect 2314 32716 2320 32768
rect 2372 32756 2378 32768
rect 2593 32759 2651 32765
rect 2593 32756 2605 32759
rect 2372 32728 2605 32756
rect 2372 32716 2378 32728
rect 2593 32725 2605 32728
rect 2639 32725 2651 32759
rect 14660 32756 14688 32796
rect 22370 32784 22376 32796
rect 22428 32784 22434 32836
rect 23934 32784 23940 32836
rect 23992 32824 23998 32836
rect 24826 32827 24884 32833
rect 24826 32824 24838 32827
rect 23992 32796 24838 32824
rect 23992 32784 23998 32796
rect 24826 32793 24838 32796
rect 24872 32793 24884 32827
rect 24964 32824 24992 32864
rect 28534 32852 28540 32904
rect 28592 32892 28598 32904
rect 31220 32901 31248 32932
rect 31478 32920 31484 32932
rect 31536 32920 31542 32972
rect 46477 32963 46535 32969
rect 46477 32929 46489 32963
rect 46523 32960 46535 32963
rect 47946 32960 47952 32972
rect 46523 32932 47952 32960
rect 46523 32929 46535 32932
rect 46477 32923 46535 32929
rect 47946 32920 47952 32932
rect 48004 32920 48010 32972
rect 28629 32895 28687 32901
rect 28629 32892 28641 32895
rect 28592 32864 28641 32892
rect 28592 32852 28598 32864
rect 28629 32861 28641 32864
rect 28675 32861 28687 32895
rect 28629 32855 28687 32861
rect 31205 32895 31263 32901
rect 31205 32861 31217 32895
rect 31251 32861 31263 32895
rect 31386 32892 31392 32904
rect 31347 32864 31392 32892
rect 31205 32855 31263 32861
rect 31386 32852 31392 32864
rect 31444 32852 31450 32904
rect 32125 32895 32183 32901
rect 32125 32861 32137 32895
rect 32171 32892 32183 32895
rect 32214 32892 32220 32904
rect 32171 32864 32220 32892
rect 32171 32861 32183 32864
rect 32125 32855 32183 32861
rect 32214 32852 32220 32864
rect 32272 32852 32278 32904
rect 31570 32824 31576 32836
rect 24964 32796 31576 32824
rect 24826 32787 24884 32793
rect 31570 32784 31576 32796
rect 31628 32784 31634 32836
rect 31849 32827 31907 32833
rect 31849 32793 31861 32827
rect 31895 32824 31907 32827
rect 33502 32824 33508 32836
rect 31895 32796 33508 32824
rect 31895 32793 31907 32796
rect 31849 32787 31907 32793
rect 33502 32784 33508 32796
rect 33560 32784 33566 32836
rect 46661 32827 46719 32833
rect 46661 32793 46673 32827
rect 46707 32824 46719 32827
rect 47854 32824 47860 32836
rect 46707 32796 47860 32824
rect 46707 32793 46719 32796
rect 46661 32787 46719 32793
rect 47854 32784 47860 32796
rect 47912 32784 47918 32836
rect 48314 32824 48320 32836
rect 48275 32796 48320 32824
rect 48314 32784 48320 32796
rect 48372 32784 48378 32836
rect 18322 32756 18328 32768
rect 14660 32728 18328 32756
rect 2593 32719 2651 32725
rect 18322 32716 18328 32728
rect 18380 32716 18386 32768
rect 18874 32756 18880 32768
rect 18835 32728 18880 32756
rect 18874 32716 18880 32728
rect 18932 32716 18938 32768
rect 21174 32716 21180 32768
rect 21232 32756 21238 32768
rect 21637 32759 21695 32765
rect 21637 32756 21649 32759
rect 21232 32728 21649 32756
rect 21232 32716 21238 32728
rect 21637 32725 21649 32728
rect 21683 32725 21695 32759
rect 21637 32719 21695 32725
rect 21726 32716 21732 32768
rect 21784 32756 21790 32768
rect 22094 32756 22100 32768
rect 21784 32728 22100 32756
rect 21784 32716 21790 32728
rect 22094 32716 22100 32728
rect 22152 32716 22158 32768
rect 23109 32759 23167 32765
rect 23109 32725 23121 32759
rect 23155 32756 23167 32759
rect 23382 32756 23388 32768
rect 23155 32728 23388 32756
rect 23155 32725 23167 32728
rect 23109 32719 23167 32725
rect 23382 32716 23388 32728
rect 23440 32716 23446 32768
rect 28445 32759 28503 32765
rect 28445 32725 28457 32759
rect 28491 32756 28503 32759
rect 29086 32756 29092 32768
rect 28491 32728 29092 32756
rect 28491 32725 28503 32728
rect 28445 32719 28503 32725
rect 29086 32716 29092 32728
rect 29144 32716 29150 32768
rect 32033 32759 32091 32765
rect 32033 32725 32045 32759
rect 32079 32756 32091 32759
rect 32122 32756 32128 32768
rect 32079 32728 32128 32756
rect 32079 32725 32091 32728
rect 32033 32719 32091 32725
rect 32122 32716 32128 32728
rect 32180 32716 32186 32768
rect 47302 32716 47308 32768
rect 47360 32756 47366 32768
rect 48130 32756 48136 32768
rect 47360 32728 48136 32756
rect 47360 32716 47366 32728
rect 48130 32716 48136 32728
rect 48188 32716 48194 32768
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 12894 32512 12900 32564
rect 12952 32552 12958 32564
rect 15194 32552 15200 32564
rect 12952 32524 15200 32552
rect 12952 32512 12958 32524
rect 15194 32512 15200 32524
rect 15252 32512 15258 32564
rect 15749 32555 15807 32561
rect 15749 32521 15761 32555
rect 15795 32552 15807 32555
rect 17126 32552 17132 32564
rect 15795 32524 17132 32552
rect 15795 32521 15807 32524
rect 15749 32515 15807 32521
rect 17126 32512 17132 32524
rect 17184 32512 17190 32564
rect 18230 32552 18236 32564
rect 18191 32524 18236 32552
rect 18230 32512 18236 32524
rect 18288 32512 18294 32564
rect 23382 32552 23388 32564
rect 23343 32524 23388 32552
rect 23382 32512 23388 32524
rect 23440 32512 23446 32564
rect 23934 32552 23940 32564
rect 23895 32524 23940 32552
rect 23934 32512 23940 32524
rect 23992 32512 23998 32564
rect 24394 32512 24400 32564
rect 24452 32552 24458 32564
rect 26418 32552 26424 32564
rect 24452 32524 26424 32552
rect 24452 32512 24458 32524
rect 26418 32512 26424 32524
rect 26476 32512 26482 32564
rect 32674 32552 32680 32564
rect 31312 32524 32680 32552
rect 2314 32484 2320 32496
rect 2275 32456 2320 32484
rect 2314 32444 2320 32456
rect 2372 32444 2378 32496
rect 18598 32484 18604 32496
rect 18511 32456 18604 32484
rect 18598 32444 18604 32456
rect 18656 32484 18662 32496
rect 26234 32484 26240 32496
rect 18656 32456 26240 32484
rect 18656 32444 18662 32456
rect 26234 32444 26240 32456
rect 26292 32444 26298 32496
rect 30282 32484 30288 32496
rect 27172 32456 30288 32484
rect 2130 32416 2136 32428
rect 2091 32388 2136 32416
rect 2130 32376 2136 32388
rect 2188 32376 2194 32428
rect 14918 32376 14924 32428
rect 14976 32416 14982 32428
rect 18417 32419 18475 32425
rect 18417 32416 18429 32419
rect 14976 32388 18429 32416
rect 14976 32376 14982 32388
rect 18417 32385 18429 32388
rect 18463 32416 18475 32419
rect 18506 32416 18512 32428
rect 18463 32388 18512 32416
rect 18463 32385 18475 32388
rect 18417 32379 18475 32385
rect 18506 32376 18512 32388
rect 18564 32376 18570 32428
rect 18616 32416 18644 32444
rect 18693 32419 18751 32425
rect 18693 32416 18705 32419
rect 18616 32388 18705 32416
rect 18693 32385 18705 32388
rect 18739 32385 18751 32419
rect 18874 32416 18880 32428
rect 18835 32388 18880 32416
rect 18693 32379 18751 32385
rect 18874 32376 18880 32388
rect 18932 32376 18938 32428
rect 22002 32416 22008 32428
rect 21963 32388 22008 32416
rect 22002 32376 22008 32388
rect 22060 32376 22066 32428
rect 22094 32376 22100 32428
rect 22152 32416 22158 32428
rect 22261 32419 22319 32425
rect 22261 32416 22273 32419
rect 22152 32388 22273 32416
rect 22152 32376 22158 32388
rect 22261 32385 22273 32388
rect 22307 32385 22319 32419
rect 22261 32379 22319 32385
rect 24121 32419 24179 32425
rect 24121 32385 24133 32419
rect 24167 32416 24179 32419
rect 24857 32419 24915 32425
rect 24857 32416 24869 32419
rect 24167 32388 24869 32416
rect 24167 32385 24179 32388
rect 24121 32379 24179 32385
rect 24857 32385 24869 32388
rect 24903 32385 24915 32419
rect 24857 32379 24915 32385
rect 24946 32376 24952 32428
rect 25004 32416 25010 32428
rect 25041 32419 25099 32425
rect 25041 32416 25053 32419
rect 25004 32388 25053 32416
rect 25004 32376 25010 32388
rect 25041 32385 25053 32388
rect 25087 32385 25099 32419
rect 25041 32379 25099 32385
rect 25222 32376 25228 32428
rect 25280 32416 25286 32428
rect 25317 32419 25375 32425
rect 25317 32416 25329 32419
rect 25280 32388 25329 32416
rect 25280 32376 25286 32388
rect 25317 32385 25329 32388
rect 25363 32385 25375 32419
rect 25317 32379 25375 32385
rect 25501 32419 25559 32425
rect 25501 32385 25513 32419
rect 25547 32416 25559 32419
rect 26326 32416 26332 32428
rect 25547 32388 26332 32416
rect 25547 32385 25559 32388
rect 25501 32379 25559 32385
rect 26326 32376 26332 32388
rect 26384 32376 26390 32428
rect 2774 32348 2780 32360
rect 2735 32320 2780 32348
rect 2774 32308 2780 32320
rect 2832 32308 2838 32360
rect 15838 32348 15844 32360
rect 15799 32320 15844 32348
rect 15838 32308 15844 32320
rect 15896 32308 15902 32360
rect 16025 32351 16083 32357
rect 16025 32317 16037 32351
rect 16071 32348 16083 32351
rect 16114 32348 16120 32360
rect 16071 32320 16120 32348
rect 16071 32317 16083 32320
rect 16025 32311 16083 32317
rect 16114 32308 16120 32320
rect 16172 32308 16178 32360
rect 16850 32308 16856 32360
rect 16908 32348 16914 32360
rect 17586 32348 17592 32360
rect 16908 32320 17592 32348
rect 16908 32308 16914 32320
rect 17586 32308 17592 32320
rect 17644 32348 17650 32360
rect 20070 32348 20076 32360
rect 17644 32320 20076 32348
rect 17644 32308 17650 32320
rect 20070 32308 20076 32320
rect 20128 32308 20134 32360
rect 24394 32348 24400 32360
rect 24355 32320 24400 32348
rect 24394 32308 24400 32320
rect 24452 32308 24458 32360
rect 24578 32308 24584 32360
rect 24636 32348 24642 32360
rect 27172 32357 27200 32456
rect 29012 32428 29040 32456
rect 30282 32444 30288 32456
rect 30340 32444 30346 32496
rect 27246 32376 27252 32428
rect 27304 32416 27310 32428
rect 27413 32419 27471 32425
rect 27413 32416 27425 32419
rect 27304 32388 27425 32416
rect 27304 32376 27310 32388
rect 27413 32385 27425 32388
rect 27459 32385 27471 32419
rect 28994 32416 29000 32428
rect 28907 32388 29000 32416
rect 27413 32379 27471 32385
rect 28994 32376 29000 32388
rect 29052 32376 29058 32428
rect 29086 32376 29092 32428
rect 29144 32416 29150 32428
rect 29253 32419 29311 32425
rect 29253 32416 29265 32419
rect 29144 32388 29265 32416
rect 29144 32376 29150 32388
rect 29253 32385 29265 32388
rect 29299 32385 29311 32419
rect 31110 32416 31116 32428
rect 31071 32388 31116 32416
rect 29253 32379 29311 32385
rect 31110 32376 31116 32388
rect 31168 32376 31174 32428
rect 31312 32425 31340 32524
rect 32674 32512 32680 32524
rect 32732 32512 32738 32564
rect 47854 32552 47860 32564
rect 47815 32524 47860 32552
rect 47854 32512 47860 32524
rect 47912 32512 47918 32564
rect 31389 32487 31447 32493
rect 31389 32453 31401 32487
rect 31435 32484 31447 32487
rect 31662 32484 31668 32496
rect 31435 32456 31668 32484
rect 31435 32453 31447 32456
rect 31389 32447 31447 32453
rect 31662 32444 31668 32456
rect 31720 32444 31726 32496
rect 36630 32484 36636 32496
rect 32324 32456 36636 32484
rect 31261 32419 31340 32425
rect 31261 32385 31273 32419
rect 31307 32388 31340 32419
rect 31481 32419 31539 32425
rect 31307 32385 31319 32388
rect 31261 32379 31319 32385
rect 31481 32385 31493 32419
rect 31527 32385 31539 32419
rect 31481 32379 31539 32385
rect 27157 32351 27215 32357
rect 27157 32348 27169 32351
rect 24636 32320 27169 32348
rect 24636 32308 24642 32320
rect 27157 32317 27169 32320
rect 27203 32317 27215 32351
rect 31496 32348 31524 32379
rect 31570 32376 31576 32428
rect 31628 32425 31634 32428
rect 32324 32425 32352 32456
rect 36630 32444 36636 32456
rect 36688 32444 36694 32496
rect 31628 32416 31636 32425
rect 32309 32419 32367 32425
rect 31628 32388 31673 32416
rect 31628 32379 31636 32388
rect 32309 32385 32321 32419
rect 32355 32385 32367 32419
rect 32565 32419 32623 32425
rect 32565 32416 32577 32419
rect 32309 32379 32367 32385
rect 32416 32388 32577 32416
rect 31628 32376 31634 32379
rect 32416 32348 32444 32388
rect 32565 32385 32577 32388
rect 32611 32385 32623 32419
rect 32565 32379 32623 32385
rect 47765 32419 47823 32425
rect 47765 32385 47777 32419
rect 47811 32416 47823 32419
rect 48130 32416 48136 32428
rect 47811 32388 48136 32416
rect 47811 32385 47823 32388
rect 47765 32379 47823 32385
rect 48130 32376 48136 32388
rect 48188 32376 48194 32428
rect 27157 32311 27215 32317
rect 30392 32320 31524 32348
rect 31772 32320 32444 32348
rect 30392 32224 30420 32320
rect 31772 32289 31800 32320
rect 31757 32283 31815 32289
rect 31757 32249 31769 32283
rect 31803 32249 31815 32283
rect 31757 32243 31815 32249
rect 15378 32212 15384 32224
rect 15339 32184 15384 32212
rect 15378 32172 15384 32184
rect 15436 32172 15442 32224
rect 24302 32212 24308 32224
rect 24263 32184 24308 32212
rect 24302 32172 24308 32184
rect 24360 32172 24366 32224
rect 27430 32172 27436 32224
rect 27488 32212 27494 32224
rect 28537 32215 28595 32221
rect 28537 32212 28549 32215
rect 27488 32184 28549 32212
rect 27488 32172 27494 32184
rect 28537 32181 28549 32184
rect 28583 32181 28595 32215
rect 30374 32212 30380 32224
rect 30335 32184 30380 32212
rect 28537 32175 28595 32181
rect 30374 32172 30380 32184
rect 30432 32172 30438 32224
rect 32674 32172 32680 32224
rect 32732 32212 32738 32224
rect 33689 32215 33747 32221
rect 33689 32212 33701 32215
rect 32732 32184 33701 32212
rect 32732 32172 32738 32184
rect 33689 32181 33701 32184
rect 33735 32181 33747 32215
rect 33689 32175 33747 32181
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 21910 32008 21916 32020
rect 21871 31980 21916 32008
rect 21910 31968 21916 31980
rect 21968 31968 21974 32020
rect 23934 32008 23940 32020
rect 23847 31980 23940 32008
rect 23934 31968 23940 31980
rect 23992 32008 23998 32020
rect 24302 32008 24308 32020
rect 23992 31980 24308 32008
rect 23992 31968 23998 31980
rect 24302 31968 24308 31980
rect 24360 31968 24366 32020
rect 24946 32008 24952 32020
rect 24412 31980 24952 32008
rect 24412 31940 24440 31980
rect 24946 31968 24952 31980
rect 25004 31968 25010 32020
rect 25314 31968 25320 32020
rect 25372 32008 25378 32020
rect 25958 32008 25964 32020
rect 25372 31980 25964 32008
rect 25372 31968 25378 31980
rect 25958 31968 25964 31980
rect 26016 31968 26022 32020
rect 27798 32008 27804 32020
rect 26068 31980 27804 32008
rect 22848 31912 24440 31940
rect 1578 31872 1584 31884
rect 1539 31844 1584 31872
rect 1578 31832 1584 31844
rect 1636 31832 1642 31884
rect 17126 31872 17132 31884
rect 16316 31844 17132 31872
rect 1857 31807 1915 31813
rect 1857 31773 1869 31807
rect 1903 31804 1915 31807
rect 6638 31804 6644 31816
rect 1903 31776 6644 31804
rect 1903 31773 1915 31776
rect 1857 31767 1915 31773
rect 6638 31764 6644 31776
rect 6696 31764 6702 31816
rect 12621 31807 12679 31813
rect 12621 31773 12633 31807
rect 12667 31804 12679 31807
rect 13814 31804 13820 31816
rect 12667 31776 13820 31804
rect 12667 31773 12679 31776
rect 12621 31767 12679 31773
rect 13814 31764 13820 31776
rect 13872 31764 13878 31816
rect 16316 31813 16344 31844
rect 17126 31832 17132 31844
rect 17184 31832 17190 31884
rect 19426 31832 19432 31884
rect 19484 31872 19490 31884
rect 20533 31875 20591 31881
rect 20533 31872 20545 31875
rect 19484 31844 20545 31872
rect 19484 31832 19490 31844
rect 20533 31841 20545 31844
rect 20579 31841 20591 31875
rect 20533 31835 20591 31841
rect 16301 31807 16359 31813
rect 16301 31773 16313 31807
rect 16347 31773 16359 31807
rect 16482 31804 16488 31816
rect 16443 31776 16488 31804
rect 16301 31767 16359 31773
rect 16482 31764 16488 31776
rect 16540 31764 16546 31816
rect 21818 31764 21824 31816
rect 21876 31804 21882 31816
rect 22649 31807 22707 31813
rect 22649 31804 22661 31807
rect 21876 31776 22661 31804
rect 21876 31764 21882 31776
rect 22649 31773 22661 31776
rect 22695 31804 22707 31807
rect 22848 31804 22876 31912
rect 23569 31875 23627 31881
rect 23569 31841 23581 31875
rect 23615 31872 23627 31875
rect 24578 31872 24584 31884
rect 23615 31844 24256 31872
rect 24539 31844 24584 31872
rect 23615 31841 23627 31844
rect 23569 31835 23627 31841
rect 22695 31776 22876 31804
rect 22925 31807 22983 31813
rect 22695 31773 22707 31776
rect 22649 31767 22707 31773
rect 22925 31773 22937 31807
rect 22971 31773 22983 31807
rect 22925 31767 22983 31773
rect 23109 31807 23167 31813
rect 23109 31773 23121 31807
rect 23155 31804 23167 31807
rect 23382 31804 23388 31816
rect 23155 31776 23388 31804
rect 23155 31773 23167 31776
rect 23109 31767 23167 31773
rect 20800 31739 20858 31745
rect 20800 31705 20812 31739
rect 20846 31736 20858 31739
rect 20990 31736 20996 31748
rect 20846 31708 20996 31736
rect 20846 31705 20858 31708
rect 20800 31699 20858 31705
rect 20990 31696 20996 31708
rect 21048 31696 21054 31748
rect 22370 31696 22376 31748
rect 22428 31736 22434 31748
rect 22940 31736 22968 31767
rect 23382 31764 23388 31776
rect 23440 31764 23446 31816
rect 23750 31804 23756 31816
rect 23711 31776 23756 31804
rect 23750 31764 23756 31776
rect 23808 31764 23814 31816
rect 24029 31807 24087 31813
rect 24029 31773 24041 31807
rect 24075 31804 24087 31807
rect 24228 31804 24256 31844
rect 24578 31832 24584 31844
rect 24636 31832 24642 31884
rect 24837 31807 24895 31813
rect 24837 31804 24849 31807
rect 24075 31776 24164 31804
rect 24228 31776 24849 31804
rect 24075 31773 24087 31776
rect 24029 31767 24087 31773
rect 22428 31708 22968 31736
rect 24136 31736 24164 31776
rect 24837 31773 24849 31776
rect 24883 31773 24895 31807
rect 26068 31804 26096 31980
rect 27798 31968 27804 31980
rect 27856 31968 27862 32020
rect 28534 32008 28540 32020
rect 28495 31980 28540 32008
rect 28534 31968 28540 31980
rect 28592 31968 28598 32020
rect 31110 31968 31116 32020
rect 31168 32008 31174 32020
rect 31665 32011 31723 32017
rect 31665 32008 31677 32011
rect 31168 31980 31677 32008
rect 31168 31968 31174 31980
rect 31665 31977 31677 31980
rect 31711 31977 31723 32011
rect 31665 31971 31723 31977
rect 32033 32011 32091 32017
rect 32033 31977 32045 32011
rect 32079 32008 32091 32011
rect 32214 32008 32220 32020
rect 32079 31980 32220 32008
rect 32079 31977 32091 31980
rect 32033 31971 32091 31977
rect 32214 31968 32220 31980
rect 32272 32008 32278 32020
rect 32272 31980 32904 32008
rect 32272 31968 32278 31980
rect 30466 31900 30472 31952
rect 30524 31940 30530 31952
rect 32585 31943 32643 31949
rect 32585 31940 32597 31943
rect 30524 31912 32597 31940
rect 30524 31900 30530 31912
rect 32585 31909 32597 31912
rect 32631 31909 32643 31943
rect 32585 31903 32643 31909
rect 27062 31832 27068 31884
rect 27120 31872 27126 31884
rect 32122 31872 32128 31884
rect 27120 31844 27292 31872
rect 32083 31844 32128 31872
rect 27120 31832 27126 31844
rect 24837 31767 24895 31773
rect 24964 31776 26096 31804
rect 24964 31736 24992 31776
rect 26878 31764 26884 31816
rect 26936 31804 26942 31816
rect 27264 31813 27292 31844
rect 32122 31832 32128 31844
rect 32180 31872 32186 31884
rect 32180 31844 32812 31872
rect 32180 31832 32186 31844
rect 32784 31816 32812 31844
rect 26973 31807 27031 31813
rect 26973 31804 26985 31807
rect 26936 31776 26985 31804
rect 26936 31764 26942 31776
rect 26973 31773 26985 31776
rect 27019 31773 27031 31807
rect 26973 31767 27031 31773
rect 27249 31807 27307 31813
rect 27249 31773 27261 31807
rect 27295 31773 27307 31807
rect 27430 31804 27436 31816
rect 27391 31776 27436 31804
rect 27249 31767 27307 31773
rect 24136 31708 24992 31736
rect 26988 31736 27016 31767
rect 27430 31764 27436 31776
rect 27488 31764 27494 31816
rect 28718 31804 28724 31816
rect 27540 31776 28724 31804
rect 27540 31736 27568 31776
rect 28718 31764 28724 31776
rect 28776 31764 28782 31816
rect 28997 31807 29055 31813
rect 28997 31773 29009 31807
rect 29043 31804 29055 31807
rect 29086 31804 29092 31816
rect 29043 31776 29092 31804
rect 29043 31773 29055 31776
rect 28997 31767 29055 31773
rect 29086 31764 29092 31776
rect 29144 31764 29150 31816
rect 29181 31807 29239 31813
rect 29181 31773 29193 31807
rect 29227 31804 29239 31807
rect 30374 31804 30380 31816
rect 29227 31776 30380 31804
rect 29227 31773 29239 31776
rect 29181 31767 29239 31773
rect 30374 31764 30380 31776
rect 30432 31764 30438 31816
rect 31846 31804 31852 31816
rect 31807 31776 31852 31804
rect 31846 31764 31852 31776
rect 31904 31764 31910 31816
rect 32766 31804 32772 31816
rect 32679 31776 32772 31804
rect 32766 31764 32772 31776
rect 32824 31764 32830 31816
rect 32876 31813 32904 31980
rect 32861 31807 32919 31813
rect 32861 31773 32873 31807
rect 32907 31773 32919 31807
rect 32861 31767 32919 31773
rect 32582 31736 32588 31748
rect 26988 31708 27568 31736
rect 32543 31708 32588 31736
rect 22428 31696 22434 31708
rect 12434 31628 12440 31680
rect 12492 31668 12498 31680
rect 16485 31671 16543 31677
rect 12492 31640 12537 31668
rect 12492 31628 12498 31640
rect 16485 31637 16497 31671
rect 16531 31668 16543 31671
rect 16758 31668 16764 31680
rect 16531 31640 16764 31668
rect 16531 31637 16543 31640
rect 16485 31631 16543 31637
rect 16758 31628 16764 31640
rect 16816 31628 16822 31680
rect 22278 31628 22284 31680
rect 22336 31668 22342 31680
rect 22465 31671 22523 31677
rect 22465 31668 22477 31671
rect 22336 31640 22477 31668
rect 22336 31628 22342 31640
rect 22465 31637 22477 31640
rect 22511 31637 22523 31671
rect 22940 31668 22968 31708
rect 32582 31696 32588 31708
rect 32640 31696 32646 31748
rect 25222 31668 25228 31680
rect 22940 31640 25228 31668
rect 22465 31631 22523 31637
rect 25222 31628 25228 31640
rect 25280 31628 25286 31680
rect 26786 31668 26792 31680
rect 26747 31640 26792 31668
rect 26786 31628 26792 31640
rect 26844 31628 26850 31680
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 13814 31464 13820 31476
rect 13775 31436 13820 31464
rect 13814 31424 13820 31436
rect 13872 31424 13878 31476
rect 14277 31467 14335 31473
rect 14277 31433 14289 31467
rect 14323 31464 14335 31467
rect 15378 31464 15384 31476
rect 14323 31436 15384 31464
rect 14323 31433 14335 31436
rect 14277 31427 14335 31433
rect 15378 31424 15384 31436
rect 15436 31424 15442 31476
rect 20990 31464 20996 31476
rect 20951 31436 20996 31464
rect 20990 31424 20996 31436
rect 21048 31424 21054 31476
rect 22094 31424 22100 31476
rect 22152 31464 22158 31476
rect 22152 31436 22197 31464
rect 22152 31424 22158 31436
rect 23750 31424 23756 31476
rect 23808 31464 23814 31476
rect 24673 31467 24731 31473
rect 24673 31464 24685 31467
rect 23808 31436 24685 31464
rect 23808 31424 23814 31436
rect 24673 31433 24685 31436
rect 24719 31433 24731 31467
rect 24673 31427 24731 31433
rect 27157 31467 27215 31473
rect 27157 31433 27169 31467
rect 27203 31464 27215 31467
rect 27246 31464 27252 31476
rect 27203 31436 27252 31464
rect 27203 31433 27215 31436
rect 27157 31427 27215 31433
rect 27246 31424 27252 31436
rect 27304 31424 27310 31476
rect 31297 31467 31355 31473
rect 31297 31433 31309 31467
rect 31343 31464 31355 31467
rect 31386 31464 31392 31476
rect 31343 31436 31392 31464
rect 31343 31433 31355 31436
rect 31297 31427 31355 31433
rect 31386 31424 31392 31436
rect 31444 31424 31450 31476
rect 12244 31399 12302 31405
rect 12244 31365 12256 31399
rect 12290 31396 12302 31399
rect 12434 31396 12440 31408
rect 12290 31368 12440 31396
rect 12290 31365 12302 31368
rect 12244 31359 12302 31365
rect 12434 31356 12440 31368
rect 12492 31356 12498 31408
rect 12618 31356 12624 31408
rect 12676 31396 12682 31408
rect 17310 31396 17316 31408
rect 12676 31368 17316 31396
rect 12676 31356 12682 31368
rect 17310 31356 17316 31368
rect 17368 31356 17374 31408
rect 4608 31331 4666 31337
rect 4608 31297 4620 31331
rect 4654 31328 4666 31331
rect 5994 31328 6000 31340
rect 4654 31300 6000 31328
rect 4654 31297 4666 31300
rect 4608 31291 4666 31297
rect 5994 31288 6000 31300
rect 6052 31288 6058 31340
rect 8386 31328 8392 31340
rect 8347 31300 8392 31328
rect 8386 31288 8392 31300
rect 8444 31288 8450 31340
rect 11790 31288 11796 31340
rect 11848 31328 11854 31340
rect 11977 31331 12035 31337
rect 11977 31328 11989 31331
rect 11848 31300 11989 31328
rect 11848 31288 11854 31300
rect 11977 31297 11989 31300
rect 12023 31297 12035 31331
rect 14185 31331 14243 31337
rect 14185 31328 14197 31331
rect 11977 31291 12035 31297
rect 13556 31300 14197 31328
rect 4341 31263 4399 31269
rect 4341 31229 4353 31263
rect 4387 31229 4399 31263
rect 4341 31223 4399 31229
rect 4356 31124 4384 31223
rect 13556 31136 13584 31300
rect 14185 31297 14197 31300
rect 14231 31297 14243 31331
rect 14185 31291 14243 31297
rect 15473 31331 15531 31337
rect 15473 31297 15485 31331
rect 15519 31328 15531 31331
rect 16850 31328 16856 31340
rect 15519 31300 16620 31328
rect 16811 31300 16856 31328
rect 15519 31297 15531 31300
rect 15473 31291 15531 31297
rect 16592 31272 16620 31300
rect 16850 31288 16856 31300
rect 16908 31288 16914 31340
rect 17034 31328 17040 31340
rect 16995 31300 17040 31328
rect 17034 31288 17040 31300
rect 17092 31288 17098 31340
rect 17586 31328 17592 31340
rect 17547 31300 17592 31328
rect 17586 31288 17592 31300
rect 17644 31288 17650 31340
rect 17773 31331 17831 31337
rect 17773 31297 17785 31331
rect 17819 31297 17831 31331
rect 21174 31328 21180 31340
rect 21135 31300 21180 31328
rect 17773 31291 17831 31297
rect 14090 31220 14096 31272
rect 14148 31260 14154 31272
rect 14458 31260 14464 31272
rect 14148 31232 14464 31260
rect 14148 31220 14154 31232
rect 14458 31220 14464 31232
rect 14516 31220 14522 31272
rect 15562 31260 15568 31272
rect 15523 31232 15568 31260
rect 15562 31220 15568 31232
rect 15620 31220 15626 31272
rect 15838 31260 15844 31272
rect 15799 31232 15844 31260
rect 15838 31220 15844 31232
rect 15896 31220 15902 31272
rect 16574 31220 16580 31272
rect 16632 31260 16638 31272
rect 17788 31260 17816 31291
rect 21174 31288 21180 31300
rect 21232 31288 21238 31340
rect 22278 31328 22284 31340
rect 22239 31300 22284 31328
rect 22278 31288 22284 31300
rect 22336 31288 22342 31340
rect 24854 31328 24860 31340
rect 24815 31300 24860 31328
rect 24854 31288 24860 31300
rect 24912 31288 24918 31340
rect 25133 31331 25191 31337
rect 25133 31297 25145 31331
rect 25179 31297 25191 31331
rect 25314 31328 25320 31340
rect 25275 31300 25320 31328
rect 25133 31291 25191 31297
rect 16632 31232 17816 31260
rect 21453 31263 21511 31269
rect 16632 31220 16638 31232
rect 21453 31229 21465 31263
rect 21499 31260 21511 31263
rect 21542 31260 21548 31272
rect 21499 31232 21548 31260
rect 21499 31229 21511 31232
rect 21453 31223 21511 31229
rect 21542 31220 21548 31232
rect 21600 31220 21606 31272
rect 22462 31220 22468 31272
rect 22520 31260 22526 31272
rect 22557 31263 22615 31269
rect 22557 31260 22569 31263
rect 22520 31232 22569 31260
rect 22520 31220 22526 31232
rect 22557 31229 22569 31232
rect 22603 31260 22615 31263
rect 23198 31260 23204 31272
rect 22603 31232 23204 31260
rect 22603 31229 22615 31232
rect 22557 31223 22615 31229
rect 23198 31220 23204 31232
rect 23256 31220 23262 31272
rect 25148 31260 25176 31291
rect 25314 31288 25320 31300
rect 25372 31288 25378 31340
rect 26786 31288 26792 31340
rect 26844 31328 26850 31340
rect 27341 31331 27399 31337
rect 27341 31328 27353 31331
rect 26844 31300 27353 31328
rect 26844 31288 26850 31300
rect 27341 31297 27353 31300
rect 27387 31297 27399 31331
rect 27341 31291 27399 31297
rect 28994 31288 29000 31340
rect 29052 31328 29058 31340
rect 30190 31337 30196 31340
rect 29917 31331 29975 31337
rect 29917 31328 29929 31331
rect 29052 31300 29929 31328
rect 29052 31288 29058 31300
rect 29917 31297 29929 31300
rect 29963 31297 29975 31331
rect 29917 31291 29975 31297
rect 30184 31291 30196 31337
rect 30248 31328 30254 31340
rect 30248 31300 30284 31328
rect 30190 31288 30196 31291
rect 30248 31288 30254 31300
rect 32122 31288 32128 31340
rect 32180 31328 32186 31340
rect 32493 31331 32551 31337
rect 32493 31328 32505 31331
rect 32180 31300 32505 31328
rect 32180 31288 32186 31300
rect 32493 31297 32505 31300
rect 32539 31297 32551 31331
rect 32493 31291 32551 31297
rect 25222 31260 25228 31272
rect 25148 31232 25228 31260
rect 25222 31220 25228 31232
rect 25280 31220 25286 31272
rect 27617 31263 27675 31269
rect 27617 31229 27629 31263
rect 27663 31260 27675 31263
rect 27798 31260 27804 31272
rect 27663 31232 27804 31260
rect 27663 31229 27675 31232
rect 27617 31223 27675 31229
rect 27798 31220 27804 31232
rect 27856 31220 27862 31272
rect 32585 31263 32643 31269
rect 32585 31229 32597 31263
rect 32631 31260 32643 31263
rect 32674 31260 32680 31272
rect 32631 31232 32680 31260
rect 32631 31229 32643 31232
rect 32585 31223 32643 31229
rect 32674 31220 32680 31232
rect 32732 31220 32738 31272
rect 32766 31220 32772 31272
rect 32824 31260 32830 31272
rect 32861 31263 32919 31269
rect 32861 31260 32873 31263
rect 32824 31232 32873 31260
rect 32824 31220 32830 31232
rect 32861 31229 32873 31232
rect 32907 31229 32919 31263
rect 32861 31223 32919 31229
rect 13630 31152 13636 31204
rect 13688 31192 13694 31204
rect 17681 31195 17739 31201
rect 13688 31164 17080 31192
rect 13688 31152 13694 31164
rect 4706 31124 4712 31136
rect 4356 31096 4712 31124
rect 4706 31084 4712 31096
rect 4764 31084 4770 31136
rect 5350 31084 5356 31136
rect 5408 31124 5414 31136
rect 5721 31127 5779 31133
rect 5721 31124 5733 31127
rect 5408 31096 5733 31124
rect 5408 31084 5414 31096
rect 5721 31093 5733 31096
rect 5767 31093 5779 31127
rect 8202 31124 8208 31136
rect 8163 31096 8208 31124
rect 5721 31087 5779 31093
rect 8202 31084 8208 31096
rect 8260 31084 8266 31136
rect 13357 31127 13415 31133
rect 13357 31093 13369 31127
rect 13403 31124 13415 31127
rect 13538 31124 13544 31136
rect 13403 31096 13544 31124
rect 13403 31093 13415 31096
rect 13357 31087 13415 31093
rect 13538 31084 13544 31096
rect 13596 31084 13602 31136
rect 16482 31084 16488 31136
rect 16540 31124 16546 31136
rect 16945 31127 17003 31133
rect 16945 31124 16957 31127
rect 16540 31096 16957 31124
rect 16540 31084 16546 31096
rect 16945 31093 16957 31096
rect 16991 31093 17003 31127
rect 17052 31124 17080 31164
rect 17681 31161 17693 31195
rect 17727 31192 17739 31195
rect 22370 31192 22376 31204
rect 17727 31164 22376 31192
rect 17727 31161 17739 31164
rect 17681 31155 17739 31161
rect 22370 31152 22376 31164
rect 22428 31152 22434 31204
rect 20438 31124 20444 31136
rect 17052 31096 20444 31124
rect 16945 31087 17003 31093
rect 20438 31084 20444 31096
rect 20496 31084 20502 31136
rect 21361 31127 21419 31133
rect 21361 31093 21373 31127
rect 21407 31124 21419 31127
rect 22465 31127 22523 31133
rect 22465 31124 22477 31127
rect 21407 31096 22477 31124
rect 21407 31093 21419 31096
rect 21361 31087 21419 31093
rect 22465 31093 22477 31096
rect 22511 31124 22523 31127
rect 23934 31124 23940 31136
rect 22511 31096 23940 31124
rect 22511 31093 22523 31096
rect 22465 31087 22523 31093
rect 23934 31084 23940 31096
rect 23992 31124 23998 31136
rect 24762 31124 24768 31136
rect 23992 31096 24768 31124
rect 23992 31084 23998 31096
rect 24762 31084 24768 31096
rect 24820 31084 24826 31136
rect 27522 31124 27528 31136
rect 27483 31096 27528 31124
rect 27522 31084 27528 31096
rect 27580 31084 27586 31136
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 5350 30920 5356 30932
rect 5311 30892 5356 30920
rect 5350 30880 5356 30892
rect 5408 30880 5414 30932
rect 5994 30920 6000 30932
rect 5955 30892 6000 30920
rect 5994 30880 6000 30892
rect 6052 30880 6058 30932
rect 12526 30920 12532 30932
rect 7208 30892 9168 30920
rect 12487 30892 12532 30920
rect 6914 30744 6920 30796
rect 6972 30784 6978 30796
rect 7208 30793 7236 30892
rect 9140 30796 9168 30892
rect 12526 30880 12532 30892
rect 12584 30880 12590 30932
rect 15562 30880 15568 30932
rect 15620 30920 15626 30932
rect 17129 30923 17187 30929
rect 17129 30920 17141 30923
rect 15620 30892 17141 30920
rect 15620 30880 15626 30892
rect 17129 30889 17141 30892
rect 17175 30889 17187 30923
rect 17129 30883 17187 30889
rect 17954 30880 17960 30932
rect 18012 30920 18018 30932
rect 18049 30923 18107 30929
rect 18049 30920 18061 30923
rect 18012 30892 18061 30920
rect 18012 30880 18018 30892
rect 18049 30889 18061 30892
rect 18095 30920 18107 30923
rect 19242 30920 19248 30932
rect 18095 30892 19248 30920
rect 18095 30889 18107 30892
rect 18049 30883 18107 30889
rect 19242 30880 19248 30892
rect 19300 30880 19306 30932
rect 32401 30923 32459 30929
rect 32401 30889 32413 30923
rect 32447 30920 32459 30923
rect 32582 30920 32588 30932
rect 32447 30892 32588 30920
rect 32447 30889 32459 30892
rect 32401 30883 32459 30889
rect 32582 30880 32588 30892
rect 32640 30880 32646 30932
rect 15105 30855 15163 30861
rect 12406 30824 12664 30852
rect 7193 30787 7251 30793
rect 7193 30784 7205 30787
rect 6972 30756 7205 30784
rect 6972 30744 6978 30756
rect 7193 30753 7205 30756
rect 7239 30753 7251 30787
rect 9122 30784 9128 30796
rect 9083 30756 9128 30784
rect 7193 30747 7251 30753
rect 9122 30744 9128 30756
rect 9180 30744 9186 30796
rect 12406 30784 12434 30824
rect 10152 30756 12434 30784
rect 5077 30719 5135 30725
rect 5077 30685 5089 30719
rect 5123 30716 5135 30719
rect 5166 30716 5172 30728
rect 5123 30688 5172 30716
rect 5123 30685 5135 30688
rect 5077 30679 5135 30685
rect 5166 30676 5172 30688
rect 5224 30676 5230 30728
rect 6178 30716 6184 30728
rect 6139 30688 6184 30716
rect 6178 30676 6184 30688
rect 6236 30676 6242 30728
rect 7460 30719 7518 30725
rect 7460 30685 7472 30719
rect 7506 30716 7518 30719
rect 8202 30716 8208 30728
rect 7506 30688 8208 30716
rect 7506 30685 7518 30688
rect 7460 30679 7518 30685
rect 8202 30676 8208 30688
rect 8260 30676 8266 30728
rect 10152 30716 10180 30756
rect 12636 30728 12664 30824
rect 15105 30821 15117 30855
rect 15151 30852 15163 30855
rect 15930 30852 15936 30864
rect 15151 30824 15936 30852
rect 15151 30821 15163 30824
rect 15105 30815 15163 30821
rect 15930 30812 15936 30824
rect 15988 30812 15994 30864
rect 16298 30852 16304 30864
rect 16259 30824 16304 30852
rect 16298 30812 16304 30824
rect 16356 30812 16362 30864
rect 16485 30855 16543 30861
rect 16485 30821 16497 30855
rect 16531 30852 16543 30855
rect 16574 30852 16580 30864
rect 16531 30824 16580 30852
rect 16531 30821 16543 30824
rect 16485 30815 16543 30821
rect 16574 30812 16580 30824
rect 16632 30812 16638 30864
rect 16758 30812 16764 30864
rect 16816 30852 16822 30864
rect 17037 30855 17095 30861
rect 17037 30852 17049 30855
rect 16816 30824 17049 30852
rect 16816 30812 16822 30824
rect 17037 30821 17049 30824
rect 17083 30821 17095 30855
rect 17037 30815 17095 30821
rect 17586 30812 17592 30864
rect 17644 30852 17650 30864
rect 17681 30855 17739 30861
rect 17681 30852 17693 30855
rect 17644 30824 17693 30852
rect 17644 30812 17650 30824
rect 17681 30821 17693 30824
rect 17727 30852 17739 30855
rect 18693 30855 18751 30861
rect 18693 30852 18705 30855
rect 17727 30824 18705 30852
rect 17727 30821 17739 30824
rect 17681 30815 17739 30821
rect 18693 30821 18705 30824
rect 18739 30821 18751 30855
rect 18693 30815 18751 30821
rect 14369 30787 14427 30793
rect 13556 30756 14320 30784
rect 13556 30728 13584 30756
rect 9324 30688 10180 30716
rect 12345 30719 12403 30725
rect 1854 30608 1860 30660
rect 1912 30648 1918 30660
rect 9324 30648 9352 30688
rect 12345 30685 12357 30719
rect 12391 30716 12403 30719
rect 12434 30716 12440 30728
rect 12391 30688 12440 30716
rect 12391 30685 12403 30688
rect 12345 30679 12403 30685
rect 12434 30676 12440 30688
rect 12492 30676 12498 30728
rect 12618 30716 12624 30728
rect 12579 30688 12624 30716
rect 12618 30676 12624 30688
rect 12676 30676 12682 30728
rect 13538 30716 13544 30728
rect 13499 30688 13544 30716
rect 13538 30676 13544 30688
rect 13596 30676 13602 30728
rect 13722 30716 13728 30728
rect 13683 30688 13728 30716
rect 13722 30676 13728 30688
rect 13780 30676 13786 30728
rect 14292 30725 14320 30756
rect 14369 30753 14381 30787
rect 14415 30784 14427 30787
rect 16025 30787 16083 30793
rect 16025 30784 16037 30787
rect 14415 30756 16037 30784
rect 14415 30753 14427 30756
rect 14369 30747 14427 30753
rect 15304 30725 15332 30756
rect 16025 30753 16037 30756
rect 16071 30753 16083 30787
rect 17221 30787 17279 30793
rect 17221 30784 17233 30787
rect 16025 30747 16083 30753
rect 16592 30756 17233 30784
rect 14277 30719 14335 30725
rect 14277 30685 14289 30719
rect 14323 30685 14335 30719
rect 14277 30679 14335 30685
rect 14461 30719 14519 30725
rect 14461 30685 14473 30719
rect 14507 30685 14519 30719
rect 14461 30679 14519 30685
rect 15289 30719 15347 30725
rect 15289 30685 15301 30719
rect 15335 30716 15347 30719
rect 15470 30716 15476 30728
rect 15335 30688 15476 30716
rect 15335 30685 15347 30688
rect 15289 30679 15347 30685
rect 1912 30620 9352 30648
rect 9392 30651 9450 30657
rect 1912 30608 1918 30620
rect 9392 30617 9404 30651
rect 9438 30648 9450 30651
rect 9490 30648 9496 30660
rect 9438 30620 9496 30648
rect 9438 30617 9450 30620
rect 9392 30611 9450 30617
rect 9490 30608 9496 30620
rect 9548 30608 9554 30660
rect 13630 30648 13636 30660
rect 9600 30620 13636 30648
rect 5534 30580 5540 30592
rect 5495 30552 5540 30580
rect 5534 30540 5540 30552
rect 5592 30540 5598 30592
rect 7834 30540 7840 30592
rect 7892 30580 7898 30592
rect 8573 30583 8631 30589
rect 8573 30580 8585 30583
rect 7892 30552 8585 30580
rect 7892 30540 7898 30552
rect 8573 30549 8585 30552
rect 8619 30549 8631 30583
rect 8573 30543 8631 30549
rect 9122 30540 9128 30592
rect 9180 30580 9186 30592
rect 9600 30580 9628 30620
rect 13630 30608 13636 30620
rect 13688 30608 13694 30660
rect 13740 30648 13768 30676
rect 14476 30648 14504 30679
rect 15470 30676 15476 30688
rect 15528 30676 15534 30728
rect 15565 30719 15623 30725
rect 15565 30685 15577 30719
rect 15611 30716 15623 30719
rect 16482 30716 16488 30728
rect 15611 30688 16488 30716
rect 15611 30685 15623 30688
rect 15565 30679 15623 30685
rect 16482 30676 16488 30688
rect 16540 30716 16546 30728
rect 16592 30716 16620 30756
rect 17221 30753 17233 30756
rect 17267 30753 17279 30787
rect 19426 30784 19432 30796
rect 19387 30756 19432 30784
rect 17221 30747 17279 30753
rect 19426 30744 19432 30756
rect 19484 30744 19490 30796
rect 28074 30744 28080 30796
rect 28132 30784 28138 30796
rect 28132 30756 28856 30784
rect 28132 30744 28138 30756
rect 16942 30716 16948 30728
rect 16540 30688 16620 30716
rect 16903 30688 16948 30716
rect 16540 30676 16546 30688
rect 16942 30676 16948 30688
rect 17000 30676 17006 30728
rect 17678 30676 17684 30728
rect 17736 30716 17742 30728
rect 28828 30725 28856 30756
rect 18693 30719 18751 30725
rect 18693 30716 18705 30719
rect 17736 30688 18705 30716
rect 17736 30676 17742 30688
rect 18693 30685 18705 30688
rect 18739 30685 18751 30719
rect 18693 30679 18751 30685
rect 18877 30719 18935 30725
rect 18877 30685 18889 30719
rect 18923 30685 18935 30719
rect 18877 30679 18935 30685
rect 28629 30719 28687 30725
rect 28629 30685 28641 30719
rect 28675 30685 28687 30719
rect 28629 30679 28687 30685
rect 28813 30719 28871 30725
rect 28813 30685 28825 30719
rect 28859 30685 28871 30719
rect 30558 30716 30564 30728
rect 30519 30688 30564 30716
rect 28813 30679 28871 30685
rect 13740 30620 14504 30648
rect 17862 30608 17868 30660
rect 17920 30648 17926 30660
rect 18892 30648 18920 30679
rect 17920 30620 18920 30648
rect 17920 30608 17926 30620
rect 19334 30608 19340 30660
rect 19392 30648 19398 30660
rect 19674 30651 19732 30657
rect 19674 30648 19686 30651
rect 19392 30620 19686 30648
rect 19392 30608 19398 30620
rect 19674 30617 19686 30620
rect 19720 30617 19732 30651
rect 28644 30648 28672 30679
rect 30558 30676 30564 30688
rect 30616 30676 30622 30728
rect 30742 30676 30748 30728
rect 30800 30716 30806 30728
rect 30837 30719 30895 30725
rect 30837 30716 30849 30719
rect 30800 30688 30849 30716
rect 30800 30676 30806 30688
rect 30837 30685 30849 30688
rect 30883 30685 30895 30719
rect 30837 30679 30895 30685
rect 31021 30719 31079 30725
rect 31021 30685 31033 30719
rect 31067 30716 31079 30719
rect 31386 30716 31392 30728
rect 31067 30688 31392 30716
rect 31067 30685 31079 30688
rect 31021 30679 31079 30685
rect 31386 30676 31392 30688
rect 31444 30676 31450 30728
rect 32122 30716 32128 30728
rect 32083 30688 32128 30716
rect 32122 30676 32128 30688
rect 32180 30676 32186 30728
rect 32217 30719 32275 30725
rect 32217 30685 32229 30719
rect 32263 30716 32275 30719
rect 32674 30716 32680 30728
rect 32263 30688 32680 30716
rect 32263 30685 32275 30688
rect 32217 30679 32275 30685
rect 32674 30676 32680 30688
rect 32732 30676 32738 30728
rect 30098 30648 30104 30660
rect 28644 30620 30104 30648
rect 19674 30611 19732 30617
rect 30098 30608 30104 30620
rect 30156 30608 30162 30660
rect 10502 30580 10508 30592
rect 9180 30552 9628 30580
rect 10463 30552 10508 30580
rect 9180 30540 9186 30552
rect 10502 30540 10508 30552
rect 10560 30540 10566 30592
rect 12161 30583 12219 30589
rect 12161 30549 12173 30583
rect 12207 30580 12219 30583
rect 12250 30580 12256 30592
rect 12207 30552 12256 30580
rect 12207 30549 12219 30552
rect 12161 30543 12219 30549
rect 12250 30540 12256 30552
rect 12308 30540 12314 30592
rect 13725 30583 13783 30589
rect 13725 30549 13737 30583
rect 13771 30580 13783 30583
rect 15194 30580 15200 30592
rect 13771 30552 15200 30580
rect 13771 30549 13783 30552
rect 13725 30543 13783 30549
rect 15194 30540 15200 30552
rect 15252 30580 15258 30592
rect 15473 30583 15531 30589
rect 15473 30580 15485 30583
rect 15252 30552 15485 30580
rect 15252 30540 15258 30552
rect 15473 30549 15485 30552
rect 15519 30580 15531 30583
rect 16298 30580 16304 30592
rect 15519 30552 16304 30580
rect 15519 30549 15531 30552
rect 15473 30543 15531 30549
rect 16298 30540 16304 30552
rect 16356 30540 16362 30592
rect 18046 30580 18052 30592
rect 18007 30552 18052 30580
rect 18046 30540 18052 30552
rect 18104 30540 18110 30592
rect 18233 30583 18291 30589
rect 18233 30549 18245 30583
rect 18279 30580 18291 30583
rect 18598 30580 18604 30592
rect 18279 30552 18604 30580
rect 18279 30549 18291 30552
rect 18233 30543 18291 30549
rect 18598 30540 18604 30552
rect 18656 30540 18662 30592
rect 18782 30540 18788 30592
rect 18840 30580 18846 30592
rect 20809 30583 20867 30589
rect 20809 30580 20821 30583
rect 18840 30552 20821 30580
rect 18840 30540 18846 30552
rect 20809 30549 20821 30552
rect 20855 30549 20867 30583
rect 28810 30580 28816 30592
rect 28771 30552 28816 30580
rect 20809 30543 20867 30549
rect 28810 30540 28816 30552
rect 28868 30540 28874 30592
rect 30374 30580 30380 30592
rect 30335 30552 30380 30580
rect 30374 30540 30380 30552
rect 30432 30540 30438 30592
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 5534 30336 5540 30388
rect 5592 30336 5598 30388
rect 5997 30379 6055 30385
rect 5997 30345 6009 30379
rect 6043 30376 6055 30379
rect 6178 30376 6184 30388
rect 6043 30348 6184 30376
rect 6043 30345 6055 30348
rect 5997 30339 6055 30345
rect 6178 30336 6184 30348
rect 6236 30336 6242 30388
rect 7392 30348 7604 30376
rect 5552 30308 5580 30336
rect 6638 30308 6644 30320
rect 5092 30280 5580 30308
rect 6551 30280 6644 30308
rect 5092 30249 5120 30280
rect 6638 30268 6644 30280
rect 6696 30308 6702 30320
rect 7392 30308 7420 30348
rect 6696 30280 7420 30308
rect 7576 30308 7604 30348
rect 8386 30336 8392 30388
rect 8444 30376 8450 30388
rect 9033 30379 9091 30385
rect 9033 30376 9045 30379
rect 8444 30348 9045 30376
rect 8444 30336 8450 30348
rect 9033 30345 9045 30348
rect 9079 30345 9091 30379
rect 9490 30376 9496 30388
rect 9451 30348 9496 30376
rect 9033 30339 9091 30345
rect 9490 30336 9496 30348
rect 9548 30336 9554 30388
rect 16942 30336 16948 30388
rect 17000 30376 17006 30388
rect 17862 30376 17868 30388
rect 17000 30348 17868 30376
rect 17000 30336 17006 30348
rect 17862 30336 17868 30348
rect 17920 30336 17926 30388
rect 19242 30336 19248 30388
rect 19300 30376 19306 30388
rect 19300 30348 23060 30376
rect 19300 30336 19306 30348
rect 23032 30320 23060 30348
rect 23290 30336 23296 30388
rect 23348 30376 23354 30388
rect 23750 30376 23756 30388
rect 23348 30348 23756 30376
rect 23348 30336 23354 30348
rect 23750 30336 23756 30348
rect 23808 30376 23814 30388
rect 24397 30379 24455 30385
rect 24397 30376 24409 30379
rect 23808 30348 24409 30376
rect 23808 30336 23814 30348
rect 24397 30345 24409 30348
rect 24443 30345 24455 30379
rect 30190 30376 30196 30388
rect 30151 30348 30196 30376
rect 24397 30339 24455 30345
rect 30190 30336 30196 30348
rect 30248 30336 30254 30388
rect 11882 30308 11888 30320
rect 7576 30280 11888 30308
rect 6696 30268 6702 30280
rect 11882 30268 11888 30280
rect 11940 30268 11946 30320
rect 17034 30308 17040 30320
rect 16995 30280 17040 30308
rect 17034 30268 17040 30280
rect 17092 30268 17098 30320
rect 17126 30268 17132 30320
rect 17184 30308 17190 30320
rect 17221 30311 17279 30317
rect 17221 30308 17233 30311
rect 17184 30280 17233 30308
rect 17184 30268 17190 30280
rect 17221 30277 17233 30280
rect 17267 30277 17279 30311
rect 17221 30271 17279 30277
rect 17773 30311 17831 30317
rect 17773 30277 17785 30311
rect 17819 30308 17831 30311
rect 18046 30308 18052 30320
rect 17819 30280 18052 30308
rect 17819 30277 17831 30280
rect 17773 30271 17831 30277
rect 18046 30268 18052 30280
rect 18104 30268 18110 30320
rect 18506 30268 18512 30320
rect 18564 30308 18570 30320
rect 18877 30311 18935 30317
rect 18877 30308 18889 30311
rect 18564 30280 18889 30308
rect 18564 30268 18570 30280
rect 18877 30277 18889 30280
rect 18923 30277 18935 30311
rect 18877 30271 18935 30277
rect 18969 30311 19027 30317
rect 18969 30277 18981 30311
rect 19015 30308 19027 30311
rect 19426 30308 19432 30320
rect 19015 30280 19432 30308
rect 19015 30277 19027 30280
rect 18969 30271 19027 30277
rect 5077 30243 5135 30249
rect 5077 30209 5089 30243
rect 5123 30209 5135 30243
rect 5077 30203 5135 30209
rect 5166 30200 5172 30252
rect 5224 30240 5230 30252
rect 5537 30243 5595 30249
rect 5537 30240 5549 30243
rect 5224 30212 5549 30240
rect 5224 30200 5230 30212
rect 5537 30209 5549 30212
rect 5583 30240 5595 30243
rect 6825 30243 6883 30249
rect 6825 30240 6837 30243
rect 5583 30212 6837 30240
rect 5583 30209 5595 30212
rect 5537 30203 5595 30209
rect 6825 30209 6837 30212
rect 6871 30240 6883 30243
rect 7374 30240 7380 30252
rect 6871 30212 7380 30240
rect 6871 30209 6883 30212
rect 6825 30203 6883 30209
rect 7374 30200 7380 30212
rect 7432 30200 7438 30252
rect 7469 30243 7527 30249
rect 7469 30209 7481 30243
rect 7515 30240 7527 30243
rect 7834 30240 7840 30252
rect 7515 30212 7840 30240
rect 7515 30209 7527 30212
rect 7469 30203 7527 30209
rect 7475 30172 7503 30203
rect 7834 30200 7840 30212
rect 7892 30200 7898 30252
rect 8573 30243 8631 30249
rect 8573 30209 8585 30243
rect 8619 30209 8631 30243
rect 8573 30203 8631 30209
rect 7742 30172 7748 30184
rect 7300 30144 7503 30172
rect 7703 30144 7748 30172
rect 4890 30036 4896 30048
rect 4851 30008 4896 30036
rect 4890 29996 4896 30008
rect 4948 29996 4954 30048
rect 5813 30039 5871 30045
rect 5813 30005 5825 30039
rect 5859 30036 5871 30039
rect 7300 30036 7328 30144
rect 7742 30132 7748 30144
rect 7800 30172 7806 30184
rect 8588 30172 8616 30203
rect 8662 30200 8668 30252
rect 8720 30240 8726 30252
rect 12250 30249 12256 30252
rect 9677 30243 9735 30249
rect 9677 30240 9689 30243
rect 8720 30212 9689 30240
rect 8720 30200 8726 30212
rect 9677 30209 9689 30212
rect 9723 30209 9735 30243
rect 12244 30240 12256 30249
rect 12211 30212 12256 30240
rect 9677 30203 9735 30209
rect 12244 30203 12256 30212
rect 12250 30200 12256 30203
rect 12308 30200 12314 30252
rect 15194 30240 15200 30252
rect 15155 30212 15200 30240
rect 15194 30200 15200 30212
rect 15252 30200 15258 30252
rect 15470 30240 15476 30252
rect 15431 30212 15476 30240
rect 15470 30200 15476 30212
rect 15528 30200 15534 30252
rect 16850 30240 16856 30252
rect 16763 30212 16856 30240
rect 16850 30200 16856 30212
rect 16908 30200 16914 30252
rect 17678 30240 17684 30252
rect 17639 30212 17684 30240
rect 17678 30200 17684 30212
rect 17736 30200 17742 30252
rect 17862 30240 17868 30252
rect 17823 30212 17868 30240
rect 17862 30200 17868 30212
rect 17920 30200 17926 30252
rect 18598 30240 18604 30252
rect 18559 30212 18604 30240
rect 18598 30200 18604 30212
rect 18656 30200 18662 30252
rect 18782 30249 18788 30252
rect 18749 30243 18788 30249
rect 18749 30209 18761 30243
rect 18749 30203 18788 30209
rect 18782 30200 18788 30203
rect 18840 30200 18846 30252
rect 11974 30172 11980 30184
rect 7800 30144 8616 30172
rect 11935 30144 11980 30172
rect 7800 30132 7806 30144
rect 11974 30132 11980 30144
rect 12032 30132 12038 30184
rect 16868 30172 16896 30200
rect 18800 30172 18828 30200
rect 16868 30144 18828 30172
rect 18892 30172 18920 30271
rect 19426 30268 19432 30280
rect 19484 30268 19490 30320
rect 22370 30308 22376 30320
rect 22331 30280 22376 30308
rect 22370 30268 22376 30280
rect 22428 30308 22434 30320
rect 22925 30311 22983 30317
rect 22925 30308 22937 30311
rect 22428 30280 22937 30308
rect 22428 30268 22434 30280
rect 22925 30277 22937 30280
rect 22971 30277 22983 30311
rect 22925 30271 22983 30277
rect 23014 30268 23020 30320
rect 23072 30268 23078 30320
rect 23141 30311 23199 30317
rect 23141 30308 23153 30311
rect 23124 30277 23153 30308
rect 23187 30308 23199 30311
rect 23566 30308 23572 30320
rect 23187 30280 23572 30308
rect 23187 30277 23199 30280
rect 23124 30271 23199 30277
rect 19058 30200 19064 30252
rect 19116 30249 19122 30252
rect 19116 30240 19124 30249
rect 19116 30212 19161 30240
rect 19116 30203 19124 30212
rect 19116 30200 19122 30203
rect 20622 30200 20628 30252
rect 20680 30240 20686 30252
rect 22189 30243 22247 30249
rect 22189 30240 22201 30243
rect 20680 30212 22201 30240
rect 20680 30200 20686 30212
rect 22189 30209 22201 30212
rect 22235 30209 22247 30243
rect 22189 30203 22247 30209
rect 20254 30172 20260 30184
rect 18892 30144 20260 30172
rect 20254 30132 20260 30144
rect 20312 30132 20318 30184
rect 22204 30172 22232 30203
rect 22462 30200 22468 30252
rect 22520 30240 22526 30252
rect 22520 30212 22565 30240
rect 22520 30200 22526 30212
rect 23124 30172 23152 30271
rect 23566 30268 23572 30280
rect 23624 30268 23630 30320
rect 24305 30311 24363 30317
rect 24305 30277 24317 30311
rect 24351 30308 24363 30311
rect 25130 30308 25136 30320
rect 24351 30280 25136 30308
rect 24351 30277 24363 30280
rect 24305 30271 24363 30277
rect 22204 30144 23152 30172
rect 7466 30064 7472 30116
rect 7524 30104 7530 30116
rect 7653 30107 7711 30113
rect 7653 30104 7665 30107
rect 7524 30076 7665 30104
rect 7524 30064 7530 30076
rect 7653 30073 7665 30076
rect 7699 30073 7711 30107
rect 16758 30104 16764 30116
rect 7653 30067 7711 30073
rect 15580 30076 16764 30104
rect 5859 30008 7328 30036
rect 7561 30039 7619 30045
rect 5859 30005 5871 30008
rect 5813 29999 5871 30005
rect 7561 30005 7573 30039
rect 7607 30036 7619 30039
rect 8386 30036 8392 30048
rect 7607 30008 8392 30036
rect 7607 30005 7619 30008
rect 7561 29999 7619 30005
rect 8386 29996 8392 30008
rect 8444 29996 8450 30048
rect 8849 30039 8907 30045
rect 8849 30005 8861 30039
rect 8895 30036 8907 30039
rect 10502 30036 10508 30048
rect 8895 30008 10508 30036
rect 8895 30005 8907 30008
rect 8849 29999 8907 30005
rect 10502 29996 10508 30008
rect 10560 29996 10566 30048
rect 13078 29996 13084 30048
rect 13136 30036 13142 30048
rect 13357 30039 13415 30045
rect 13357 30036 13369 30039
rect 13136 30008 13369 30036
rect 13136 29996 13142 30008
rect 13357 30005 13369 30008
rect 13403 30036 13415 30039
rect 13722 30036 13728 30048
rect 13403 30008 13728 30036
rect 13403 30005 13415 30008
rect 13357 29999 13415 30005
rect 13722 29996 13728 30008
rect 13780 29996 13786 30048
rect 15580 30045 15608 30076
rect 16758 30064 16764 30076
rect 16816 30104 16822 30116
rect 17678 30104 17684 30116
rect 16816 30076 17684 30104
rect 16816 30064 16822 30076
rect 17678 30064 17684 30076
rect 17736 30064 17742 30116
rect 19245 30107 19303 30113
rect 19245 30073 19257 30107
rect 19291 30104 19303 30107
rect 19334 30104 19340 30116
rect 19291 30076 19340 30104
rect 19291 30073 19303 30076
rect 19245 30067 19303 30073
rect 19334 30064 19340 30076
rect 19392 30064 19398 30116
rect 19518 30064 19524 30116
rect 19576 30104 19582 30116
rect 22554 30104 22560 30116
rect 19576 30076 22560 30104
rect 19576 30064 19582 30076
rect 22554 30064 22560 30076
rect 22612 30064 22618 30116
rect 22646 30064 22652 30116
rect 22704 30104 22710 30116
rect 24320 30104 24348 30271
rect 25130 30268 25136 30280
rect 25188 30308 25194 30320
rect 26602 30308 26608 30320
rect 25188 30280 26608 30308
rect 25188 30268 25194 30280
rect 26602 30268 26608 30280
rect 26660 30268 26666 30320
rect 27890 30308 27896 30320
rect 27851 30280 27896 30308
rect 27890 30268 27896 30280
rect 27948 30268 27954 30320
rect 41322 30268 41328 30320
rect 41380 30308 41386 30320
rect 47670 30308 47676 30320
rect 41380 30280 47676 30308
rect 41380 30268 41386 30280
rect 47670 30268 47676 30280
rect 47728 30268 47734 30320
rect 25682 30200 25688 30252
rect 25740 30240 25746 30252
rect 26053 30243 26111 30249
rect 26053 30240 26065 30243
rect 25740 30212 26065 30240
rect 25740 30200 25746 30212
rect 26053 30209 26065 30212
rect 26099 30209 26111 30243
rect 26053 30203 26111 30209
rect 26234 30200 26240 30252
rect 26292 30240 26298 30252
rect 26329 30243 26387 30249
rect 26329 30240 26341 30243
rect 26292 30212 26341 30240
rect 26292 30200 26298 30212
rect 26329 30209 26341 30212
rect 26375 30209 26387 30243
rect 26510 30240 26516 30252
rect 26471 30212 26516 30240
rect 26329 30203 26387 30209
rect 26510 30200 26516 30212
rect 26568 30200 26574 30252
rect 28074 30240 28080 30252
rect 28035 30212 28080 30240
rect 28074 30200 28080 30212
rect 28132 30200 28138 30252
rect 28353 30243 28411 30249
rect 28353 30209 28365 30243
rect 28399 30240 28411 30243
rect 28810 30240 28816 30252
rect 28399 30212 28816 30240
rect 28399 30209 28411 30212
rect 28353 30203 28411 30209
rect 28810 30200 28816 30212
rect 28868 30240 28874 30252
rect 28997 30243 29055 30249
rect 28997 30240 29009 30243
rect 28868 30212 29009 30240
rect 28868 30200 28874 30212
rect 28997 30209 29009 30212
rect 29043 30209 29055 30243
rect 30374 30240 30380 30252
rect 30335 30212 30380 30240
rect 28997 30203 29055 30209
rect 30374 30200 30380 30212
rect 30432 30200 30438 30252
rect 30653 30243 30711 30249
rect 30653 30209 30665 30243
rect 30699 30240 30711 30243
rect 30834 30240 30840 30252
rect 30699 30212 30840 30240
rect 30699 30209 30711 30212
rect 30653 30203 30711 30209
rect 30834 30200 30840 30212
rect 30892 30240 30898 30252
rect 30892 30212 31754 30240
rect 30892 30200 30898 30212
rect 28261 30175 28319 30181
rect 28261 30141 28273 30175
rect 28307 30172 28319 30175
rect 29089 30175 29147 30181
rect 29089 30172 29101 30175
rect 28307 30144 29101 30172
rect 28307 30141 28319 30144
rect 28261 30135 28319 30141
rect 29089 30141 29101 30144
rect 29135 30172 29147 30175
rect 30466 30172 30472 30184
rect 29135 30144 30472 30172
rect 29135 30141 29147 30144
rect 29089 30135 29147 30141
rect 30466 30132 30472 30144
rect 30524 30132 30530 30184
rect 31726 30172 31754 30212
rect 32858 30200 32864 30252
rect 32916 30240 32922 30252
rect 47302 30240 47308 30252
rect 32916 30212 47308 30240
rect 32916 30200 32922 30212
rect 47302 30200 47308 30212
rect 47360 30240 47366 30252
rect 47765 30243 47823 30249
rect 47765 30240 47777 30243
rect 47360 30212 47777 30240
rect 47360 30200 47366 30212
rect 47765 30209 47777 30212
rect 47811 30209 47823 30243
rect 47765 30203 47823 30209
rect 31846 30172 31852 30184
rect 31726 30144 31852 30172
rect 31846 30132 31852 30144
rect 31904 30132 31910 30184
rect 22704 30076 24348 30104
rect 22704 30064 22710 30076
rect 15565 30039 15623 30045
rect 15565 30005 15577 30039
rect 15611 30005 15623 30039
rect 15746 30036 15752 30048
rect 15707 30008 15752 30036
rect 15565 29999 15623 30005
rect 15746 29996 15752 30008
rect 15804 29996 15810 30048
rect 15930 29996 15936 30048
rect 15988 30036 15994 30048
rect 21634 30036 21640 30048
rect 15988 30008 21640 30036
rect 15988 29996 15994 30008
rect 21634 29996 21640 30008
rect 21692 29996 21698 30048
rect 22005 30039 22063 30045
rect 22005 30005 22017 30039
rect 22051 30036 22063 30039
rect 22370 30036 22376 30048
rect 22051 30008 22376 30036
rect 22051 30005 22063 30008
rect 22005 29999 22063 30005
rect 22370 29996 22376 30008
rect 22428 29996 22434 30048
rect 22462 29996 22468 30048
rect 22520 30036 22526 30048
rect 23109 30039 23167 30045
rect 23109 30036 23121 30039
rect 22520 30008 23121 30036
rect 22520 29996 22526 30008
rect 23109 30005 23121 30008
rect 23155 30005 23167 30039
rect 23290 30036 23296 30048
rect 23251 30008 23296 30036
rect 23109 29999 23167 30005
rect 23290 29996 23296 30008
rect 23348 29996 23354 30048
rect 25869 30039 25927 30045
rect 25869 30005 25881 30039
rect 25915 30036 25927 30039
rect 26326 30036 26332 30048
rect 25915 30008 26332 30036
rect 25915 30005 25927 30008
rect 25869 29999 25927 30005
rect 26326 29996 26332 30008
rect 26384 29996 26390 30048
rect 29270 29996 29276 30048
rect 29328 30036 29334 30048
rect 29365 30039 29423 30045
rect 29365 30036 29377 30039
rect 29328 30008 29377 30036
rect 29328 29996 29334 30008
rect 29365 30005 29377 30008
rect 29411 30005 29423 30039
rect 29365 29999 29423 30005
rect 30561 30039 30619 30045
rect 30561 30005 30573 30039
rect 30607 30036 30619 30039
rect 31018 30036 31024 30048
rect 30607 30008 31024 30036
rect 30607 30005 30619 30008
rect 30561 29999 30619 30005
rect 31018 29996 31024 30008
rect 31076 29996 31082 30048
rect 46474 29996 46480 30048
rect 46532 30036 46538 30048
rect 47213 30039 47271 30045
rect 47213 30036 47225 30039
rect 46532 30008 47225 30036
rect 46532 29996 46538 30008
rect 47213 30005 47225 30008
rect 47259 30005 47271 30039
rect 47854 30036 47860 30048
rect 47815 30008 47860 30036
rect 47213 29999 47271 30005
rect 47854 29996 47860 30008
rect 47912 29996 47918 30048
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 12434 29792 12440 29844
rect 12492 29832 12498 29844
rect 15746 29832 15752 29844
rect 12492 29804 12537 29832
rect 15707 29804 15752 29832
rect 12492 29792 12498 29804
rect 15746 29792 15752 29804
rect 15804 29792 15810 29844
rect 20622 29832 20628 29844
rect 20583 29804 20628 29832
rect 20622 29792 20628 29804
rect 20680 29792 20686 29844
rect 22097 29835 22155 29841
rect 22097 29801 22109 29835
rect 22143 29832 22155 29835
rect 22186 29832 22192 29844
rect 22143 29804 22192 29832
rect 22143 29801 22155 29804
rect 22097 29795 22155 29801
rect 22186 29792 22192 29804
rect 22244 29792 22250 29844
rect 22370 29792 22376 29844
rect 22428 29832 22434 29844
rect 23109 29835 23167 29841
rect 23109 29832 23121 29835
rect 22428 29804 23121 29832
rect 22428 29792 22434 29804
rect 23109 29801 23121 29804
rect 23155 29801 23167 29835
rect 23109 29795 23167 29801
rect 23474 29792 23480 29844
rect 23532 29832 23538 29844
rect 30098 29832 30104 29844
rect 23532 29804 28994 29832
rect 30059 29804 30104 29832
rect 23532 29792 23538 29804
rect 15841 29767 15899 29773
rect 15841 29733 15853 29767
rect 15887 29764 15899 29767
rect 20901 29767 20959 29773
rect 20901 29764 20913 29767
rect 15887 29736 20913 29764
rect 15887 29733 15899 29736
rect 15841 29727 15899 29733
rect 20901 29733 20913 29736
rect 20947 29733 20959 29767
rect 22462 29764 22468 29776
rect 20901 29727 20959 29733
rect 21652 29736 22468 29764
rect 6914 29696 6920 29708
rect 6875 29668 6920 29696
rect 6914 29656 6920 29668
rect 6972 29656 6978 29708
rect 15473 29699 15531 29705
rect 15473 29665 15485 29699
rect 15519 29696 15531 29699
rect 19518 29696 19524 29708
rect 15519 29668 19524 29696
rect 15519 29665 15531 29668
rect 15473 29659 15531 29665
rect 19518 29656 19524 29668
rect 19576 29656 19582 29708
rect 20916 29696 20944 29727
rect 21652 29708 21680 29736
rect 22462 29724 22468 29736
rect 22520 29724 22526 29776
rect 22741 29767 22799 29773
rect 22741 29733 22753 29767
rect 22787 29764 22799 29767
rect 23290 29764 23296 29776
rect 22787 29736 23296 29764
rect 22787 29733 22799 29736
rect 22741 29727 22799 29733
rect 23290 29724 23296 29736
rect 23348 29724 23354 29776
rect 28966 29764 28994 29804
rect 30098 29792 30104 29804
rect 30156 29792 30162 29844
rect 31662 29764 31668 29776
rect 28966 29736 31668 29764
rect 31662 29724 31668 29736
rect 31720 29724 31726 29776
rect 20916 29668 21588 29696
rect 4341 29631 4399 29637
rect 4341 29597 4353 29631
rect 4387 29597 4399 29631
rect 4341 29591 4399 29597
rect 4608 29631 4666 29637
rect 4608 29597 4620 29631
rect 4654 29628 4666 29631
rect 4890 29628 4896 29640
rect 4654 29600 4896 29628
rect 4654 29597 4666 29600
rect 4608 29591 4666 29597
rect 4356 29560 4384 29591
rect 4890 29588 4896 29600
rect 4948 29588 4954 29640
rect 12621 29631 12679 29637
rect 12621 29597 12633 29631
rect 12667 29628 12679 29631
rect 12710 29628 12716 29640
rect 12667 29600 12716 29628
rect 12667 29597 12679 29600
rect 12621 29591 12679 29597
rect 12710 29588 12716 29600
rect 12768 29588 12774 29640
rect 12894 29628 12900 29640
rect 12855 29600 12900 29628
rect 12894 29588 12900 29600
rect 12952 29588 12958 29640
rect 13078 29628 13084 29640
rect 13039 29600 13084 29628
rect 13078 29588 13084 29600
rect 13136 29588 13142 29640
rect 15930 29628 15936 29640
rect 15891 29600 15936 29628
rect 15930 29588 15936 29600
rect 15988 29588 15994 29640
rect 16022 29588 16028 29640
rect 16080 29628 16086 29640
rect 16209 29631 16267 29637
rect 16209 29628 16221 29631
rect 16080 29600 16221 29628
rect 16080 29588 16086 29600
rect 16209 29597 16221 29600
rect 16255 29597 16267 29631
rect 16209 29591 16267 29597
rect 20349 29631 20407 29637
rect 20349 29597 20361 29631
rect 20395 29597 20407 29631
rect 20714 29628 20720 29640
rect 20675 29600 20720 29628
rect 20349 29591 20407 29597
rect 4706 29560 4712 29572
rect 4356 29532 4712 29560
rect 4706 29520 4712 29532
rect 4764 29560 4770 29572
rect 6914 29560 6920 29572
rect 4764 29532 6920 29560
rect 4764 29520 4770 29532
rect 6914 29520 6920 29532
rect 6972 29520 6978 29572
rect 7184 29563 7242 29569
rect 7184 29529 7196 29563
rect 7230 29560 7242 29563
rect 7282 29560 7288 29572
rect 7230 29532 7288 29560
rect 7230 29529 7242 29532
rect 7184 29523 7242 29529
rect 7282 29520 7288 29532
rect 7340 29520 7346 29572
rect 20364 29560 20392 29591
rect 20714 29588 20720 29600
rect 20772 29588 20778 29640
rect 21266 29588 21272 29640
rect 21324 29628 21330 29640
rect 21560 29637 21588 29668
rect 21634 29656 21640 29708
rect 21692 29696 21698 29708
rect 23658 29696 23664 29708
rect 21692 29668 21737 29696
rect 21836 29668 23664 29696
rect 21692 29656 21698 29668
rect 21361 29631 21419 29637
rect 21361 29628 21373 29631
rect 21324 29600 21373 29628
rect 21324 29588 21330 29600
rect 21361 29597 21373 29600
rect 21407 29597 21419 29631
rect 21361 29591 21419 29597
rect 21545 29631 21603 29637
rect 21545 29597 21557 29631
rect 21591 29597 21603 29631
rect 21545 29591 21603 29597
rect 21729 29631 21787 29637
rect 21729 29597 21741 29631
rect 21775 29628 21787 29631
rect 21836 29628 21864 29668
rect 23658 29656 23664 29668
rect 23716 29656 23722 29708
rect 24578 29656 24584 29708
rect 24636 29696 24642 29708
rect 25409 29699 25467 29705
rect 25409 29696 25421 29699
rect 24636 29668 25421 29696
rect 24636 29656 24642 29668
rect 25409 29665 25421 29668
rect 25455 29665 25467 29699
rect 46474 29696 46480 29708
rect 46435 29668 46480 29696
rect 25409 29659 25467 29665
rect 21775 29600 21864 29628
rect 21913 29631 21971 29637
rect 21775 29597 21787 29600
rect 21729 29591 21787 29597
rect 21913 29597 21925 29631
rect 21959 29597 21971 29631
rect 21913 29591 21971 29597
rect 21284 29560 21312 29588
rect 20364 29532 21312 29560
rect 5718 29492 5724 29504
rect 5679 29464 5724 29492
rect 5718 29452 5724 29464
rect 5776 29452 5782 29504
rect 8294 29492 8300 29504
rect 8255 29464 8300 29492
rect 8294 29452 8300 29464
rect 8352 29452 8358 29504
rect 16117 29495 16175 29501
rect 16117 29461 16129 29495
rect 16163 29492 16175 29495
rect 16666 29492 16672 29504
rect 16163 29464 16672 29492
rect 16163 29461 16175 29464
rect 16117 29455 16175 29461
rect 16666 29452 16672 29464
rect 16724 29452 16730 29504
rect 20714 29452 20720 29504
rect 20772 29492 20778 29504
rect 21358 29492 21364 29504
rect 20772 29464 21364 29492
rect 20772 29452 20778 29464
rect 21358 29452 21364 29464
rect 21416 29492 21422 29504
rect 21928 29492 21956 29591
rect 22830 29588 22836 29640
rect 22888 29628 22894 29640
rect 23750 29628 23756 29640
rect 22888 29600 23756 29628
rect 22888 29588 22894 29600
rect 23750 29588 23756 29600
rect 23808 29588 23814 29640
rect 23845 29631 23903 29637
rect 23845 29597 23857 29631
rect 23891 29597 23903 29631
rect 23845 29591 23903 29597
rect 24029 29631 24087 29637
rect 24029 29597 24041 29631
rect 24075 29628 24087 29631
rect 24765 29631 24823 29637
rect 24765 29628 24777 29631
rect 24075 29600 24777 29628
rect 24075 29597 24087 29600
rect 24029 29591 24087 29597
rect 24765 29597 24777 29600
rect 24811 29597 24823 29631
rect 25424 29628 25452 29659
rect 46474 29656 46480 29668
rect 46532 29656 46538 29708
rect 46661 29699 46719 29705
rect 46661 29665 46673 29699
rect 46707 29696 46719 29699
rect 47854 29696 47860 29708
rect 46707 29668 47860 29696
rect 46707 29665 46719 29668
rect 46661 29659 46719 29665
rect 47854 29656 47860 29668
rect 47912 29656 47918 29708
rect 27341 29631 27399 29637
rect 27341 29628 27353 29631
rect 25424 29600 27353 29628
rect 24765 29591 24823 29597
rect 27341 29597 27353 29600
rect 27387 29597 27399 29631
rect 27341 29591 27399 29597
rect 23014 29520 23020 29572
rect 23072 29560 23078 29572
rect 23109 29563 23167 29569
rect 23109 29560 23121 29563
rect 23072 29532 23121 29560
rect 23072 29520 23078 29532
rect 23109 29529 23121 29532
rect 23155 29529 23167 29563
rect 23109 29523 23167 29529
rect 23382 29520 23388 29572
rect 23440 29560 23446 29572
rect 23860 29560 23888 29591
rect 24581 29563 24639 29569
rect 24581 29560 24593 29563
rect 23440 29532 24593 29560
rect 23440 29520 23446 29532
rect 24581 29529 24593 29532
rect 24627 29560 24639 29563
rect 24670 29560 24676 29572
rect 24627 29532 24676 29560
rect 24627 29529 24639 29532
rect 24581 29523 24639 29529
rect 24670 29520 24676 29532
rect 24728 29520 24734 29572
rect 24780 29560 24808 29591
rect 28534 29588 28540 29640
rect 28592 29628 28598 29640
rect 29917 29631 29975 29637
rect 29917 29628 29929 29631
rect 28592 29600 29929 29628
rect 28592 29588 28598 29600
rect 29917 29597 29929 29600
rect 29963 29597 29975 29631
rect 29917 29591 29975 29597
rect 25676 29563 25734 29569
rect 24780 29532 25544 29560
rect 21416 29464 21956 29492
rect 21416 29452 21422 29464
rect 23198 29452 23204 29504
rect 23256 29492 23262 29504
rect 23293 29495 23351 29501
rect 23293 29492 23305 29495
rect 23256 29464 23305 29492
rect 23256 29452 23262 29464
rect 23293 29461 23305 29464
rect 23339 29461 23351 29495
rect 23293 29455 23351 29461
rect 23658 29452 23664 29504
rect 23716 29492 23722 29504
rect 23937 29495 23995 29501
rect 23937 29492 23949 29495
rect 23716 29464 23949 29492
rect 23716 29452 23722 29464
rect 23937 29461 23949 29464
rect 23983 29461 23995 29495
rect 24946 29492 24952 29504
rect 24907 29464 24952 29492
rect 23937 29455 23995 29461
rect 24946 29452 24952 29464
rect 25004 29452 25010 29504
rect 25516 29492 25544 29532
rect 25676 29529 25688 29563
rect 25722 29560 25734 29563
rect 26142 29560 26148 29572
rect 25722 29532 26148 29560
rect 25722 29529 25734 29532
rect 25676 29523 25734 29529
rect 26142 29520 26148 29532
rect 26200 29520 26206 29572
rect 27614 29569 27620 29572
rect 27608 29523 27620 29569
rect 27672 29560 27678 29572
rect 29733 29563 29791 29569
rect 29733 29560 29745 29563
rect 27672 29532 27708 29560
rect 28736 29532 29745 29560
rect 27614 29520 27620 29523
rect 27672 29520 27678 29532
rect 26510 29492 26516 29504
rect 25516 29464 26516 29492
rect 26510 29452 26516 29464
rect 26568 29492 26574 29504
rect 26789 29495 26847 29501
rect 26789 29492 26801 29495
rect 26568 29464 26801 29492
rect 26568 29452 26574 29464
rect 26789 29461 26801 29464
rect 26835 29461 26847 29495
rect 26789 29455 26847 29461
rect 27982 29452 27988 29504
rect 28040 29492 28046 29504
rect 28736 29501 28764 29532
rect 29733 29529 29745 29532
rect 29779 29529 29791 29563
rect 48314 29560 48320 29572
rect 48275 29532 48320 29560
rect 29733 29523 29791 29529
rect 48314 29520 48320 29532
rect 48372 29520 48378 29572
rect 28721 29495 28779 29501
rect 28721 29492 28733 29495
rect 28040 29464 28733 29492
rect 28040 29452 28046 29464
rect 28721 29461 28733 29464
rect 28767 29461 28779 29495
rect 28721 29455 28779 29461
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 7282 29288 7288 29300
rect 7243 29260 7288 29288
rect 7282 29248 7288 29260
rect 7340 29248 7346 29300
rect 7653 29291 7711 29297
rect 7653 29257 7665 29291
rect 7699 29288 7711 29291
rect 7834 29288 7840 29300
rect 7699 29260 7840 29288
rect 7699 29257 7711 29260
rect 7653 29251 7711 29257
rect 7834 29248 7840 29260
rect 7892 29248 7898 29300
rect 8662 29288 8668 29300
rect 8623 29260 8668 29288
rect 8662 29248 8668 29260
rect 8720 29248 8726 29300
rect 16574 29248 16580 29300
rect 16632 29288 16638 29300
rect 17053 29291 17111 29297
rect 17053 29288 17065 29291
rect 16632 29260 17065 29288
rect 16632 29248 16638 29260
rect 17053 29257 17065 29260
rect 17099 29257 17111 29291
rect 17053 29251 17111 29257
rect 19058 29248 19064 29300
rect 19116 29288 19122 29300
rect 22830 29288 22836 29300
rect 19116 29260 22836 29288
rect 19116 29248 19122 29260
rect 22830 29248 22836 29260
rect 22888 29248 22894 29300
rect 23581 29260 24624 29288
rect 16117 29223 16175 29229
rect 16117 29189 16129 29223
rect 16163 29220 16175 29223
rect 16666 29220 16672 29232
rect 16163 29192 16672 29220
rect 16163 29189 16175 29192
rect 16117 29183 16175 29189
rect 16666 29180 16672 29192
rect 16724 29220 16730 29232
rect 16853 29223 16911 29229
rect 16853 29220 16865 29223
rect 16724 29192 16865 29220
rect 16724 29180 16730 29192
rect 16853 29189 16865 29192
rect 16899 29189 16911 29223
rect 16853 29183 16911 29189
rect 20714 29180 20720 29232
rect 20772 29220 20778 29232
rect 23581 29229 23609 29260
rect 20993 29223 21051 29229
rect 20993 29220 21005 29223
rect 20772 29192 21005 29220
rect 20772 29180 20778 29192
rect 20993 29189 21005 29192
rect 21039 29189 21051 29223
rect 23569 29223 23627 29229
rect 20993 29183 21051 29189
rect 22204 29192 23520 29220
rect 5166 29152 5172 29164
rect 5127 29124 5172 29152
rect 5166 29112 5172 29124
rect 5224 29112 5230 29164
rect 7466 29152 7472 29164
rect 7427 29124 7472 29152
rect 7466 29112 7472 29124
rect 7524 29112 7530 29164
rect 7745 29155 7803 29161
rect 7745 29121 7757 29155
rect 7791 29121 7803 29155
rect 7745 29115 7803 29121
rect 7760 29084 7788 29115
rect 7834 29112 7840 29164
rect 7892 29152 7898 29164
rect 8205 29155 8263 29161
rect 8205 29152 8217 29155
rect 7892 29124 8217 29152
rect 7892 29112 7898 29124
rect 8205 29121 8217 29124
rect 8251 29121 8263 29155
rect 8205 29115 8263 29121
rect 15378 29112 15384 29164
rect 15436 29152 15442 29164
rect 15930 29152 15936 29164
rect 15436 29124 15936 29152
rect 15436 29112 15442 29124
rect 15930 29112 15936 29124
rect 15988 29112 15994 29164
rect 16022 29112 16028 29164
rect 16080 29152 16086 29164
rect 16209 29155 16267 29161
rect 16209 29152 16221 29155
rect 16080 29124 16221 29152
rect 16080 29112 16086 29124
rect 16209 29121 16221 29124
rect 16255 29121 16267 29155
rect 16209 29115 16267 29121
rect 18506 29112 18512 29164
rect 18564 29152 18570 29164
rect 22204 29152 22232 29192
rect 23492 29164 23520 29192
rect 23569 29189 23581 29223
rect 23615 29189 23627 29223
rect 24394 29220 24400 29232
rect 23569 29183 23627 29189
rect 24320 29192 24400 29220
rect 22370 29152 22376 29164
rect 18564 29124 22232 29152
rect 22331 29124 22376 29152
rect 18564 29112 18570 29124
rect 22370 29112 22376 29124
rect 22428 29112 22434 29164
rect 22646 29152 22652 29164
rect 22607 29124 22652 29152
rect 22646 29112 22652 29124
rect 22704 29112 22710 29164
rect 23198 29152 23204 29164
rect 23159 29124 23204 29152
rect 23198 29112 23204 29124
rect 23256 29112 23262 29164
rect 23382 29161 23388 29164
rect 23349 29155 23388 29161
rect 23349 29121 23361 29155
rect 23349 29115 23388 29121
rect 23382 29112 23388 29115
rect 23440 29112 23446 29164
rect 23474 29112 23480 29164
rect 23532 29152 23538 29164
rect 23750 29161 23756 29164
rect 23707 29155 23756 29161
rect 23532 29124 23577 29152
rect 23532 29112 23538 29124
rect 23707 29121 23719 29155
rect 23753 29121 23756 29155
rect 23707 29115 23756 29121
rect 23750 29112 23756 29115
rect 23808 29112 23814 29164
rect 24320 29161 24348 29192
rect 24394 29180 24400 29192
rect 24452 29180 24458 29232
rect 24596 29220 24624 29260
rect 24670 29248 24676 29300
rect 24728 29288 24734 29300
rect 25685 29291 25743 29297
rect 25685 29288 25697 29291
rect 24728 29260 25697 29288
rect 24728 29248 24734 29260
rect 25685 29257 25697 29260
rect 25731 29257 25743 29291
rect 26142 29288 26148 29300
rect 26103 29260 26148 29288
rect 25685 29251 25743 29257
rect 26142 29248 26148 29260
rect 26200 29248 26206 29300
rect 27982 29288 27988 29300
rect 27943 29260 27988 29288
rect 27982 29248 27988 29260
rect 28040 29248 28046 29300
rect 28077 29291 28135 29297
rect 28077 29257 28089 29291
rect 28123 29288 28135 29291
rect 28813 29291 28871 29297
rect 28813 29288 28825 29291
rect 28123 29260 28825 29288
rect 28123 29257 28135 29260
rect 28077 29251 28135 29257
rect 28813 29257 28825 29260
rect 28859 29257 28871 29291
rect 29270 29288 29276 29300
rect 29231 29260 29276 29288
rect 28813 29251 28871 29257
rect 29270 29248 29276 29260
rect 29328 29248 29334 29300
rect 25038 29220 25044 29232
rect 24596 29192 25044 29220
rect 25038 29180 25044 29192
rect 25096 29180 25102 29232
rect 24305 29155 24363 29161
rect 24305 29121 24317 29155
rect 24351 29121 24363 29155
rect 24561 29155 24619 29161
rect 24561 29152 24573 29155
rect 24305 29115 24363 29121
rect 24412 29124 24573 29152
rect 8386 29084 8392 29096
rect 7760 29056 8392 29084
rect 8386 29044 8392 29056
rect 8444 29084 8450 29096
rect 9214 29084 9220 29096
rect 8444 29056 9220 29084
rect 8444 29044 8450 29056
rect 9214 29044 9220 29056
rect 9272 29044 9278 29096
rect 15749 29087 15807 29093
rect 15749 29053 15761 29087
rect 15795 29084 15807 29087
rect 16942 29084 16948 29096
rect 15795 29056 16948 29084
rect 15795 29053 15807 29056
rect 15749 29047 15807 29053
rect 16942 29044 16948 29056
rect 17000 29044 17006 29096
rect 22465 29087 22523 29093
rect 22465 29053 22477 29087
rect 22511 29053 22523 29087
rect 22465 29047 22523 29053
rect 22557 29087 22615 29093
rect 22557 29053 22569 29087
rect 22603 29053 22615 29087
rect 24412 29084 24440 29124
rect 24561 29121 24573 29124
rect 24607 29121 24619 29155
rect 26326 29152 26332 29164
rect 26287 29124 26332 29152
rect 24561 29115 24619 29121
rect 26326 29112 26332 29124
rect 26384 29112 26390 29164
rect 26513 29155 26571 29161
rect 26513 29121 26525 29155
rect 26559 29152 26571 29155
rect 27522 29152 27528 29164
rect 26559 29124 27528 29152
rect 26559 29121 26571 29124
rect 26513 29115 26571 29121
rect 27522 29112 27528 29124
rect 27580 29152 27586 29164
rect 27890 29152 27896 29164
rect 27580 29124 27896 29152
rect 27580 29112 27586 29124
rect 27890 29112 27896 29124
rect 27948 29112 27954 29164
rect 29178 29152 29184 29164
rect 29139 29124 29184 29152
rect 29178 29112 29184 29124
rect 29236 29112 29242 29164
rect 30834 29152 30840 29164
rect 30795 29124 30840 29152
rect 30834 29112 30840 29124
rect 30892 29112 30898 29164
rect 33410 29152 33416 29164
rect 31726 29124 33416 29152
rect 26605 29087 26663 29093
rect 26605 29084 26617 29087
rect 22557 29047 22615 29053
rect 23860 29056 24440 29084
rect 26252 29056 26617 29084
rect 5718 29016 5724 29028
rect 5460 28988 5724 29016
rect 5460 28957 5488 28988
rect 5718 28976 5724 28988
rect 5776 28976 5782 29028
rect 21266 29016 21272 29028
rect 21227 28988 21272 29016
rect 21266 28976 21272 28988
rect 21324 28976 21330 29028
rect 21453 29019 21511 29025
rect 21453 28985 21465 29019
rect 21499 29016 21511 29019
rect 22094 29016 22100 29028
rect 21499 28988 22100 29016
rect 21499 28985 21511 28988
rect 21453 28979 21511 28985
rect 22094 28976 22100 28988
rect 22152 29016 22158 29028
rect 22480 29016 22508 29047
rect 22152 28988 22508 29016
rect 22572 29016 22600 29047
rect 23658 29016 23664 29028
rect 22572 28988 23664 29016
rect 22152 28976 22158 28988
rect 23658 28976 23664 28988
rect 23716 28976 23722 29028
rect 23860 29025 23888 29056
rect 23845 29019 23903 29025
rect 23845 28985 23857 29019
rect 23891 28985 23903 29019
rect 23845 28979 23903 28985
rect 5445 28951 5503 28957
rect 5445 28917 5457 28951
rect 5491 28917 5503 28951
rect 5626 28948 5632 28960
rect 5587 28920 5632 28948
rect 5445 28911 5503 28917
rect 5626 28908 5632 28920
rect 5684 28908 5690 28960
rect 8294 28948 8300 28960
rect 8255 28920 8300 28948
rect 8294 28908 8300 28920
rect 8352 28908 8358 28960
rect 16942 28908 16948 28960
rect 17000 28948 17006 28960
rect 17037 28951 17095 28957
rect 17037 28948 17049 28951
rect 17000 28920 17049 28948
rect 17000 28908 17006 28920
rect 17037 28917 17049 28920
rect 17083 28917 17095 28951
rect 17218 28948 17224 28960
rect 17179 28920 17224 28948
rect 17037 28911 17095 28917
rect 17218 28908 17224 28920
rect 17276 28908 17282 28960
rect 22189 28951 22247 28957
rect 22189 28917 22201 28951
rect 22235 28948 22247 28951
rect 22370 28948 22376 28960
rect 22235 28920 22376 28948
rect 22235 28917 22247 28920
rect 22189 28911 22247 28917
rect 22370 28908 22376 28920
rect 22428 28908 22434 28960
rect 25406 28908 25412 28960
rect 25464 28948 25470 28960
rect 26252 28948 26280 29056
rect 26605 29053 26617 29056
rect 26651 29053 26663 29087
rect 26605 29047 26663 29053
rect 28166 29044 28172 29096
rect 28224 29084 28230 29096
rect 29365 29087 29423 29093
rect 28224 29056 28269 29084
rect 28224 29044 28230 29056
rect 29365 29053 29377 29087
rect 29411 29053 29423 29087
rect 29365 29047 29423 29053
rect 29380 29016 29408 29047
rect 30650 29044 30656 29096
rect 30708 29084 30714 29096
rect 31113 29087 31171 29093
rect 31113 29084 31125 29087
rect 30708 29056 31125 29084
rect 30708 29044 30714 29056
rect 31113 29053 31125 29056
rect 31159 29084 31171 29087
rect 31726 29084 31754 29124
rect 33410 29112 33416 29124
rect 33468 29152 33474 29164
rect 38010 29152 38016 29164
rect 33468 29124 38016 29152
rect 33468 29112 33474 29124
rect 38010 29112 38016 29124
rect 38068 29112 38074 29164
rect 47670 29112 47676 29164
rect 47728 29152 47734 29164
rect 47765 29155 47823 29161
rect 47765 29152 47777 29155
rect 47728 29124 47777 29152
rect 47728 29112 47734 29124
rect 47765 29121 47777 29124
rect 47811 29121 47823 29155
rect 47765 29115 47823 29121
rect 31159 29056 31754 29084
rect 31159 29053 31171 29056
rect 31113 29047 31171 29053
rect 31018 29016 31024 29028
rect 27540 28988 29408 29016
rect 30979 28988 31024 29016
rect 25464 28920 26280 28948
rect 25464 28908 25470 28920
rect 26694 28908 26700 28960
rect 26752 28948 26758 28960
rect 27540 28948 27568 28988
rect 31018 28976 31024 28988
rect 31076 28976 31082 29028
rect 31846 28976 31852 29028
rect 31904 29016 31910 29028
rect 38470 29016 38476 29028
rect 31904 28988 38476 29016
rect 31904 28976 31910 28988
rect 38470 28976 38476 28988
rect 38528 28976 38534 29028
rect 26752 28920 27568 28948
rect 27617 28951 27675 28957
rect 26752 28908 26758 28920
rect 27617 28917 27629 28951
rect 27663 28948 27675 28951
rect 27706 28948 27712 28960
rect 27663 28920 27712 28948
rect 27663 28917 27675 28920
rect 27617 28911 27675 28917
rect 27706 28908 27712 28920
rect 27764 28908 27770 28960
rect 30650 28948 30656 28960
rect 30611 28920 30656 28948
rect 30650 28908 30656 28920
rect 30708 28908 30714 28960
rect 47210 28948 47216 28960
rect 47171 28920 47216 28948
rect 47210 28908 47216 28920
rect 47268 28908 47274 28960
rect 47854 28948 47860 28960
rect 47815 28920 47860 28948
rect 47854 28908 47860 28920
rect 47912 28908 47918 28960
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 9214 28744 9220 28756
rect 9175 28716 9220 28744
rect 9214 28704 9220 28716
rect 9272 28704 9278 28756
rect 13814 28704 13820 28756
rect 13872 28744 13878 28756
rect 14458 28744 14464 28756
rect 13872 28716 14464 28744
rect 13872 28704 13878 28716
rect 14458 28704 14464 28716
rect 14516 28744 14522 28756
rect 23566 28744 23572 28756
rect 14516 28716 21036 28744
rect 23527 28716 23572 28744
rect 14516 28704 14522 28716
rect 14550 28568 14556 28620
rect 14608 28608 14614 28620
rect 21008 28617 21036 28716
rect 23566 28704 23572 28716
rect 23624 28704 23630 28756
rect 27525 28747 27583 28753
rect 27525 28713 27537 28747
rect 27571 28744 27583 28747
rect 27614 28744 27620 28756
rect 27571 28716 27620 28744
rect 27571 28713 27583 28716
rect 27525 28707 27583 28713
rect 27614 28704 27620 28716
rect 27672 28704 27678 28756
rect 28074 28704 28080 28756
rect 28132 28744 28138 28756
rect 28445 28747 28503 28753
rect 28445 28744 28457 28747
rect 28132 28716 28457 28744
rect 28132 28704 28138 28716
rect 28445 28713 28457 28716
rect 28491 28713 28503 28747
rect 32122 28744 32128 28756
rect 32083 28716 32128 28744
rect 28445 28707 28503 28713
rect 32122 28704 32128 28716
rect 32180 28704 32186 28756
rect 15473 28611 15531 28617
rect 15473 28608 15485 28611
rect 14608 28580 15485 28608
rect 14608 28568 14614 28580
rect 15473 28577 15485 28580
rect 15519 28577 15531 28611
rect 15473 28571 15531 28577
rect 15657 28611 15715 28617
rect 15657 28577 15669 28611
rect 15703 28608 15715 28611
rect 20993 28611 21051 28617
rect 15703 28580 17632 28608
rect 15703 28577 15715 28580
rect 15657 28571 15715 28577
rect 5169 28543 5227 28549
rect 5169 28509 5181 28543
rect 5215 28540 5227 28543
rect 5626 28540 5632 28552
rect 5215 28512 5632 28540
rect 5215 28509 5227 28512
rect 5169 28503 5227 28509
rect 5626 28500 5632 28512
rect 5684 28500 5690 28552
rect 9125 28543 9183 28549
rect 9125 28509 9137 28543
rect 9171 28540 9183 28543
rect 9398 28540 9404 28552
rect 9171 28512 9404 28540
rect 9171 28509 9183 28512
rect 9125 28503 9183 28509
rect 9398 28500 9404 28512
rect 9456 28500 9462 28552
rect 13446 28540 13452 28552
rect 13407 28512 13452 28540
rect 13446 28500 13452 28512
rect 13504 28500 13510 28552
rect 13630 28540 13636 28552
rect 13591 28512 13636 28540
rect 13630 28500 13636 28512
rect 13688 28500 13694 28552
rect 15381 28543 15439 28549
rect 15381 28509 15393 28543
rect 15427 28509 15439 28543
rect 15381 28503 15439 28509
rect 15565 28543 15623 28549
rect 15565 28509 15577 28543
rect 15611 28540 15623 28543
rect 15746 28540 15752 28552
rect 15611 28512 15752 28540
rect 15611 28509 15623 28512
rect 15565 28503 15623 28509
rect 14826 28432 14832 28484
rect 14884 28472 14890 28484
rect 15396 28472 15424 28503
rect 15746 28500 15752 28512
rect 15804 28500 15810 28552
rect 15838 28500 15844 28552
rect 15896 28540 15902 28552
rect 16393 28543 16451 28549
rect 15896 28512 16335 28540
rect 15896 28500 15902 28512
rect 16307 28472 16335 28512
rect 16393 28509 16405 28543
rect 16439 28540 16451 28543
rect 16574 28540 16580 28552
rect 16439 28512 16580 28540
rect 16439 28509 16451 28512
rect 16393 28503 16451 28509
rect 16574 28500 16580 28512
rect 16632 28500 16638 28552
rect 16669 28543 16727 28549
rect 16669 28509 16681 28543
rect 16715 28540 16727 28543
rect 16942 28540 16948 28552
rect 16715 28512 16948 28540
rect 16715 28509 16727 28512
rect 16669 28503 16727 28509
rect 16684 28472 16712 28503
rect 16942 28500 16948 28512
rect 17000 28500 17006 28552
rect 17402 28500 17408 28552
rect 17460 28540 17466 28552
rect 17497 28543 17555 28549
rect 17497 28540 17509 28543
rect 17460 28512 17509 28540
rect 17460 28500 17466 28512
rect 17497 28509 17509 28512
rect 17543 28509 17555 28543
rect 17604 28540 17632 28580
rect 20993 28577 21005 28611
rect 21039 28577 21051 28611
rect 22646 28608 22652 28620
rect 20993 28571 21051 28577
rect 21100 28580 22652 28608
rect 21100 28540 21128 28580
rect 22646 28568 22652 28580
rect 22704 28568 22710 28620
rect 24946 28608 24952 28620
rect 23492 28580 24952 28608
rect 17604 28512 21128 28540
rect 17497 28503 17555 28509
rect 22094 28500 22100 28552
rect 22152 28540 22158 28552
rect 22152 28512 22197 28540
rect 22152 28500 22158 28512
rect 22278 28500 22284 28552
rect 22336 28540 22342 28552
rect 23492 28549 23520 28580
rect 24946 28568 24952 28580
rect 25004 28568 25010 28620
rect 27154 28568 27160 28620
rect 27212 28608 27218 28620
rect 30745 28611 30803 28617
rect 30745 28608 30757 28611
rect 27212 28580 30757 28608
rect 27212 28568 27218 28580
rect 30745 28577 30757 28580
rect 30791 28577 30803 28611
rect 30745 28571 30803 28577
rect 46477 28611 46535 28617
rect 46477 28577 46489 28611
rect 46523 28608 46535 28611
rect 47210 28608 47216 28620
rect 46523 28580 47216 28608
rect 46523 28577 46535 28580
rect 46477 28571 46535 28577
rect 47210 28568 47216 28580
rect 47268 28568 47274 28620
rect 48222 28608 48228 28620
rect 48183 28580 48228 28608
rect 48222 28568 48228 28580
rect 48280 28568 48286 28620
rect 22373 28543 22431 28549
rect 22373 28540 22385 28543
rect 22336 28512 22385 28540
rect 22336 28500 22342 28512
rect 22373 28509 22385 28512
rect 22419 28509 22431 28543
rect 22373 28503 22431 28509
rect 23477 28543 23535 28549
rect 23477 28509 23489 28543
rect 23523 28509 23535 28543
rect 23658 28540 23664 28552
rect 23619 28512 23664 28540
rect 23477 28503 23535 28509
rect 23658 28500 23664 28512
rect 23716 28500 23722 28552
rect 27706 28540 27712 28552
rect 27667 28512 27712 28540
rect 27706 28500 27712 28512
rect 27764 28500 27770 28552
rect 27982 28500 27988 28552
rect 28040 28540 28046 28552
rect 28353 28543 28411 28549
rect 28353 28540 28365 28543
rect 28040 28512 28365 28540
rect 28040 28500 28046 28512
rect 28353 28509 28365 28512
rect 28399 28509 28411 28543
rect 28534 28540 28540 28552
rect 28495 28512 28540 28540
rect 28353 28503 28411 28509
rect 28534 28500 28540 28512
rect 28592 28500 28598 28552
rect 30650 28500 30656 28552
rect 30708 28540 30714 28552
rect 31001 28543 31059 28549
rect 31001 28540 31013 28543
rect 30708 28512 31013 28540
rect 30708 28500 30714 28512
rect 31001 28509 31013 28512
rect 31047 28509 31059 28543
rect 31001 28503 31059 28509
rect 35894 28500 35900 28552
rect 35952 28540 35958 28552
rect 36541 28543 36599 28549
rect 36541 28540 36553 28543
rect 35952 28512 36553 28540
rect 35952 28500 35958 28512
rect 36541 28509 36553 28512
rect 36587 28509 36599 28543
rect 36541 28503 36599 28509
rect 14884 28444 16252 28472
rect 16307 28444 16712 28472
rect 17764 28475 17822 28481
rect 14884 28432 14890 28444
rect 16224 28416 16252 28444
rect 17764 28441 17776 28475
rect 17810 28472 17822 28475
rect 18782 28472 18788 28484
rect 17810 28444 18788 28472
rect 17810 28441 17822 28444
rect 17764 28435 17822 28441
rect 18782 28432 18788 28444
rect 18840 28432 18846 28484
rect 23676 28472 23704 28500
rect 22296 28444 23704 28472
rect 37369 28475 37427 28481
rect 4982 28404 4988 28416
rect 4943 28376 4988 28404
rect 4982 28364 4988 28376
rect 5040 28364 5046 28416
rect 13538 28404 13544 28416
rect 13499 28376 13544 28404
rect 13538 28364 13544 28376
rect 13596 28364 13602 28416
rect 15194 28404 15200 28416
rect 15155 28376 15200 28404
rect 15194 28364 15200 28376
rect 15252 28364 15258 28416
rect 16206 28404 16212 28416
rect 16167 28376 16212 28404
rect 16206 28364 16212 28376
rect 16264 28364 16270 28416
rect 16577 28407 16635 28413
rect 16577 28373 16589 28407
rect 16623 28404 16635 28407
rect 16666 28404 16672 28416
rect 16623 28376 16672 28404
rect 16623 28373 16635 28376
rect 16577 28367 16635 28373
rect 16666 28364 16672 28376
rect 16724 28364 16730 28416
rect 17494 28364 17500 28416
rect 17552 28404 17558 28416
rect 18414 28404 18420 28416
rect 17552 28376 18420 28404
rect 17552 28364 17558 28376
rect 18414 28364 18420 28376
rect 18472 28404 18478 28416
rect 18877 28407 18935 28413
rect 18877 28404 18889 28407
rect 18472 28376 18889 28404
rect 18472 28364 18478 28376
rect 18877 28373 18889 28376
rect 18923 28373 18935 28407
rect 18877 28367 18935 28373
rect 20162 28364 20168 28416
rect 20220 28404 20226 28416
rect 20441 28407 20499 28413
rect 20441 28404 20453 28407
rect 20220 28376 20453 28404
rect 20220 28364 20226 28376
rect 20441 28373 20453 28376
rect 20487 28373 20499 28407
rect 20806 28404 20812 28416
rect 20767 28376 20812 28404
rect 20441 28367 20499 28373
rect 20806 28364 20812 28376
rect 20864 28364 20870 28416
rect 20898 28364 20904 28416
rect 20956 28404 20962 28416
rect 22186 28404 22192 28416
rect 22244 28413 22250 28416
rect 22296 28413 22324 28444
rect 37369 28441 37381 28475
rect 37415 28472 37427 28475
rect 38102 28472 38108 28484
rect 37415 28444 38108 28472
rect 37415 28441 37427 28444
rect 37369 28435 37427 28441
rect 38102 28432 38108 28444
rect 38160 28432 38166 28484
rect 46661 28475 46719 28481
rect 46661 28441 46673 28475
rect 46707 28472 46719 28475
rect 47854 28472 47860 28484
rect 46707 28444 47860 28472
rect 46707 28441 46719 28444
rect 46661 28435 46719 28441
rect 47854 28432 47860 28444
rect 47912 28432 47918 28484
rect 20956 28376 21001 28404
rect 22153 28376 22192 28404
rect 20956 28364 20962 28376
rect 22186 28364 22192 28376
rect 22244 28367 22253 28413
rect 22281 28407 22339 28413
rect 22281 28373 22293 28407
rect 22327 28373 22339 28407
rect 22281 28367 22339 28373
rect 22244 28364 22250 28367
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 4706 28200 4712 28212
rect 4540 28172 4712 28200
rect 4341 28067 4399 28073
rect 4341 28033 4353 28067
rect 4387 28064 4399 28067
rect 4540 28064 4568 28172
rect 4706 28160 4712 28172
rect 4764 28160 4770 28212
rect 13357 28203 13415 28209
rect 13357 28169 13369 28203
rect 13403 28200 13415 28203
rect 13446 28200 13452 28212
rect 13403 28172 13452 28200
rect 13403 28169 13415 28172
rect 13357 28163 13415 28169
rect 13446 28160 13452 28172
rect 13504 28160 13510 28212
rect 15289 28203 15347 28209
rect 15289 28169 15301 28203
rect 15335 28200 15347 28203
rect 16022 28200 16028 28212
rect 15335 28172 16028 28200
rect 15335 28169 15347 28172
rect 15289 28163 15347 28169
rect 16022 28160 16028 28172
rect 16080 28160 16086 28212
rect 17589 28203 17647 28209
rect 17589 28169 17601 28203
rect 17635 28200 17647 28203
rect 17635 28172 18276 28200
rect 17635 28169 17647 28172
rect 17589 28163 17647 28169
rect 4608 28135 4666 28141
rect 4608 28101 4620 28135
rect 4654 28132 4666 28135
rect 4982 28132 4988 28144
rect 4654 28104 4988 28132
rect 4654 28101 4666 28104
rect 4608 28095 4666 28101
rect 4982 28092 4988 28104
rect 5040 28092 5046 28144
rect 6914 28092 6920 28144
rect 6972 28132 6978 28144
rect 7929 28135 7987 28141
rect 7929 28132 7941 28135
rect 6972 28104 7941 28132
rect 6972 28092 6978 28104
rect 7929 28101 7941 28104
rect 7975 28101 7987 28135
rect 14550 28132 14556 28144
rect 14511 28104 14556 28132
rect 7929 28095 7987 28101
rect 14550 28092 14556 28104
rect 14608 28092 14614 28144
rect 15470 28092 15476 28144
rect 15528 28132 15534 28144
rect 17405 28135 17463 28141
rect 15528 28104 15608 28132
rect 15528 28092 15534 28104
rect 4387 28036 4568 28064
rect 8941 28067 8999 28073
rect 4387 28033 4399 28036
rect 4341 28027 4399 28033
rect 8941 28033 8953 28067
rect 8987 28064 8999 28067
rect 9398 28064 9404 28076
rect 8987 28036 9404 28064
rect 8987 28033 8999 28036
rect 8941 28027 8999 28033
rect 9398 28024 9404 28036
rect 9456 28024 9462 28076
rect 12802 28024 12808 28076
rect 12860 28064 12866 28076
rect 12986 28064 12992 28076
rect 12860 28036 12992 28064
rect 12860 28024 12866 28036
rect 12986 28024 12992 28036
rect 13044 28024 13050 28076
rect 13449 28067 13507 28073
rect 13449 28033 13461 28067
rect 13495 28064 13507 28067
rect 14366 28064 14372 28076
rect 13495 28036 14372 28064
rect 13495 28033 13507 28036
rect 13449 28027 13507 28033
rect 14366 28024 14372 28036
rect 14424 28024 14430 28076
rect 14737 28067 14795 28073
rect 14737 28033 14749 28067
rect 14783 28033 14795 28067
rect 14737 28027 14795 28033
rect 8846 27996 8852 28008
rect 8807 27968 8852 27996
rect 8846 27956 8852 27968
rect 8904 27956 8910 28008
rect 13633 27999 13691 28005
rect 13633 27965 13645 27999
rect 13679 27996 13691 27999
rect 13814 27996 13820 28008
rect 13679 27968 13820 27996
rect 13679 27965 13691 27968
rect 13633 27959 13691 27965
rect 13814 27956 13820 27968
rect 13872 27956 13878 28008
rect 14752 27996 14780 28027
rect 14826 28024 14832 28076
rect 14884 28064 14890 28076
rect 15580 28073 15608 28104
rect 17405 28101 17417 28135
rect 17451 28132 17463 28135
rect 17954 28132 17960 28144
rect 17451 28104 17960 28132
rect 17451 28101 17463 28104
rect 17405 28095 17463 28101
rect 17954 28092 17960 28104
rect 18012 28092 18018 28144
rect 15565 28067 15623 28073
rect 14884 28036 14929 28064
rect 14884 28024 14890 28036
rect 15565 28033 15577 28067
rect 15611 28033 15623 28067
rect 15565 28027 15623 28033
rect 15654 28067 15712 28073
rect 15654 28033 15666 28067
rect 15700 28033 15712 28067
rect 15654 28027 15712 28033
rect 15749 28070 15807 28076
rect 15749 28036 15761 28070
rect 15795 28036 15807 28070
rect 15749 28030 15807 28036
rect 15933 28067 15991 28073
rect 15933 28033 15945 28067
rect 15979 28033 15991 28067
rect 14752 27968 14872 27996
rect 9309 27931 9367 27937
rect 9309 27897 9321 27931
rect 9355 27928 9367 27931
rect 9582 27928 9588 27940
rect 9355 27900 9588 27928
rect 9355 27897 9367 27900
rect 9309 27891 9367 27897
rect 9582 27888 9588 27900
rect 9640 27888 9646 27940
rect 14844 27928 14872 27968
rect 15672 27928 15700 28027
rect 15764 27996 15792 28030
rect 15933 28027 15991 28033
rect 17037 28067 17095 28073
rect 17037 28033 17049 28067
rect 17083 28064 17095 28067
rect 17218 28064 17224 28076
rect 17083 28036 17224 28064
rect 17083 28033 17095 28036
rect 17037 28027 17095 28033
rect 15838 27996 15844 28008
rect 15764 27968 15844 27996
rect 15838 27956 15844 27968
rect 15896 27956 15902 28008
rect 15746 27928 15752 27940
rect 14844 27900 15752 27928
rect 15746 27888 15752 27900
rect 15804 27888 15810 27940
rect 4982 27820 4988 27872
rect 5040 27860 5046 27872
rect 5721 27863 5779 27869
rect 5721 27860 5733 27863
rect 5040 27832 5733 27860
rect 5040 27820 5046 27832
rect 5721 27829 5733 27832
rect 5767 27829 5779 27863
rect 8018 27860 8024 27872
rect 7979 27832 8024 27860
rect 5721 27823 5779 27829
rect 8018 27820 8024 27832
rect 8076 27820 8082 27872
rect 12710 27820 12716 27872
rect 12768 27860 12774 27872
rect 12989 27863 13047 27869
rect 12989 27860 13001 27863
rect 12768 27832 13001 27860
rect 12768 27820 12774 27832
rect 12989 27829 13001 27832
rect 13035 27829 13047 27863
rect 14550 27860 14556 27872
rect 14511 27832 14556 27860
rect 12989 27823 13047 27829
rect 14550 27820 14556 27832
rect 14608 27820 14614 27872
rect 15562 27820 15568 27872
rect 15620 27860 15626 27872
rect 15948 27860 15976 28027
rect 17218 28024 17224 28036
rect 17276 28024 17282 28076
rect 18248 28073 18276 28172
rect 18782 28160 18788 28212
rect 18840 28200 18846 28212
rect 18877 28203 18935 28209
rect 18877 28200 18889 28203
rect 18840 28172 18889 28200
rect 18840 28160 18846 28172
rect 18877 28169 18889 28172
rect 18923 28169 18935 28203
rect 20806 28200 20812 28212
rect 20767 28172 20812 28200
rect 18877 28163 18935 28169
rect 20806 28160 20812 28172
rect 20864 28160 20870 28212
rect 20898 28160 20904 28212
rect 20956 28200 20962 28212
rect 22097 28203 22155 28209
rect 22097 28200 22109 28203
rect 20956 28172 22109 28200
rect 20956 28160 20962 28172
rect 22097 28169 22109 28172
rect 22143 28169 22155 28203
rect 22097 28163 22155 28169
rect 30653 28203 30711 28209
rect 30653 28169 30665 28203
rect 30699 28200 30711 28203
rect 30834 28200 30840 28212
rect 30699 28172 30840 28200
rect 30699 28169 30711 28172
rect 30653 28163 30711 28169
rect 30834 28160 30840 28172
rect 30892 28160 30898 28212
rect 18506 28132 18512 28144
rect 18467 28104 18512 28132
rect 18506 28092 18512 28104
rect 18564 28092 18570 28144
rect 18601 28135 18659 28141
rect 18601 28101 18613 28135
rect 18647 28132 18659 28135
rect 18647 28104 20760 28132
rect 18647 28101 18659 28104
rect 18601 28095 18659 28101
rect 18414 28073 18420 28076
rect 18233 28067 18291 28073
rect 18233 28033 18245 28067
rect 18279 28033 18291 28067
rect 18233 28027 18291 28033
rect 18381 28067 18420 28073
rect 18381 28033 18393 28067
rect 18381 28027 18420 28033
rect 18414 28024 18420 28027
rect 18472 28024 18478 28076
rect 18739 28067 18797 28073
rect 18739 28033 18751 28067
rect 18785 28064 18797 28067
rect 19058 28064 19064 28076
rect 18785 28036 19064 28064
rect 18785 28033 18797 28036
rect 18739 28027 18797 28033
rect 19058 28024 19064 28036
rect 19116 28024 19122 28076
rect 19696 28067 19754 28073
rect 19696 28033 19708 28067
rect 19742 28064 19754 28067
rect 19978 28064 19984 28076
rect 19742 28036 19984 28064
rect 19742 28033 19754 28036
rect 19696 28027 19754 28033
rect 19978 28024 19984 28036
rect 20036 28024 20042 28076
rect 17402 27956 17408 28008
rect 17460 27996 17466 28008
rect 19426 27996 19432 28008
rect 17460 27968 19432 27996
rect 17460 27956 17466 27968
rect 19426 27956 19432 27968
rect 19484 27956 19490 28008
rect 20732 27996 20760 28104
rect 20824 28064 20852 28160
rect 21358 28132 21364 28144
rect 21319 28104 21364 28132
rect 21358 28092 21364 28104
rect 21416 28092 21422 28144
rect 30742 28092 30748 28144
rect 30800 28132 30806 28144
rect 30800 28104 31156 28132
rect 30800 28092 30806 28104
rect 21269 28067 21327 28073
rect 21269 28064 21281 28067
rect 20824 28036 21281 28064
rect 21269 28033 21281 28036
rect 21315 28033 21327 28067
rect 21450 28064 21456 28076
rect 21411 28036 21456 28064
rect 21269 28027 21327 28033
rect 21450 28024 21456 28036
rect 21508 28024 21514 28076
rect 22186 28024 22192 28076
rect 22244 28064 22250 28076
rect 22281 28067 22339 28073
rect 22281 28064 22293 28067
rect 22244 28036 22293 28064
rect 22244 28024 22250 28036
rect 22281 28033 22293 28036
rect 22327 28033 22339 28067
rect 22281 28027 22339 28033
rect 22370 28024 22376 28076
rect 22428 28064 22434 28076
rect 22646 28064 22652 28076
rect 22428 28036 22473 28064
rect 22607 28036 22652 28064
rect 22428 28024 22434 28036
rect 22646 28024 22652 28036
rect 22704 28024 22710 28076
rect 24578 28064 24584 28076
rect 24539 28036 24584 28064
rect 24578 28024 24584 28036
rect 24636 28024 24642 28076
rect 26694 28064 26700 28076
rect 24780 28036 26700 28064
rect 21358 27996 21364 28008
rect 20732 27968 21364 27996
rect 21358 27956 21364 27968
rect 21416 27956 21422 28008
rect 22554 27996 22560 28008
rect 22467 27968 22560 27996
rect 22554 27956 22560 27968
rect 22612 27996 22618 28008
rect 24780 27996 24808 28036
rect 26694 28024 26700 28036
rect 26752 28024 26758 28076
rect 30466 28024 30472 28076
rect 30524 28064 30530 28076
rect 31128 28073 31156 28104
rect 30837 28067 30895 28073
rect 30837 28064 30849 28067
rect 30524 28036 30849 28064
rect 30524 28024 30530 28036
rect 30837 28033 30849 28036
rect 30883 28033 30895 28067
rect 30837 28027 30895 28033
rect 31113 28067 31171 28073
rect 31113 28033 31125 28067
rect 31159 28033 31171 28067
rect 31113 28027 31171 28033
rect 31297 28067 31355 28073
rect 31297 28033 31309 28067
rect 31343 28064 31355 28067
rect 32122 28064 32128 28076
rect 31343 28036 32128 28064
rect 31343 28033 31355 28036
rect 31297 28027 31355 28033
rect 32122 28024 32128 28036
rect 32180 28024 32186 28076
rect 47486 28024 47492 28076
rect 47544 28064 47550 28076
rect 47762 28064 47768 28076
rect 47544 28036 47768 28064
rect 47544 28024 47550 28036
rect 47762 28024 47768 28036
rect 47820 28024 47826 28076
rect 22612 27968 24808 27996
rect 24857 27999 24915 28005
rect 22612 27956 22618 27968
rect 24857 27965 24869 27999
rect 24903 27996 24915 27999
rect 25406 27996 25412 28008
rect 24903 27968 25412 27996
rect 24903 27965 24915 27968
rect 24857 27959 24915 27965
rect 25406 27956 25412 27968
rect 25464 27956 25470 28008
rect 24397 27931 24455 27937
rect 24397 27897 24409 27931
rect 24443 27928 24455 27931
rect 24443 27900 24900 27928
rect 24443 27897 24455 27900
rect 24397 27891 24455 27897
rect 24872 27872 24900 27900
rect 15620 27832 15976 27860
rect 15620 27820 15626 27832
rect 16206 27820 16212 27872
rect 16264 27860 16270 27872
rect 17405 27863 17463 27869
rect 17405 27860 17417 27863
rect 16264 27832 17417 27860
rect 16264 27820 16270 27832
rect 17405 27829 17417 27832
rect 17451 27829 17463 27863
rect 24762 27860 24768 27872
rect 24723 27832 24768 27860
rect 17405 27823 17463 27829
rect 24762 27820 24768 27832
rect 24820 27820 24826 27872
rect 24854 27820 24860 27872
rect 24912 27820 24918 27872
rect 47210 27860 47216 27872
rect 47171 27832 47216 27860
rect 47210 27820 47216 27832
rect 47268 27820 47274 27872
rect 47854 27860 47860 27872
rect 47815 27832 47860 27860
rect 47854 27820 47860 27832
rect 47912 27820 47918 27872
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 4801 27659 4859 27665
rect 4801 27625 4813 27659
rect 4847 27656 4859 27659
rect 4982 27656 4988 27668
rect 4847 27628 4988 27656
rect 4847 27625 4859 27628
rect 4801 27619 4859 27625
rect 4982 27616 4988 27628
rect 5040 27616 5046 27668
rect 5718 27656 5724 27668
rect 5679 27628 5724 27656
rect 5718 27616 5724 27628
rect 5776 27616 5782 27668
rect 8386 27656 8392 27668
rect 8347 27628 8392 27656
rect 8386 27616 8392 27628
rect 8444 27616 8450 27668
rect 19978 27656 19984 27668
rect 16500 27628 18276 27656
rect 19939 27628 19984 27656
rect 14366 27588 14372 27600
rect 14327 27560 14372 27588
rect 14366 27548 14372 27560
rect 14424 27548 14430 27600
rect 15378 27588 15384 27600
rect 15339 27560 15384 27588
rect 15378 27548 15384 27560
rect 15436 27548 15442 27600
rect 16114 27588 16120 27600
rect 15672 27560 16120 27588
rect 4985 27523 5043 27529
rect 4985 27489 4997 27523
rect 5031 27520 5043 27523
rect 5031 27492 6592 27520
rect 5031 27489 5043 27492
rect 4985 27483 5043 27489
rect 4525 27455 4583 27461
rect 4525 27421 4537 27455
rect 4571 27452 4583 27455
rect 5166 27452 5172 27464
rect 4571 27424 5172 27452
rect 4571 27421 4583 27424
rect 4525 27415 4583 27421
rect 5166 27412 5172 27424
rect 5224 27452 5230 27464
rect 6564 27461 6592 27492
rect 11974 27480 11980 27532
rect 12032 27520 12038 27532
rect 12069 27523 12127 27529
rect 12069 27520 12081 27523
rect 12032 27492 12081 27520
rect 12032 27480 12038 27492
rect 12069 27489 12081 27492
rect 12115 27489 12127 27523
rect 12069 27483 12127 27489
rect 14829 27523 14887 27529
rect 14829 27489 14841 27523
rect 14875 27520 14887 27523
rect 15672 27520 15700 27560
rect 16114 27548 16120 27560
rect 16172 27588 16178 27600
rect 16500 27588 16528 27628
rect 16172 27560 16528 27588
rect 16172 27548 16178 27560
rect 16574 27548 16580 27600
rect 16632 27588 16638 27600
rect 18141 27591 18199 27597
rect 18141 27588 18153 27591
rect 16632 27560 18153 27588
rect 16632 27548 16638 27560
rect 18141 27557 18153 27560
rect 18187 27557 18199 27591
rect 18141 27551 18199 27557
rect 14875 27492 15700 27520
rect 15749 27523 15807 27529
rect 14875 27489 14887 27492
rect 14829 27483 14887 27489
rect 15749 27489 15761 27523
rect 15795 27520 15807 27523
rect 16850 27520 16856 27532
rect 15795 27492 16856 27520
rect 15795 27489 15807 27492
rect 15749 27483 15807 27489
rect 16850 27480 16856 27492
rect 16908 27480 16914 27532
rect 16945 27523 17003 27529
rect 16945 27489 16957 27523
rect 16991 27520 17003 27523
rect 18248 27520 18276 27628
rect 19978 27616 19984 27628
rect 20036 27616 20042 27668
rect 20993 27591 21051 27597
rect 20993 27557 21005 27591
rect 21039 27588 21051 27591
rect 21266 27588 21272 27600
rect 21039 27560 21272 27588
rect 21039 27557 21051 27560
rect 20993 27551 21051 27557
rect 21266 27548 21272 27560
rect 21324 27548 21330 27600
rect 26602 27588 26608 27600
rect 26563 27560 26608 27588
rect 26602 27548 26608 27560
rect 26660 27548 26666 27600
rect 29089 27591 29147 27597
rect 29089 27557 29101 27591
rect 29135 27588 29147 27591
rect 29362 27588 29368 27600
rect 29135 27560 29368 27588
rect 29135 27557 29147 27560
rect 29089 27551 29147 27557
rect 29362 27548 29368 27560
rect 29420 27548 29426 27600
rect 22554 27520 22560 27532
rect 16991 27492 18092 27520
rect 18248 27492 22560 27520
rect 16991 27489 17003 27492
rect 16945 27483 17003 27489
rect 5445 27455 5503 27461
rect 5445 27452 5457 27455
rect 5224 27424 5457 27452
rect 5224 27412 5230 27424
rect 5445 27421 5457 27424
rect 5491 27421 5503 27455
rect 5445 27415 5503 27421
rect 6549 27455 6607 27461
rect 6549 27421 6561 27455
rect 6595 27421 6607 27455
rect 6549 27415 6607 27421
rect 8113 27455 8171 27461
rect 8113 27421 8125 27455
rect 8159 27421 8171 27455
rect 14550 27452 14556 27464
rect 14511 27424 14556 27452
rect 8113 27415 8171 27421
rect 5460 27384 5488 27415
rect 7006 27384 7012 27396
rect 5460 27356 7012 27384
rect 7006 27344 7012 27356
rect 7064 27384 7070 27396
rect 8128 27384 8156 27415
rect 14550 27412 14556 27424
rect 14608 27412 14614 27464
rect 14645 27455 14703 27461
rect 14645 27421 14657 27455
rect 14691 27421 14703 27455
rect 14645 27415 14703 27421
rect 14921 27455 14979 27461
rect 14921 27421 14933 27455
rect 14967 27452 14979 27455
rect 15286 27452 15292 27464
rect 14967 27424 15292 27452
rect 14967 27421 14979 27424
rect 14921 27415 14979 27421
rect 7064 27356 8156 27384
rect 12336 27387 12394 27393
rect 7064 27344 7070 27356
rect 12336 27353 12348 27387
rect 12382 27384 12394 27387
rect 12526 27384 12532 27396
rect 12382 27356 12532 27384
rect 12382 27353 12394 27356
rect 12336 27347 12394 27353
rect 12526 27344 12532 27356
rect 12584 27344 12590 27396
rect 14660 27384 14688 27415
rect 15286 27412 15292 27424
rect 15344 27412 15350 27464
rect 15562 27452 15568 27464
rect 15523 27424 15568 27452
rect 15562 27412 15568 27424
rect 15620 27412 15626 27464
rect 15654 27412 15660 27464
rect 15712 27452 15718 27464
rect 15841 27455 15899 27461
rect 15712 27424 15757 27452
rect 15712 27412 15718 27424
rect 15841 27421 15853 27455
rect 15887 27421 15899 27455
rect 16574 27452 16580 27464
rect 16487 27424 16580 27452
rect 15841 27415 15899 27421
rect 15194 27384 15200 27396
rect 14660 27356 15200 27384
rect 15194 27344 15200 27356
rect 15252 27344 15258 27396
rect 15856 27384 15884 27415
rect 16574 27412 16580 27424
rect 16632 27452 16638 27464
rect 17405 27455 17463 27461
rect 17405 27452 17417 27455
rect 16632 27424 17417 27452
rect 16632 27412 16638 27424
rect 17405 27421 17417 27424
rect 17451 27452 17463 27455
rect 17494 27452 17500 27464
rect 17451 27424 17500 27452
rect 17451 27421 17463 27424
rect 17405 27415 17463 27421
rect 17494 27412 17500 27424
rect 17552 27412 17558 27464
rect 18064 27461 18092 27492
rect 22554 27480 22560 27492
rect 22612 27480 22618 27532
rect 46477 27523 46535 27529
rect 46477 27489 46489 27523
rect 46523 27520 46535 27523
rect 47210 27520 47216 27532
rect 46523 27492 47216 27520
rect 46523 27489 46535 27492
rect 46477 27483 46535 27489
rect 47210 27480 47216 27492
rect 47268 27480 47274 27532
rect 48222 27520 48228 27532
rect 48183 27492 48228 27520
rect 48222 27480 48228 27492
rect 48280 27480 48286 27532
rect 17589 27455 17647 27461
rect 17589 27421 17601 27455
rect 17635 27421 17647 27455
rect 17589 27415 17647 27421
rect 18049 27455 18107 27461
rect 18049 27421 18061 27455
rect 18095 27421 18107 27455
rect 18049 27415 18107 27421
rect 18233 27455 18291 27461
rect 18233 27421 18245 27455
rect 18279 27421 18291 27455
rect 20162 27452 20168 27464
rect 20123 27424 20168 27452
rect 18233 27415 18291 27421
rect 15672 27356 15884 27384
rect 16761 27387 16819 27393
rect 5902 27316 5908 27328
rect 5863 27288 5908 27316
rect 5902 27276 5908 27288
rect 5960 27276 5966 27328
rect 6362 27316 6368 27328
rect 6323 27288 6368 27316
rect 6362 27276 6368 27288
rect 6420 27276 6426 27328
rect 7558 27276 7564 27328
rect 7616 27316 7622 27328
rect 8573 27319 8631 27325
rect 8573 27316 8585 27319
rect 7616 27288 8585 27316
rect 7616 27276 7622 27288
rect 8573 27285 8585 27288
rect 8619 27285 8631 27319
rect 13446 27316 13452 27328
rect 13407 27288 13452 27316
rect 8573 27279 8631 27285
rect 13446 27276 13452 27288
rect 13504 27276 13510 27328
rect 13538 27276 13544 27328
rect 13596 27316 13602 27328
rect 15470 27316 15476 27328
rect 13596 27288 15476 27316
rect 13596 27276 13602 27288
rect 15470 27276 15476 27288
rect 15528 27316 15534 27328
rect 15672 27316 15700 27356
rect 16761 27353 16773 27387
rect 16807 27384 16819 27387
rect 17218 27384 17224 27396
rect 16807 27356 17224 27384
rect 16807 27353 16819 27356
rect 16761 27347 16819 27353
rect 17218 27344 17224 27356
rect 17276 27384 17282 27396
rect 17604 27384 17632 27415
rect 17276 27356 17632 27384
rect 17276 27344 17282 27356
rect 15528 27288 15700 27316
rect 15528 27276 15534 27288
rect 15746 27276 15752 27328
rect 15804 27316 15810 27328
rect 17589 27319 17647 27325
rect 17589 27316 17601 27319
rect 15804 27288 17601 27316
rect 15804 27276 15810 27288
rect 17589 27285 17601 27288
rect 17635 27316 17647 27319
rect 18248 27316 18276 27415
rect 20162 27412 20168 27424
rect 20220 27412 20226 27464
rect 20806 27412 20812 27464
rect 20864 27452 20870 27464
rect 20901 27455 20959 27461
rect 20901 27452 20913 27455
rect 20864 27424 20913 27452
rect 20864 27412 20870 27424
rect 20901 27421 20913 27424
rect 20947 27421 20959 27455
rect 20901 27415 20959 27421
rect 21082 27412 21088 27464
rect 21140 27452 21146 27464
rect 21450 27452 21456 27464
rect 21140 27424 21456 27452
rect 21140 27412 21146 27424
rect 21450 27412 21456 27424
rect 21508 27412 21514 27464
rect 24581 27455 24639 27461
rect 24581 27421 24593 27455
rect 24627 27452 24639 27455
rect 26418 27452 26424 27464
rect 24627 27424 26188 27452
rect 26379 27424 26424 27452
rect 24627 27421 24639 27424
rect 24581 27415 24639 27421
rect 24854 27393 24860 27396
rect 24848 27384 24860 27393
rect 24815 27356 24860 27384
rect 24848 27347 24860 27356
rect 24854 27344 24860 27347
rect 24912 27344 24918 27396
rect 26160 27384 26188 27424
rect 26418 27412 26424 27424
rect 26476 27412 26482 27464
rect 28534 27412 28540 27464
rect 28592 27452 28598 27464
rect 28905 27455 28963 27461
rect 28905 27452 28917 27455
rect 28592 27424 28917 27452
rect 28592 27412 28598 27424
rect 28905 27421 28917 27424
rect 28951 27421 28963 27455
rect 28905 27415 28963 27421
rect 29181 27455 29239 27461
rect 29181 27421 29193 27455
rect 29227 27452 29239 27455
rect 29270 27452 29276 27464
rect 29227 27424 29276 27452
rect 29227 27421 29239 27424
rect 29181 27415 29239 27421
rect 29270 27412 29276 27424
rect 29328 27412 29334 27464
rect 31202 27452 31208 27464
rect 31115 27424 31208 27452
rect 31202 27412 31208 27424
rect 31260 27452 31266 27464
rect 32766 27452 32772 27464
rect 31260 27424 32772 27452
rect 31260 27412 31266 27424
rect 32766 27412 32772 27424
rect 32824 27412 32830 27464
rect 33594 27452 33600 27464
rect 33555 27424 33600 27452
rect 33594 27412 33600 27424
rect 33652 27412 33658 27464
rect 34882 27452 34888 27464
rect 34843 27424 34888 27452
rect 34882 27412 34888 27424
rect 34940 27412 34946 27464
rect 35066 27452 35072 27464
rect 35027 27424 35072 27452
rect 35066 27412 35072 27424
rect 35124 27412 35130 27464
rect 35710 27452 35716 27464
rect 35671 27424 35716 27452
rect 35710 27412 35716 27424
rect 35768 27412 35774 27464
rect 35897 27455 35955 27461
rect 35897 27421 35909 27455
rect 35943 27452 35955 27455
rect 36170 27452 36176 27464
rect 35943 27424 36176 27452
rect 35943 27421 35955 27424
rect 35897 27415 35955 27421
rect 36170 27412 36176 27424
rect 36228 27412 36234 27464
rect 38102 27452 38108 27464
rect 38063 27424 38108 27452
rect 38102 27412 38108 27424
rect 38160 27412 38166 27464
rect 26234 27384 26240 27396
rect 26147 27356 26240 27384
rect 26234 27344 26240 27356
rect 26292 27384 26298 27396
rect 27154 27384 27160 27396
rect 26292 27356 27160 27384
rect 26292 27344 26298 27356
rect 27154 27344 27160 27356
rect 27212 27344 27218 27396
rect 31294 27344 31300 27396
rect 31352 27384 31358 27396
rect 31450 27387 31508 27393
rect 31450 27384 31462 27387
rect 31352 27356 31462 27384
rect 31352 27344 31358 27356
rect 31450 27353 31462 27356
rect 31496 27353 31508 27387
rect 31450 27347 31508 27353
rect 35253 27387 35311 27393
rect 35253 27353 35265 27387
rect 35299 27384 35311 27387
rect 36446 27384 36452 27396
rect 35299 27356 36452 27384
rect 35299 27353 35311 27356
rect 35253 27347 35311 27353
rect 36446 27344 36452 27356
rect 36504 27344 36510 27396
rect 38372 27387 38430 27393
rect 38372 27353 38384 27387
rect 38418 27384 38430 27387
rect 38562 27384 38568 27396
rect 38418 27356 38568 27384
rect 38418 27353 38430 27356
rect 38372 27347 38430 27353
rect 38562 27344 38568 27356
rect 38620 27344 38626 27396
rect 46661 27387 46719 27393
rect 46661 27353 46673 27387
rect 46707 27384 46719 27387
rect 47854 27384 47860 27396
rect 46707 27356 47860 27384
rect 46707 27353 46719 27356
rect 46661 27347 46719 27353
rect 47854 27344 47860 27356
rect 47912 27344 47918 27396
rect 17635 27288 18276 27316
rect 17635 27285 17647 27288
rect 17589 27279 17647 27285
rect 25038 27276 25044 27328
rect 25096 27316 25102 27328
rect 25961 27319 26019 27325
rect 25961 27316 25973 27319
rect 25096 27288 25973 27316
rect 25096 27276 25102 27288
rect 25961 27285 25973 27288
rect 26007 27285 26019 27319
rect 28718 27316 28724 27328
rect 28679 27288 28724 27316
rect 25961 27279 26019 27285
rect 28718 27276 28724 27288
rect 28776 27276 28782 27328
rect 32122 27276 32128 27328
rect 32180 27316 32186 27328
rect 32585 27319 32643 27325
rect 32585 27316 32597 27319
rect 32180 27288 32597 27316
rect 32180 27276 32186 27288
rect 32585 27285 32597 27288
rect 32631 27285 32643 27319
rect 32585 27279 32643 27285
rect 33413 27319 33471 27325
rect 33413 27285 33425 27319
rect 33459 27316 33471 27319
rect 33502 27316 33508 27328
rect 33459 27288 33508 27316
rect 33459 27285 33471 27288
rect 33413 27279 33471 27285
rect 33502 27276 33508 27288
rect 33560 27276 33566 27328
rect 35802 27316 35808 27328
rect 35763 27288 35808 27316
rect 35802 27276 35808 27288
rect 35860 27276 35866 27328
rect 39482 27316 39488 27328
rect 39443 27288 39488 27316
rect 39482 27276 39488 27288
rect 39540 27276 39546 27328
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 5718 27112 5724 27124
rect 5679 27084 5724 27112
rect 5718 27072 5724 27084
rect 5776 27072 5782 27124
rect 7377 27115 7435 27121
rect 7377 27081 7389 27115
rect 7423 27081 7435 27115
rect 9398 27112 9404 27124
rect 9359 27084 9404 27112
rect 7377 27075 7435 27081
rect 4608 27047 4666 27053
rect 4608 27013 4620 27047
rect 4654 27044 4666 27047
rect 6362 27044 6368 27056
rect 4654 27016 6368 27044
rect 4654 27013 4666 27016
rect 4608 27007 4666 27013
rect 6362 27004 6368 27016
rect 6420 27004 6426 27056
rect 7392 27044 7420 27075
rect 9398 27072 9404 27084
rect 9456 27072 9462 27124
rect 12526 27112 12532 27124
rect 12487 27084 12532 27112
rect 12526 27072 12532 27084
rect 12584 27072 12590 27124
rect 14553 27115 14611 27121
rect 14553 27081 14565 27115
rect 14599 27112 14611 27115
rect 14642 27112 14648 27124
rect 14599 27084 14648 27112
rect 14599 27081 14611 27084
rect 14553 27075 14611 27081
rect 14642 27072 14648 27084
rect 14700 27072 14706 27124
rect 15654 27072 15660 27124
rect 15712 27112 15718 27124
rect 16025 27115 16083 27121
rect 16025 27112 16037 27115
rect 15712 27084 16037 27112
rect 15712 27072 15718 27084
rect 16025 27081 16037 27084
rect 16071 27081 16083 27115
rect 16025 27075 16083 27081
rect 16850 27072 16856 27124
rect 16908 27112 16914 27124
rect 17313 27115 17371 27121
rect 17313 27112 17325 27115
rect 16908 27084 17325 27112
rect 16908 27072 16914 27084
rect 17313 27081 17325 27084
rect 17359 27112 17371 27115
rect 18598 27112 18604 27124
rect 17359 27084 18604 27112
rect 17359 27081 17371 27084
rect 17313 27075 17371 27081
rect 18598 27072 18604 27084
rect 18656 27072 18662 27124
rect 24397 27115 24455 27121
rect 24397 27081 24409 27115
rect 24443 27112 24455 27115
rect 24578 27112 24584 27124
rect 24443 27084 24584 27112
rect 24443 27081 24455 27084
rect 24397 27075 24455 27081
rect 24578 27072 24584 27084
rect 24636 27072 24642 27124
rect 28537 27115 28595 27121
rect 28537 27081 28549 27115
rect 28583 27112 28595 27115
rect 28626 27112 28632 27124
rect 28583 27084 28632 27112
rect 28583 27081 28595 27084
rect 28537 27075 28595 27081
rect 28626 27072 28632 27084
rect 28684 27072 28690 27124
rect 32122 27072 32128 27124
rect 32180 27112 32186 27124
rect 34882 27112 34888 27124
rect 32180 27084 34888 27112
rect 32180 27072 32186 27084
rect 34882 27072 34888 27084
rect 34940 27112 34946 27124
rect 34940 27084 35296 27112
rect 34940 27072 34946 27084
rect 8266 27047 8324 27053
rect 8266 27044 8278 27047
rect 7392 27016 8278 27044
rect 8266 27013 8278 27016
rect 8312 27013 8324 27047
rect 25222 27044 25228 27056
rect 8266 27007 8324 27013
rect 24872 27016 25228 27044
rect 4341 26979 4399 26985
rect 4341 26945 4353 26979
rect 4387 26976 4399 26979
rect 5166 26976 5172 26988
rect 4387 26948 5172 26976
rect 4387 26945 4399 26948
rect 4341 26939 4399 26945
rect 5166 26936 5172 26948
rect 5224 26936 5230 26988
rect 5902 26936 5908 26988
rect 5960 26976 5966 26988
rect 6733 26979 6791 26985
rect 6733 26976 6745 26979
rect 5960 26948 6745 26976
rect 5960 26936 5966 26948
rect 6733 26945 6745 26948
rect 6779 26945 6791 26979
rect 7558 26976 7564 26988
rect 7519 26948 7564 26976
rect 6733 26939 6791 26945
rect 7558 26936 7564 26948
rect 7616 26936 7622 26988
rect 12710 26976 12716 26988
rect 12671 26948 12716 26976
rect 12710 26936 12716 26948
rect 12768 26936 12774 26988
rect 13538 26976 13544 26988
rect 13499 26948 13544 26976
rect 13538 26936 13544 26948
rect 13596 26936 13602 26988
rect 13725 26979 13783 26985
rect 13725 26945 13737 26979
rect 13771 26976 13783 26979
rect 14369 26979 14427 26985
rect 14369 26976 14381 26979
rect 13771 26948 14381 26976
rect 13771 26945 13783 26948
rect 13725 26939 13783 26945
rect 14369 26945 14381 26948
rect 14415 26945 14427 26979
rect 14369 26939 14427 26945
rect 15933 26979 15991 26985
rect 15933 26945 15945 26979
rect 15979 26976 15991 26979
rect 16574 26976 16580 26988
rect 15979 26948 16580 26976
rect 15979 26945 15991 26948
rect 15933 26939 15991 26945
rect 16574 26936 16580 26948
rect 16632 26936 16638 26988
rect 17218 26976 17224 26988
rect 17179 26948 17224 26976
rect 17218 26936 17224 26948
rect 17276 26936 17282 26988
rect 20530 26976 20536 26988
rect 20491 26948 20536 26976
rect 20530 26936 20536 26948
rect 20588 26936 20594 26988
rect 20714 26976 20720 26988
rect 20675 26948 20720 26976
rect 20714 26936 20720 26948
rect 20772 26936 20778 26988
rect 22462 26976 22468 26988
rect 22423 26948 22468 26976
rect 22462 26936 22468 26948
rect 22520 26936 22526 26988
rect 24581 26979 24639 26985
rect 24581 26945 24593 26979
rect 24627 26945 24639 26979
rect 24581 26939 24639 26945
rect 7098 26868 7104 26920
rect 7156 26908 7162 26920
rect 8018 26908 8024 26920
rect 7156 26880 8024 26908
rect 7156 26868 7162 26880
rect 8018 26868 8024 26880
rect 8076 26868 8082 26920
rect 14182 26908 14188 26920
rect 14143 26880 14188 26908
rect 14182 26868 14188 26880
rect 14240 26908 14246 26920
rect 15562 26908 15568 26920
rect 14240 26880 15568 26908
rect 14240 26868 14246 26880
rect 15562 26868 15568 26880
rect 15620 26868 15626 26920
rect 20732 26840 20760 26936
rect 20809 26911 20867 26917
rect 20809 26877 20821 26911
rect 20855 26908 20867 26911
rect 22554 26908 22560 26920
rect 20855 26880 22560 26908
rect 20855 26877 20867 26880
rect 20809 26871 20867 26877
rect 22554 26868 22560 26880
rect 22612 26908 22618 26920
rect 22741 26911 22799 26917
rect 22741 26908 22753 26911
rect 22612 26880 22753 26908
rect 22612 26868 22618 26880
rect 22741 26877 22753 26880
rect 22787 26877 22799 26911
rect 24596 26908 24624 26939
rect 24670 26936 24676 26988
rect 24728 26976 24734 26988
rect 24872 26985 24900 27016
rect 25222 27004 25228 27016
rect 25280 27004 25286 27056
rect 26605 27047 26663 27053
rect 26605 27013 26617 27047
rect 26651 27044 26663 27047
rect 26694 27044 26700 27056
rect 26651 27016 26700 27044
rect 26651 27013 26663 27016
rect 26605 27007 26663 27013
rect 26694 27004 26700 27016
rect 26752 27004 26758 27056
rect 28718 27004 28724 27056
rect 28776 27044 28782 27056
rect 29242 27047 29300 27053
rect 29242 27044 29254 27047
rect 28776 27016 29254 27044
rect 28776 27004 28782 27016
rect 29242 27013 29254 27016
rect 29288 27013 29300 27047
rect 29242 27007 29300 27013
rect 29454 27004 29460 27056
rect 29512 27004 29518 27056
rect 35268 27053 35296 27084
rect 35710 27072 35716 27124
rect 35768 27112 35774 27124
rect 35989 27115 36047 27121
rect 35989 27112 36001 27115
rect 35768 27084 36001 27112
rect 35768 27072 35774 27084
rect 35989 27081 36001 27084
rect 36035 27081 36047 27115
rect 38562 27112 38568 27124
rect 38523 27084 38568 27112
rect 35989 27075 36047 27081
rect 38562 27072 38568 27084
rect 38620 27072 38626 27124
rect 35253 27047 35311 27053
rect 31588 27016 34376 27044
rect 24857 26979 24915 26985
rect 24857 26976 24869 26979
rect 24728 26948 24869 26976
rect 24728 26936 24734 26948
rect 24857 26945 24869 26948
rect 24903 26945 24915 26979
rect 25038 26976 25044 26988
rect 24999 26948 25044 26976
rect 24857 26939 24915 26945
rect 25038 26936 25044 26948
rect 25096 26936 25102 26988
rect 25866 26976 25872 26988
rect 25827 26948 25872 26976
rect 25866 26936 25872 26948
rect 25924 26936 25930 26988
rect 26329 26979 26387 26985
rect 26329 26945 26341 26979
rect 26375 26945 26387 26979
rect 27154 26976 27160 26988
rect 27115 26948 27160 26976
rect 26329 26939 26387 26945
rect 24946 26908 24952 26920
rect 24596 26880 24952 26908
rect 22741 26871 22799 26877
rect 24946 26868 24952 26880
rect 25004 26868 25010 26920
rect 25590 26868 25596 26920
rect 25648 26908 25654 26920
rect 26344 26908 26372 26939
rect 27154 26936 27160 26948
rect 27212 26936 27218 26988
rect 27246 26936 27252 26988
rect 27304 26976 27310 26988
rect 27413 26979 27471 26985
rect 27413 26976 27425 26979
rect 27304 26948 27425 26976
rect 27304 26936 27310 26948
rect 27413 26945 27425 26948
rect 27459 26945 27471 26979
rect 27413 26939 27471 26945
rect 28997 26979 29055 26985
rect 28997 26945 29009 26979
rect 29043 26976 29055 26979
rect 29472 26976 29500 27004
rect 31588 26988 31616 27016
rect 31202 26976 31208 26988
rect 29043 26948 31208 26976
rect 29043 26945 29055 26948
rect 28997 26939 29055 26945
rect 31202 26936 31208 26948
rect 31260 26936 31266 26988
rect 31297 26979 31355 26985
rect 31297 26945 31309 26979
rect 31343 26945 31355 26979
rect 31570 26976 31576 26988
rect 31531 26948 31576 26976
rect 31297 26939 31355 26945
rect 25648 26880 26372 26908
rect 31312 26908 31340 26939
rect 31570 26936 31576 26948
rect 31628 26936 31634 26988
rect 31754 26936 31760 26988
rect 31812 26976 31818 26988
rect 33502 26985 33508 26988
rect 33496 26976 33508 26985
rect 31812 26948 31857 26976
rect 33463 26948 33508 26976
rect 31812 26936 31818 26948
rect 33496 26939 33508 26948
rect 33502 26936 33508 26939
rect 33560 26936 33566 26988
rect 32398 26908 32404 26920
rect 31312 26880 32404 26908
rect 25648 26868 25654 26880
rect 32398 26868 32404 26880
rect 32456 26868 32462 26920
rect 32766 26868 32772 26920
rect 32824 26908 32830 26920
rect 33229 26911 33287 26917
rect 33229 26908 33241 26911
rect 32824 26880 33241 26908
rect 32824 26868 32830 26880
rect 33229 26877 33241 26880
rect 33275 26877 33287 26911
rect 33229 26871 33287 26877
rect 23658 26840 23664 26852
rect 20732 26812 23664 26840
rect 23658 26800 23664 26812
rect 23716 26800 23722 26852
rect 34348 26840 34376 27016
rect 35253 27013 35265 27047
rect 35299 27044 35311 27047
rect 38378 27044 38384 27056
rect 35299 27016 36124 27044
rect 35299 27013 35311 27016
rect 35253 27007 35311 27013
rect 34606 26936 34612 26988
rect 34664 26976 34670 26988
rect 35066 26976 35072 26988
rect 34664 26948 35072 26976
rect 34664 26936 34670 26948
rect 35066 26936 35072 26948
rect 35124 26936 35130 26988
rect 36096 26985 36124 27016
rect 37292 27016 38384 27044
rect 35897 26979 35955 26985
rect 35897 26945 35909 26979
rect 35943 26945 35955 26979
rect 35897 26939 35955 26945
rect 36081 26979 36139 26985
rect 36081 26945 36093 26979
rect 36127 26945 36139 26979
rect 36081 26939 36139 26945
rect 35084 26908 35112 26936
rect 35912 26908 35940 26939
rect 35084 26880 35940 26908
rect 37292 26840 37320 27016
rect 37642 26976 37648 26988
rect 37603 26948 37648 26976
rect 37642 26936 37648 26948
rect 37700 26936 37706 26988
rect 37936 26985 37964 27016
rect 38378 27004 38384 27016
rect 38436 27004 38442 27056
rect 37921 26979 37979 26985
rect 37921 26945 37933 26979
rect 37967 26945 37979 26979
rect 37921 26939 37979 26945
rect 38010 26936 38016 26988
rect 38068 26976 38074 26988
rect 38105 26979 38163 26985
rect 38105 26976 38117 26979
rect 38068 26948 38117 26976
rect 38068 26936 38074 26948
rect 38105 26945 38117 26948
rect 38151 26945 38163 26979
rect 38105 26939 38163 26945
rect 38749 26979 38807 26985
rect 38749 26945 38761 26979
rect 38795 26945 38807 26979
rect 38749 26939 38807 26945
rect 37461 26911 37519 26917
rect 37461 26877 37473 26911
rect 37507 26908 37519 26911
rect 38764 26908 38792 26939
rect 38930 26936 38936 26988
rect 38988 26976 38994 26988
rect 39025 26979 39083 26985
rect 39025 26976 39037 26979
rect 38988 26948 39037 26976
rect 38988 26936 38994 26948
rect 39025 26945 39037 26948
rect 39071 26976 39083 26979
rect 39482 26976 39488 26988
rect 39071 26948 39488 26976
rect 39071 26945 39083 26948
rect 39025 26939 39083 26945
rect 39482 26936 39488 26948
rect 39540 26936 39546 26988
rect 37507 26880 38792 26908
rect 37507 26877 37519 26880
rect 37461 26871 37519 26877
rect 34348 26812 37320 26840
rect 6546 26772 6552 26784
rect 6507 26744 6552 26772
rect 6546 26732 6552 26744
rect 6604 26732 6610 26784
rect 20346 26772 20352 26784
rect 20307 26744 20352 26772
rect 20346 26732 20352 26744
rect 20404 26732 20410 26784
rect 22278 26772 22284 26784
rect 22239 26744 22284 26772
rect 22278 26732 22284 26744
rect 22336 26732 22342 26784
rect 22649 26775 22707 26781
rect 22649 26741 22661 26775
rect 22695 26772 22707 26775
rect 24578 26772 24584 26784
rect 22695 26744 24584 26772
rect 22695 26741 22707 26744
rect 22649 26735 22707 26741
rect 24578 26732 24584 26744
rect 24636 26772 24642 26784
rect 24762 26772 24768 26784
rect 24636 26744 24768 26772
rect 24636 26732 24642 26744
rect 24762 26732 24768 26744
rect 24820 26732 24826 26784
rect 25130 26732 25136 26784
rect 25188 26772 25194 26784
rect 25774 26772 25780 26784
rect 25188 26744 25780 26772
rect 25188 26732 25194 26744
rect 25774 26732 25780 26744
rect 25832 26772 25838 26784
rect 28902 26772 28908 26784
rect 25832 26744 28908 26772
rect 25832 26732 25838 26744
rect 28902 26732 28908 26744
rect 28960 26732 28966 26784
rect 29178 26732 29184 26784
rect 29236 26772 29242 26784
rect 30377 26775 30435 26781
rect 30377 26772 30389 26775
rect 29236 26744 30389 26772
rect 29236 26732 29242 26744
rect 30377 26741 30389 26744
rect 30423 26741 30435 26775
rect 30377 26735 30435 26741
rect 31113 26775 31171 26781
rect 31113 26741 31125 26775
rect 31159 26772 31171 26775
rect 31478 26772 31484 26784
rect 31159 26744 31484 26772
rect 31159 26741 31171 26744
rect 31113 26735 31171 26741
rect 31478 26732 31484 26744
rect 31536 26732 31542 26784
rect 34606 26772 34612 26784
rect 34567 26744 34612 26772
rect 34606 26732 34612 26744
rect 34664 26732 34670 26784
rect 35437 26775 35495 26781
rect 35437 26741 35449 26775
rect 35483 26772 35495 26775
rect 36170 26772 36176 26784
rect 35483 26744 36176 26772
rect 35483 26741 35495 26744
rect 35437 26735 35495 26741
rect 36170 26732 36176 26744
rect 36228 26732 36234 26784
rect 38838 26732 38844 26784
rect 38896 26772 38902 26784
rect 38933 26775 38991 26781
rect 38933 26772 38945 26775
rect 38896 26744 38945 26772
rect 38896 26732 38902 26744
rect 38933 26741 38945 26744
rect 38979 26741 38991 26775
rect 38933 26735 38991 26741
rect 46474 26732 46480 26784
rect 46532 26772 46538 26784
rect 47949 26775 48007 26781
rect 47949 26772 47961 26775
rect 46532 26744 47961 26772
rect 46532 26732 46538 26744
rect 47949 26741 47961 26744
rect 47995 26741 48007 26775
rect 47949 26735 48007 26741
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 8386 26528 8392 26580
rect 8444 26568 8450 26580
rect 8481 26571 8539 26577
rect 8481 26568 8493 26571
rect 8444 26540 8493 26568
rect 8444 26528 8450 26540
rect 8481 26537 8493 26540
rect 8527 26537 8539 26571
rect 8481 26531 8539 26537
rect 13541 26571 13599 26577
rect 13541 26537 13553 26571
rect 13587 26568 13599 26571
rect 14182 26568 14188 26580
rect 13587 26540 14188 26568
rect 13587 26537 13599 26540
rect 13541 26531 13599 26537
rect 14182 26528 14188 26540
rect 14240 26528 14246 26580
rect 17218 26528 17224 26580
rect 17276 26568 17282 26580
rect 17957 26571 18015 26577
rect 17957 26568 17969 26571
rect 17276 26540 17969 26568
rect 17276 26528 17282 26540
rect 17957 26537 17969 26540
rect 18003 26537 18015 26571
rect 20714 26568 20720 26580
rect 17957 26531 18015 26537
rect 18708 26540 20720 26568
rect 6641 26503 6699 26509
rect 6641 26469 6653 26503
rect 6687 26500 6699 26503
rect 6914 26500 6920 26512
rect 6687 26472 6920 26500
rect 6687 26469 6699 26472
rect 6641 26463 6699 26469
rect 6914 26460 6920 26472
rect 6972 26460 6978 26512
rect 18046 26460 18052 26512
rect 18104 26500 18110 26512
rect 18417 26503 18475 26509
rect 18417 26500 18429 26503
rect 18104 26472 18429 26500
rect 18104 26460 18110 26472
rect 18417 26469 18429 26472
rect 18463 26469 18475 26503
rect 18417 26463 18475 26469
rect 5258 26364 5264 26376
rect 5219 26336 5264 26364
rect 5258 26324 5264 26336
rect 5316 26324 5322 26376
rect 5528 26367 5586 26373
rect 5528 26333 5540 26367
rect 5574 26364 5586 26367
rect 6546 26364 6552 26376
rect 5574 26336 6552 26364
rect 5574 26333 5586 26336
rect 5528 26327 5586 26333
rect 6546 26324 6552 26336
rect 6604 26324 6610 26376
rect 7098 26364 7104 26376
rect 7011 26336 7104 26364
rect 7098 26324 7104 26336
rect 7156 26324 7162 26376
rect 13446 26364 13452 26376
rect 13407 26336 13452 26364
rect 13446 26324 13452 26336
rect 13504 26324 13510 26376
rect 13630 26364 13636 26376
rect 13591 26336 13636 26364
rect 13630 26324 13636 26336
rect 13688 26324 13694 26376
rect 16577 26367 16635 26373
rect 16577 26333 16589 26367
rect 16623 26364 16635 26367
rect 17402 26364 17408 26376
rect 16623 26336 17408 26364
rect 16623 26333 16635 26336
rect 16577 26327 16635 26333
rect 5276 26296 5304 26324
rect 7116 26296 7144 26324
rect 5276 26268 7144 26296
rect 7368 26299 7426 26305
rect 7368 26265 7380 26299
rect 7414 26296 7426 26299
rect 7742 26296 7748 26308
rect 7414 26268 7748 26296
rect 7414 26265 7426 26268
rect 7368 26259 7426 26265
rect 7742 26256 7748 26268
rect 7800 26256 7806 26308
rect 16592 26296 16620 26327
rect 17402 26324 17408 26336
rect 17460 26324 17466 26376
rect 18598 26364 18604 26376
rect 18559 26336 18604 26364
rect 18598 26324 18604 26336
rect 18656 26324 18662 26376
rect 18708 26373 18736 26540
rect 20714 26528 20720 26540
rect 20772 26528 20778 26580
rect 21082 26568 21088 26580
rect 21043 26540 21088 26568
rect 21082 26528 21088 26540
rect 21140 26528 21146 26580
rect 22646 26528 22652 26580
rect 22704 26568 22710 26580
rect 23106 26568 23112 26580
rect 22704 26540 23112 26568
rect 22704 26528 22710 26540
rect 23106 26528 23112 26540
rect 23164 26568 23170 26580
rect 23385 26571 23443 26577
rect 23385 26568 23397 26571
rect 23164 26540 23397 26568
rect 23164 26528 23170 26540
rect 23385 26537 23397 26540
rect 23431 26537 23443 26571
rect 23385 26531 23443 26537
rect 24949 26571 25007 26577
rect 24949 26537 24961 26571
rect 24995 26568 25007 26571
rect 25130 26568 25136 26580
rect 24995 26540 25136 26568
rect 24995 26537 25007 26540
rect 24949 26531 25007 26537
rect 25130 26528 25136 26540
rect 25188 26528 25194 26580
rect 25498 26528 25504 26580
rect 25556 26568 25562 26580
rect 30374 26568 30380 26580
rect 25556 26540 30380 26568
rect 25556 26528 25562 26540
rect 30374 26528 30380 26540
rect 30432 26568 30438 26580
rect 31021 26571 31079 26577
rect 31021 26568 31033 26571
rect 30432 26540 31033 26568
rect 30432 26528 30438 26540
rect 31021 26537 31033 26540
rect 31067 26568 31079 26571
rect 31067 26540 31754 26568
rect 31067 26537 31079 26540
rect 31021 26531 31079 26537
rect 25682 26500 25688 26512
rect 25643 26472 25688 26500
rect 25682 26460 25688 26472
rect 25740 26460 25746 26512
rect 26326 26460 26332 26512
rect 26384 26500 26390 26512
rect 26513 26503 26571 26509
rect 26513 26500 26525 26503
rect 26384 26472 26525 26500
rect 26384 26460 26390 26472
rect 26513 26469 26525 26472
rect 26559 26469 26571 26503
rect 28534 26500 28540 26512
rect 28495 26472 28540 26500
rect 26513 26463 26571 26469
rect 19426 26392 19432 26444
rect 19484 26432 19490 26444
rect 19705 26435 19763 26441
rect 19705 26432 19717 26435
rect 19484 26404 19717 26432
rect 19484 26392 19490 26404
rect 19705 26401 19717 26404
rect 19751 26401 19763 26435
rect 26234 26432 26240 26444
rect 19705 26395 19763 26401
rect 23768 26404 26240 26432
rect 18693 26367 18751 26373
rect 18693 26333 18705 26367
rect 18739 26333 18751 26367
rect 18693 26327 18751 26333
rect 19972 26367 20030 26373
rect 19972 26333 19984 26367
rect 20018 26364 20030 26367
rect 20346 26364 20352 26376
rect 20018 26336 20352 26364
rect 20018 26333 20030 26336
rect 19972 26327 20030 26333
rect 20346 26324 20352 26336
rect 20404 26324 20410 26376
rect 22005 26367 22063 26373
rect 22005 26333 22017 26367
rect 22051 26364 22063 26367
rect 23768 26364 23796 26404
rect 26234 26392 26240 26404
rect 26292 26392 26298 26444
rect 26528 26432 26556 26463
rect 28534 26460 28540 26472
rect 28592 26460 28598 26512
rect 31726 26500 31754 26540
rect 31938 26500 31944 26512
rect 31726 26472 31944 26500
rect 31938 26460 31944 26472
rect 31996 26460 32002 26512
rect 35894 26500 35900 26512
rect 33888 26472 35900 26500
rect 32766 26432 32772 26444
rect 26528 26404 27660 26432
rect 32727 26404 32772 26432
rect 24670 26364 24676 26376
rect 22051 26336 23796 26364
rect 24631 26336 24676 26364
rect 22051 26333 22063 26336
rect 22005 26327 22063 26333
rect 16500 26268 16620 26296
rect 16844 26299 16902 26305
rect 14826 26188 14832 26240
rect 14884 26228 14890 26240
rect 16500 26228 16528 26268
rect 16844 26265 16856 26299
rect 16890 26296 16902 26299
rect 17862 26296 17868 26308
rect 16890 26268 17868 26296
rect 16890 26265 16902 26268
rect 16844 26259 16902 26265
rect 17862 26256 17868 26268
rect 17920 26256 17926 26308
rect 18417 26299 18475 26305
rect 18417 26265 18429 26299
rect 18463 26296 18475 26299
rect 18506 26296 18512 26308
rect 18463 26268 18512 26296
rect 18463 26265 18475 26268
rect 18417 26259 18475 26265
rect 18506 26256 18512 26268
rect 18564 26256 18570 26308
rect 20622 26256 20628 26308
rect 20680 26296 20686 26308
rect 22020 26296 22048 26327
rect 24670 26324 24676 26336
rect 24728 26324 24734 26376
rect 25501 26367 25559 26373
rect 25501 26333 25513 26367
rect 25547 26364 25559 26367
rect 25590 26364 25596 26376
rect 25547 26336 25596 26364
rect 25547 26333 25559 26336
rect 25501 26327 25559 26333
rect 25590 26324 25596 26336
rect 25648 26324 25654 26376
rect 25682 26324 25688 26376
rect 25740 26364 25746 26376
rect 27632 26373 27660 26404
rect 32766 26392 32772 26404
rect 32824 26392 32830 26444
rect 27341 26367 27399 26373
rect 27341 26364 27353 26367
rect 25740 26336 27353 26364
rect 25740 26324 25746 26336
rect 27341 26333 27353 26336
rect 27387 26333 27399 26367
rect 27341 26327 27399 26333
rect 27617 26367 27675 26373
rect 27617 26333 27629 26367
rect 27663 26333 27675 26367
rect 27617 26327 27675 26333
rect 27801 26367 27859 26373
rect 27801 26333 27813 26367
rect 27847 26364 27859 26367
rect 28626 26364 28632 26376
rect 27847 26336 28632 26364
rect 27847 26333 27859 26336
rect 27801 26327 27859 26333
rect 22278 26305 22284 26308
rect 22272 26296 22284 26305
rect 20680 26268 22048 26296
rect 22239 26268 22284 26296
rect 20680 26256 20686 26268
rect 22272 26259 22284 26268
rect 22278 26256 22284 26259
rect 22336 26256 22342 26308
rect 25130 26296 25136 26308
rect 24964 26268 25136 26296
rect 14884 26200 16528 26228
rect 14884 26188 14890 26200
rect 19978 26188 19984 26240
rect 20036 26228 20042 26240
rect 24964 26228 24992 26268
rect 25130 26256 25136 26268
rect 25188 26256 25194 26308
rect 26329 26299 26387 26305
rect 26329 26296 26341 26299
rect 26160 26268 26341 26296
rect 20036 26200 24992 26228
rect 20036 26188 20042 26200
rect 25038 26188 25044 26240
rect 25096 26228 25102 26240
rect 26160 26228 26188 26268
rect 26329 26265 26341 26268
rect 26375 26296 26387 26299
rect 27062 26296 27068 26308
rect 26375 26268 27068 26296
rect 26375 26265 26387 26268
rect 26329 26259 26387 26265
rect 27062 26256 27068 26268
rect 27120 26256 27126 26308
rect 27632 26296 27660 26327
rect 28626 26324 28632 26336
rect 28684 26324 28690 26376
rect 28718 26324 28724 26376
rect 28776 26364 28782 26376
rect 28776 26336 28821 26364
rect 28776 26324 28782 26336
rect 28902 26324 28908 26376
rect 28960 26364 28966 26376
rect 28997 26367 29055 26373
rect 28997 26364 29009 26367
rect 28960 26336 29009 26364
rect 28960 26324 28966 26336
rect 28997 26333 29009 26336
rect 29043 26333 29055 26367
rect 29178 26364 29184 26376
rect 29139 26336 29184 26364
rect 28997 26327 29055 26333
rect 29178 26324 29184 26336
rect 29236 26324 29242 26376
rect 30742 26364 30748 26376
rect 29564 26336 30748 26364
rect 29564 26296 29592 26336
rect 30742 26324 30748 26336
rect 30800 26324 30806 26376
rect 31938 26364 31944 26376
rect 31851 26336 31944 26364
rect 31938 26324 31944 26336
rect 31996 26364 32002 26376
rect 33321 26367 33379 26373
rect 33321 26364 33333 26367
rect 31996 26336 33333 26364
rect 31996 26324 32002 26336
rect 33321 26333 33333 26336
rect 33367 26364 33379 26367
rect 33888 26364 33916 26472
rect 35894 26460 35900 26472
rect 35952 26460 35958 26512
rect 38838 26460 38844 26512
rect 38896 26500 38902 26512
rect 39393 26503 39451 26509
rect 39393 26500 39405 26503
rect 38896 26472 39405 26500
rect 38896 26460 38902 26472
rect 39393 26469 39405 26472
rect 39439 26469 39451 26503
rect 39393 26463 39451 26469
rect 35161 26435 35219 26441
rect 35161 26401 35173 26435
rect 35207 26432 35219 26435
rect 35710 26432 35716 26444
rect 35207 26404 35716 26432
rect 35207 26401 35219 26404
rect 35161 26395 35219 26401
rect 35710 26392 35716 26404
rect 35768 26392 35774 26444
rect 37921 26435 37979 26441
rect 37921 26401 37933 26435
rect 37967 26432 37979 26435
rect 46474 26432 46480 26444
rect 37967 26404 39252 26432
rect 46435 26404 46480 26432
rect 37967 26401 37979 26404
rect 37921 26395 37979 26401
rect 33367 26336 33916 26364
rect 35069 26367 35127 26373
rect 33367 26333 33379 26336
rect 33321 26327 33379 26333
rect 35069 26333 35081 26367
rect 35115 26364 35127 26367
rect 35802 26364 35808 26376
rect 35115 26336 35808 26364
rect 35115 26333 35127 26336
rect 35069 26327 35127 26333
rect 35802 26324 35808 26336
rect 35860 26324 35866 26376
rect 36078 26324 36084 26376
rect 36136 26364 36142 26376
rect 36357 26367 36415 26373
rect 36357 26364 36369 26367
rect 36136 26336 36369 26364
rect 36136 26324 36142 26336
rect 36357 26333 36369 26336
rect 36403 26333 36415 26367
rect 36538 26364 36544 26376
rect 36499 26336 36544 26364
rect 36357 26327 36415 26333
rect 36538 26324 36544 26336
rect 36596 26324 36602 26376
rect 37642 26324 37648 26376
rect 37700 26364 37706 26376
rect 38105 26367 38163 26373
rect 38105 26364 38117 26367
rect 37700 26336 38117 26364
rect 37700 26324 37706 26336
rect 38105 26333 38117 26336
rect 38151 26364 38163 26367
rect 38286 26364 38292 26376
rect 38151 26336 38292 26364
rect 38151 26333 38163 26336
rect 38105 26327 38163 26333
rect 38286 26324 38292 26336
rect 38344 26324 38350 26376
rect 38378 26324 38384 26376
rect 38436 26364 38442 26376
rect 38436 26336 38481 26364
rect 38436 26324 38442 26336
rect 38562 26324 38568 26376
rect 38620 26364 38626 26376
rect 39224 26373 39252 26404
rect 46474 26392 46480 26404
rect 46532 26392 46538 26444
rect 48222 26432 48228 26444
rect 48183 26404 48228 26432
rect 48222 26392 48228 26404
rect 48280 26392 48286 26444
rect 39209 26367 39267 26373
rect 38620 26336 38665 26364
rect 38620 26324 38626 26336
rect 39209 26333 39221 26367
rect 39255 26333 39267 26367
rect 39209 26327 39267 26333
rect 39485 26367 39543 26373
rect 39485 26333 39497 26367
rect 39531 26364 39543 26367
rect 40678 26364 40684 26376
rect 39531 26336 40684 26364
rect 39531 26333 39543 26336
rect 39485 26327 39543 26333
rect 40678 26324 40684 26336
rect 40736 26324 40742 26376
rect 29730 26296 29736 26308
rect 27632 26268 29592 26296
rect 29691 26268 29736 26296
rect 29730 26256 29736 26268
rect 29788 26256 29794 26308
rect 33778 26256 33784 26308
rect 33836 26296 33842 26308
rect 34057 26299 34115 26305
rect 34057 26296 34069 26299
rect 33836 26268 34069 26296
rect 33836 26256 33842 26268
rect 34057 26265 34069 26268
rect 34103 26265 34115 26299
rect 34057 26259 34115 26265
rect 35986 26256 35992 26308
rect 36044 26296 36050 26308
rect 36725 26299 36783 26305
rect 36725 26296 36737 26299
rect 36044 26268 36737 26296
rect 36044 26256 36050 26268
rect 36725 26265 36737 26268
rect 36771 26265 36783 26299
rect 36725 26259 36783 26265
rect 46661 26299 46719 26305
rect 46661 26265 46673 26299
rect 46707 26296 46719 26299
rect 47854 26296 47860 26308
rect 46707 26268 47860 26296
rect 46707 26265 46719 26268
rect 46661 26259 46719 26265
rect 47854 26256 47860 26268
rect 47912 26256 47918 26308
rect 25096 26200 26188 26228
rect 27157 26231 27215 26237
rect 25096 26188 25102 26200
rect 27157 26197 27169 26231
rect 27203 26228 27215 26231
rect 27338 26228 27344 26240
rect 27203 26200 27344 26228
rect 27203 26197 27215 26200
rect 27157 26191 27215 26197
rect 27338 26188 27344 26200
rect 27396 26188 27402 26240
rect 35434 26228 35440 26240
rect 35395 26200 35440 26228
rect 35434 26188 35440 26200
rect 35492 26188 35498 26240
rect 39022 26228 39028 26240
rect 38983 26200 39028 26228
rect 39022 26188 39028 26200
rect 39080 26188 39086 26240
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 7742 26024 7748 26036
rect 7703 25996 7748 26024
rect 7742 25984 7748 25996
rect 7800 25984 7806 26036
rect 17862 26024 17868 26036
rect 17823 25996 17868 26024
rect 17862 25984 17868 25996
rect 17920 25984 17926 26036
rect 20530 26024 20536 26036
rect 20491 25996 20536 26024
rect 20530 25984 20536 25996
rect 20588 25984 20594 26036
rect 22462 26024 22468 26036
rect 22423 25996 22468 26024
rect 22462 25984 22468 25996
rect 22520 25984 22526 26036
rect 25682 26024 25688 26036
rect 22848 25996 25688 26024
rect 12894 25916 12900 25968
rect 12952 25956 12958 25968
rect 22848 25956 22876 25996
rect 25682 25984 25688 25996
rect 25740 25984 25746 26036
rect 26053 26027 26111 26033
rect 26053 25993 26065 26027
rect 26099 26024 26111 26027
rect 26418 26024 26424 26036
rect 26099 25996 26424 26024
rect 26099 25993 26111 25996
rect 26053 25987 26111 25993
rect 26418 25984 26424 25996
rect 26476 25984 26482 26036
rect 27157 26027 27215 26033
rect 27157 25993 27169 26027
rect 27203 26024 27215 26027
rect 27246 26024 27252 26036
rect 27203 25996 27252 26024
rect 27203 25993 27215 25996
rect 27157 25987 27215 25993
rect 27246 25984 27252 25996
rect 27304 25984 27310 26036
rect 31294 26024 31300 26036
rect 31255 25996 31300 26024
rect 31294 25984 31300 25996
rect 31352 25984 31358 26036
rect 33505 26027 33563 26033
rect 33505 25993 33517 26027
rect 33551 26024 33563 26027
rect 33594 26024 33600 26036
rect 33551 25996 33600 26024
rect 33551 25993 33563 25996
rect 33505 25987 33563 25993
rect 33594 25984 33600 25996
rect 33652 25984 33658 26036
rect 33965 26027 34023 26033
rect 33965 25993 33977 26027
rect 34011 26024 34023 26027
rect 34701 26027 34759 26033
rect 34701 26024 34713 26027
rect 34011 25996 34713 26024
rect 34011 25993 34023 25996
rect 33965 25987 34023 25993
rect 34701 25993 34713 25996
rect 34747 25993 34759 26027
rect 34701 25987 34759 25993
rect 35161 26027 35219 26033
rect 35161 25993 35173 26027
rect 35207 26024 35219 26027
rect 35434 26024 35440 26036
rect 35207 25996 35440 26024
rect 35207 25993 35219 25996
rect 35161 25987 35219 25993
rect 35434 25984 35440 25996
rect 35492 25984 35498 26036
rect 40678 26024 40684 26036
rect 40639 25996 40684 26024
rect 40678 25984 40684 25996
rect 40736 25984 40742 26036
rect 47854 26024 47860 26036
rect 47815 25996 47860 26024
rect 47854 25984 47860 25996
rect 47912 25984 47918 26036
rect 23750 25956 23756 25968
rect 12952 25928 15976 25956
rect 12952 25916 12958 25928
rect 2222 25888 2228 25900
rect 2183 25860 2228 25888
rect 2222 25848 2228 25860
rect 2280 25848 2286 25900
rect 6825 25891 6883 25897
rect 6825 25857 6837 25891
rect 6871 25888 6883 25891
rect 7006 25888 7012 25900
rect 6871 25860 7012 25888
rect 6871 25857 6883 25860
rect 6825 25851 6883 25857
rect 7006 25848 7012 25860
rect 7064 25848 7070 25900
rect 7929 25891 7987 25897
rect 7929 25888 7941 25891
rect 7300 25860 7941 25888
rect 7300 25829 7328 25860
rect 7929 25857 7941 25860
rect 7975 25857 7987 25891
rect 7929 25851 7987 25857
rect 12713 25891 12771 25897
rect 12713 25857 12725 25891
rect 12759 25888 12771 25891
rect 12802 25888 12808 25900
rect 12759 25860 12808 25888
rect 12759 25857 12771 25860
rect 12713 25851 12771 25857
rect 12802 25848 12808 25860
rect 12860 25848 12866 25900
rect 13004 25897 13032 25928
rect 12989 25891 13047 25897
rect 12989 25857 13001 25891
rect 13035 25857 13047 25891
rect 12989 25851 13047 25857
rect 13173 25891 13231 25897
rect 13173 25857 13185 25891
rect 13219 25888 13231 25891
rect 13630 25888 13636 25900
rect 13219 25860 13636 25888
rect 13219 25857 13231 25860
rect 13173 25851 13231 25857
rect 13630 25848 13636 25860
rect 13688 25848 13694 25900
rect 15948 25897 15976 25928
rect 20732 25928 22876 25956
rect 22940 25928 23756 25956
rect 15657 25891 15715 25897
rect 15657 25857 15669 25891
rect 15703 25857 15715 25891
rect 15657 25851 15715 25857
rect 15933 25891 15991 25897
rect 15933 25857 15945 25891
rect 15979 25857 15991 25891
rect 15933 25851 15991 25857
rect 16117 25891 16175 25897
rect 16117 25857 16129 25891
rect 16163 25888 16175 25891
rect 16574 25888 16580 25900
rect 16163 25860 16580 25888
rect 16163 25857 16175 25860
rect 16117 25851 16175 25857
rect 7285 25823 7343 25829
rect 7285 25789 7297 25823
rect 7331 25789 7343 25823
rect 12820 25820 12848 25848
rect 15672 25820 15700 25851
rect 16574 25848 16580 25860
rect 16632 25888 16638 25900
rect 17034 25888 17040 25900
rect 16632 25860 17040 25888
rect 16632 25848 16638 25860
rect 17034 25848 17040 25860
rect 17092 25848 17098 25900
rect 18046 25888 18052 25900
rect 18007 25860 18052 25888
rect 18046 25848 18052 25860
rect 18104 25848 18110 25900
rect 20732 25897 20760 25928
rect 20717 25891 20775 25897
rect 20717 25888 20729 25891
rect 18156 25860 20729 25888
rect 18156 25820 18184 25860
rect 20717 25857 20729 25860
rect 20763 25857 20775 25891
rect 20717 25851 20775 25857
rect 20993 25891 21051 25897
rect 20993 25857 21005 25891
rect 21039 25857 21051 25891
rect 20993 25851 21051 25857
rect 12820 25792 18184 25820
rect 18325 25823 18383 25829
rect 7285 25783 7343 25789
rect 18325 25789 18337 25823
rect 18371 25789 18383 25823
rect 18325 25783 18383 25789
rect 1762 25644 1768 25696
rect 1820 25684 1826 25696
rect 2317 25687 2375 25693
rect 2317 25684 2329 25687
rect 1820 25656 2329 25684
rect 1820 25644 1826 25656
rect 2317 25653 2329 25656
rect 2363 25653 2375 25687
rect 6914 25684 6920 25696
rect 6875 25656 6920 25684
rect 2317 25647 2375 25653
rect 6914 25644 6920 25656
rect 6972 25644 6978 25696
rect 12526 25684 12532 25696
rect 12487 25656 12532 25684
rect 12526 25644 12532 25656
rect 12584 25644 12590 25696
rect 15473 25687 15531 25693
rect 15473 25653 15485 25687
rect 15519 25684 15531 25687
rect 16850 25684 16856 25696
rect 15519 25656 16856 25684
rect 15519 25653 15531 25656
rect 15473 25647 15531 25653
rect 16850 25644 16856 25656
rect 16908 25644 16914 25696
rect 17034 25644 17040 25696
rect 17092 25684 17098 25696
rect 18230 25684 18236 25696
rect 17092 25656 18236 25684
rect 17092 25644 17098 25656
rect 18230 25644 18236 25656
rect 18288 25644 18294 25696
rect 18340 25684 18368 25783
rect 21008 25752 21036 25851
rect 21082 25848 21088 25900
rect 21140 25888 21146 25900
rect 21177 25891 21235 25897
rect 21177 25888 21189 25891
rect 21140 25860 21189 25888
rect 21140 25848 21146 25860
rect 21177 25857 21189 25860
rect 21223 25857 21235 25891
rect 21177 25851 21235 25857
rect 21910 25848 21916 25900
rect 21968 25888 21974 25900
rect 22940 25897 22968 25928
rect 23750 25916 23756 25928
rect 23808 25956 23814 25968
rect 24670 25956 24676 25968
rect 23808 25928 24676 25956
rect 23808 25916 23814 25928
rect 24670 25916 24676 25928
rect 24728 25916 24734 25968
rect 25866 25956 25872 25968
rect 25827 25928 25872 25956
rect 25866 25916 25872 25928
rect 25924 25916 25930 25968
rect 32490 25916 32496 25968
rect 32548 25956 32554 25968
rect 35069 25959 35127 25965
rect 35069 25956 35081 25959
rect 32548 25928 35081 25956
rect 32548 25916 32554 25928
rect 35069 25925 35081 25928
rect 35115 25925 35127 25959
rect 35069 25919 35127 25925
rect 35989 25959 36047 25965
rect 35989 25925 36001 25959
rect 36035 25956 36047 25959
rect 36078 25956 36084 25968
rect 36035 25928 36084 25956
rect 36035 25925 36047 25928
rect 35989 25919 36047 25925
rect 36078 25916 36084 25928
rect 36136 25916 36142 25968
rect 36170 25916 36176 25968
rect 36228 25965 36234 25968
rect 36228 25959 36247 25965
rect 36235 25925 36247 25959
rect 36228 25919 36247 25925
rect 36228 25916 36234 25919
rect 39022 25916 39028 25968
rect 39080 25956 39086 25968
rect 39546 25959 39604 25965
rect 39546 25956 39558 25959
rect 39080 25928 39558 25956
rect 39080 25916 39086 25928
rect 39546 25925 39558 25928
rect 39592 25925 39604 25959
rect 39546 25919 39604 25925
rect 22649 25891 22707 25897
rect 22649 25888 22661 25891
rect 21968 25860 22661 25888
rect 21968 25848 21974 25860
rect 22649 25857 22661 25860
rect 22695 25857 22707 25891
rect 22649 25851 22707 25857
rect 22925 25891 22983 25897
rect 22925 25857 22937 25891
rect 22971 25857 22983 25891
rect 23106 25888 23112 25900
rect 23067 25860 23112 25888
rect 22925 25851 22983 25857
rect 23106 25848 23112 25860
rect 23164 25848 23170 25900
rect 25682 25888 25688 25900
rect 25643 25860 25688 25888
rect 25682 25848 25688 25860
rect 25740 25848 25746 25900
rect 27338 25888 27344 25900
rect 27299 25860 27344 25888
rect 27338 25848 27344 25860
rect 27396 25848 27402 25900
rect 27890 25888 27896 25900
rect 27448 25860 27896 25888
rect 23658 25780 23664 25832
rect 23716 25820 23722 25832
rect 27448 25820 27476 25860
rect 27890 25848 27896 25860
rect 27948 25888 27954 25900
rect 28169 25891 28227 25897
rect 28169 25888 28181 25891
rect 27948 25860 28181 25888
rect 27948 25848 27954 25860
rect 28169 25857 28181 25860
rect 28215 25857 28227 25891
rect 28169 25851 28227 25857
rect 28350 25848 28356 25900
rect 28408 25888 28414 25900
rect 30101 25891 30159 25897
rect 30101 25888 30113 25891
rect 28408 25860 30113 25888
rect 28408 25848 28414 25860
rect 30101 25857 30113 25860
rect 30147 25888 30159 25891
rect 31478 25888 31484 25900
rect 30147 25860 30871 25888
rect 31439 25860 31484 25888
rect 30147 25857 30159 25860
rect 30101 25851 30159 25857
rect 23716 25792 27476 25820
rect 27617 25823 27675 25829
rect 23716 25780 23722 25792
rect 27617 25789 27629 25823
rect 27663 25820 27675 25823
rect 27982 25820 27988 25832
rect 27663 25792 27988 25820
rect 27663 25789 27675 25792
rect 27617 25783 27675 25789
rect 27982 25780 27988 25792
rect 28040 25820 28046 25832
rect 29270 25820 29276 25832
rect 28040 25792 29276 25820
rect 28040 25780 28046 25792
rect 29270 25780 29276 25792
rect 29328 25820 29334 25832
rect 30843 25820 30871 25860
rect 31478 25848 31484 25860
rect 31536 25848 31542 25900
rect 31769 25891 31827 25897
rect 31769 25857 31781 25891
rect 31815 25888 31827 25891
rect 32122 25888 32128 25900
rect 31815 25860 32128 25888
rect 31815 25857 31827 25860
rect 31769 25851 31827 25857
rect 32122 25848 32128 25860
rect 32180 25848 32186 25900
rect 32214 25848 32220 25900
rect 32272 25888 32278 25900
rect 32309 25891 32367 25897
rect 32309 25888 32321 25891
rect 32272 25860 32321 25888
rect 32272 25848 32278 25860
rect 32309 25857 32321 25860
rect 32355 25857 32367 25891
rect 32309 25851 32367 25857
rect 33873 25891 33931 25897
rect 33873 25857 33885 25891
rect 33919 25888 33931 25891
rect 34606 25888 34612 25900
rect 33919 25860 34612 25888
rect 33919 25857 33931 25860
rect 33873 25851 33931 25857
rect 34606 25848 34612 25860
rect 34664 25848 34670 25900
rect 38286 25888 38292 25900
rect 35636 25860 38292 25888
rect 32232 25820 32260 25848
rect 29328 25792 30788 25820
rect 30843 25792 32260 25820
rect 34149 25823 34207 25829
rect 29328 25780 29334 25792
rect 25038 25752 25044 25764
rect 21008 25724 25044 25752
rect 25038 25712 25044 25724
rect 25096 25712 25102 25764
rect 30190 25712 30196 25764
rect 30248 25752 30254 25764
rect 30760 25752 30788 25792
rect 34149 25789 34161 25823
rect 34195 25820 34207 25823
rect 34238 25820 34244 25832
rect 34195 25792 34244 25820
rect 34195 25789 34207 25792
rect 34149 25783 34207 25789
rect 34238 25780 34244 25792
rect 34296 25780 34302 25832
rect 35345 25823 35403 25829
rect 35345 25789 35357 25823
rect 35391 25820 35403 25823
rect 35434 25820 35440 25832
rect 35391 25792 35440 25820
rect 35391 25789 35403 25792
rect 35345 25783 35403 25789
rect 35434 25780 35440 25792
rect 35492 25780 35498 25832
rect 33502 25752 33508 25764
rect 30248 25724 30696 25752
rect 30760 25724 33508 25752
rect 30248 25712 30254 25724
rect 22462 25684 22468 25696
rect 18340 25656 22468 25684
rect 22462 25644 22468 25656
rect 22520 25644 22526 25696
rect 27522 25684 27528 25696
rect 27483 25656 27528 25684
rect 27522 25644 27528 25656
rect 27580 25684 27586 25696
rect 28261 25687 28319 25693
rect 28261 25684 28273 25687
rect 27580 25656 28273 25684
rect 27580 25644 27586 25656
rect 28261 25653 28273 25656
rect 28307 25653 28319 25687
rect 28261 25647 28319 25653
rect 30285 25687 30343 25693
rect 30285 25653 30297 25687
rect 30331 25684 30343 25687
rect 30466 25684 30472 25696
rect 30331 25656 30472 25684
rect 30331 25653 30343 25656
rect 30285 25647 30343 25653
rect 30466 25644 30472 25656
rect 30524 25644 30530 25696
rect 30668 25684 30696 25724
rect 33502 25712 33508 25724
rect 33560 25712 33566 25764
rect 31665 25687 31723 25693
rect 31665 25684 31677 25687
rect 30668 25656 31677 25684
rect 31665 25653 31677 25656
rect 31711 25653 31723 25687
rect 31665 25647 31723 25653
rect 32398 25644 32404 25696
rect 32456 25684 32462 25696
rect 32493 25687 32551 25693
rect 32493 25684 32505 25687
rect 32456 25656 32505 25684
rect 32456 25644 32462 25656
rect 32493 25653 32505 25656
rect 32539 25684 32551 25687
rect 35636 25684 35664 25860
rect 38286 25848 38292 25860
rect 38344 25848 38350 25900
rect 38378 25848 38384 25900
rect 38436 25888 38442 25900
rect 38562 25888 38568 25900
rect 38436 25860 38568 25888
rect 38436 25848 38442 25860
rect 38562 25848 38568 25860
rect 38620 25848 38626 25900
rect 38746 25888 38752 25900
rect 38707 25860 38752 25888
rect 38746 25848 38752 25860
rect 38804 25848 38810 25900
rect 47762 25888 47768 25900
rect 47723 25860 47768 25888
rect 47762 25848 47768 25860
rect 47820 25848 47826 25900
rect 37274 25780 37280 25832
rect 37332 25820 37338 25832
rect 38102 25820 38108 25832
rect 37332 25792 38108 25820
rect 37332 25780 37338 25792
rect 38102 25780 38108 25792
rect 38160 25820 38166 25832
rect 39301 25823 39359 25829
rect 39301 25820 39313 25823
rect 38160 25792 39313 25820
rect 38160 25780 38166 25792
rect 39301 25789 39313 25792
rect 39347 25789 39359 25823
rect 39301 25783 39359 25789
rect 36538 25752 36544 25764
rect 36188 25724 36544 25752
rect 36188 25693 36216 25724
rect 36538 25712 36544 25724
rect 36596 25752 36602 25764
rect 36722 25752 36728 25764
rect 36596 25724 36728 25752
rect 36596 25712 36602 25724
rect 36722 25712 36728 25724
rect 36780 25712 36786 25764
rect 32539 25656 35664 25684
rect 36173 25687 36231 25693
rect 32539 25653 32551 25656
rect 32493 25647 32551 25653
rect 36173 25653 36185 25687
rect 36219 25653 36231 25687
rect 36173 25647 36231 25653
rect 36357 25687 36415 25693
rect 36357 25653 36369 25687
rect 36403 25684 36415 25687
rect 36906 25684 36912 25696
rect 36403 25656 36912 25684
rect 36403 25653 36415 25656
rect 36357 25647 36415 25653
rect 36906 25644 36912 25656
rect 36964 25644 36970 25696
rect 38105 25687 38163 25693
rect 38105 25653 38117 25687
rect 38151 25684 38163 25687
rect 38194 25684 38200 25696
rect 38151 25656 38200 25684
rect 38151 25653 38163 25656
rect 38105 25647 38163 25653
rect 38194 25644 38200 25656
rect 38252 25644 38258 25696
rect 46474 25644 46480 25696
rect 46532 25684 46538 25696
rect 47213 25687 47271 25693
rect 47213 25684 47225 25687
rect 46532 25656 47225 25684
rect 46532 25644 46538 25656
rect 47213 25653 47225 25656
rect 47259 25653 47271 25687
rect 47213 25647 47271 25653
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 13449 25483 13507 25489
rect 13449 25449 13461 25483
rect 13495 25480 13507 25483
rect 13630 25480 13636 25492
rect 13495 25452 13636 25480
rect 13495 25449 13507 25452
rect 13449 25443 13507 25449
rect 13630 25440 13636 25452
rect 13688 25440 13694 25492
rect 16209 25483 16267 25489
rect 16209 25449 16221 25483
rect 16255 25480 16267 25483
rect 16574 25480 16580 25492
rect 16255 25452 16580 25480
rect 16255 25449 16267 25452
rect 16209 25443 16267 25449
rect 16574 25440 16580 25452
rect 16632 25440 16638 25492
rect 17310 25440 17316 25492
rect 17368 25480 17374 25492
rect 18782 25480 18788 25492
rect 17368 25452 18788 25480
rect 17368 25440 17374 25452
rect 18782 25440 18788 25452
rect 18840 25440 18846 25492
rect 20806 25440 20812 25492
rect 20864 25480 20870 25492
rect 21910 25480 21916 25492
rect 20864 25452 21916 25480
rect 20864 25440 20870 25452
rect 21910 25440 21916 25452
rect 21968 25480 21974 25492
rect 24946 25480 24952 25492
rect 21968 25452 24952 25480
rect 21968 25440 21974 25452
rect 24946 25440 24952 25452
rect 25004 25480 25010 25492
rect 25685 25483 25743 25489
rect 25685 25480 25697 25483
rect 25004 25452 25697 25480
rect 25004 25440 25010 25452
rect 25685 25449 25697 25452
rect 25731 25449 25743 25483
rect 32490 25480 32496 25492
rect 32451 25452 32496 25480
rect 25685 25443 25743 25449
rect 32490 25440 32496 25452
rect 32548 25440 32554 25492
rect 18230 25372 18236 25424
rect 18288 25412 18294 25424
rect 27522 25412 27528 25424
rect 18288 25384 27528 25412
rect 18288 25372 18294 25384
rect 27522 25372 27528 25384
rect 27580 25412 27586 25424
rect 31018 25412 31024 25424
rect 27580 25384 31024 25412
rect 27580 25372 27586 25384
rect 31018 25372 31024 25384
rect 31076 25372 31082 25424
rect 1762 25344 1768 25356
rect 1723 25316 1768 25344
rect 1762 25304 1768 25316
rect 1820 25304 1826 25356
rect 2774 25304 2780 25356
rect 2832 25344 2838 25356
rect 2832 25316 2877 25344
rect 2832 25304 2838 25316
rect 11974 25304 11980 25356
rect 12032 25344 12038 25356
rect 12069 25347 12127 25353
rect 12069 25344 12081 25347
rect 12032 25316 12081 25344
rect 12032 25304 12038 25316
rect 12069 25313 12081 25316
rect 12115 25313 12127 25347
rect 18877 25347 18935 25353
rect 18877 25344 18889 25347
rect 12069 25307 12127 25313
rect 17604 25316 18889 25344
rect 1578 25276 1584 25288
rect 1539 25248 1584 25276
rect 1578 25236 1584 25248
rect 1636 25236 1642 25288
rect 12084 25276 12112 25307
rect 17604 25288 17632 25316
rect 18877 25313 18889 25316
rect 18923 25313 18935 25347
rect 18877 25307 18935 25313
rect 19334 25304 19340 25356
rect 19392 25344 19398 25356
rect 23658 25344 23664 25356
rect 19392 25316 20116 25344
rect 23619 25316 23664 25344
rect 19392 25304 19398 25316
rect 13814 25276 13820 25288
rect 12084 25248 13820 25276
rect 13814 25236 13820 25248
rect 13872 25276 13878 25288
rect 14826 25276 14832 25288
rect 13872 25248 14832 25276
rect 13872 25236 13878 25248
rect 14826 25236 14832 25248
rect 14884 25236 14890 25288
rect 16850 25276 16856 25288
rect 16811 25248 16856 25276
rect 16850 25236 16856 25248
rect 16908 25236 16914 25288
rect 17034 25276 17040 25288
rect 16995 25248 17040 25276
rect 17034 25236 17040 25248
rect 17092 25236 17098 25288
rect 17129 25279 17187 25285
rect 17129 25245 17141 25279
rect 17175 25276 17187 25279
rect 17586 25276 17592 25288
rect 17175 25248 17592 25276
rect 17175 25245 17187 25248
rect 17129 25239 17187 25245
rect 17586 25236 17592 25248
rect 17644 25236 17650 25288
rect 18601 25279 18659 25285
rect 18601 25245 18613 25279
rect 18647 25245 18659 25279
rect 18601 25239 18659 25245
rect 12342 25217 12348 25220
rect 12336 25208 12348 25217
rect 12303 25180 12348 25208
rect 12336 25171 12348 25180
rect 12342 25168 12348 25171
rect 12400 25168 12406 25220
rect 15096 25211 15154 25217
rect 15096 25177 15108 25211
rect 15142 25208 15154 25211
rect 16669 25211 16727 25217
rect 16669 25208 16681 25211
rect 15142 25180 16681 25208
rect 15142 25177 15154 25180
rect 15096 25171 15154 25177
rect 16669 25177 16681 25180
rect 16715 25177 16727 25211
rect 18616 25208 18644 25239
rect 19242 25236 19248 25288
rect 19300 25276 19306 25288
rect 19613 25279 19671 25285
rect 19613 25276 19625 25279
rect 19300 25248 19625 25276
rect 19300 25236 19306 25248
rect 19613 25245 19625 25248
rect 19659 25245 19671 25279
rect 19613 25239 19671 25245
rect 19889 25279 19947 25285
rect 19889 25245 19901 25279
rect 19935 25276 19947 25279
rect 19978 25276 19984 25288
rect 19935 25248 19984 25276
rect 19935 25245 19947 25248
rect 19889 25239 19947 25245
rect 19429 25211 19487 25217
rect 19429 25208 19441 25211
rect 18616 25180 19441 25208
rect 16669 25171 16727 25177
rect 19429 25177 19441 25180
rect 19475 25177 19487 25211
rect 19628 25208 19656 25239
rect 19978 25236 19984 25248
rect 20036 25236 20042 25288
rect 20088 25285 20116 25316
rect 23658 25304 23664 25316
rect 23716 25304 23722 25356
rect 24949 25347 25007 25353
rect 24949 25313 24961 25347
rect 24995 25344 25007 25347
rect 29362 25344 29368 25356
rect 24995 25316 29368 25344
rect 24995 25313 25007 25316
rect 24949 25307 25007 25313
rect 20073 25279 20131 25285
rect 20073 25245 20085 25279
rect 20119 25245 20131 25279
rect 20073 25239 20131 25245
rect 21358 25236 21364 25288
rect 21416 25276 21422 25288
rect 21545 25279 21603 25285
rect 21545 25276 21557 25279
rect 21416 25248 21557 25276
rect 21416 25236 21422 25248
rect 21545 25245 21557 25248
rect 21591 25245 21603 25279
rect 22370 25276 22376 25288
rect 21545 25239 21603 25245
rect 22066 25248 22376 25276
rect 20806 25208 20812 25220
rect 19628 25180 20812 25208
rect 19429 25171 19487 25177
rect 20806 25168 20812 25180
rect 20864 25168 20870 25220
rect 22066 25208 22094 25248
rect 22370 25236 22376 25248
rect 22428 25276 22434 25288
rect 24964 25276 24992 25307
rect 29362 25304 29368 25316
rect 29420 25304 29426 25356
rect 36170 25344 36176 25356
rect 35636 25316 36176 25344
rect 22428 25248 24992 25276
rect 25501 25279 25559 25285
rect 22428 25236 22434 25248
rect 25501 25245 25513 25279
rect 25547 25276 25559 25279
rect 25682 25276 25688 25288
rect 25547 25248 25688 25276
rect 25547 25245 25559 25248
rect 25501 25239 25559 25245
rect 25682 25236 25688 25248
rect 25740 25276 25746 25288
rect 27706 25276 27712 25288
rect 25740 25248 27712 25276
rect 25740 25236 25746 25248
rect 27706 25236 27712 25248
rect 27764 25276 27770 25288
rect 28350 25276 28356 25288
rect 27764 25248 28356 25276
rect 27764 25236 27770 25248
rect 28350 25236 28356 25248
rect 28408 25236 28414 25288
rect 30098 25276 30104 25288
rect 30059 25248 30104 25276
rect 30098 25236 30104 25248
rect 30156 25236 30162 25288
rect 30190 25236 30196 25288
rect 30248 25276 30254 25288
rect 30285 25279 30343 25285
rect 30285 25276 30297 25279
rect 30248 25248 30297 25276
rect 30248 25236 30254 25248
rect 30285 25245 30297 25248
rect 30331 25245 30343 25279
rect 30285 25239 30343 25245
rect 30377 25279 30435 25285
rect 30377 25245 30389 25279
rect 30423 25276 30435 25279
rect 30834 25276 30840 25288
rect 30423 25248 30840 25276
rect 30423 25245 30435 25248
rect 30377 25239 30435 25245
rect 30834 25236 30840 25248
rect 30892 25236 30898 25288
rect 31113 25279 31171 25285
rect 31113 25245 31125 25279
rect 31159 25276 31171 25279
rect 33778 25276 33784 25288
rect 31159 25248 33784 25276
rect 31159 25245 31171 25248
rect 31113 25239 31171 25245
rect 33778 25236 33784 25248
rect 33836 25236 33842 25288
rect 35636 25285 35664 25316
rect 36170 25304 36176 25316
rect 36228 25304 36234 25356
rect 36446 25344 36452 25356
rect 36407 25316 36452 25344
rect 36446 25304 36452 25316
rect 36504 25304 36510 25356
rect 46474 25344 46480 25356
rect 46435 25316 46480 25344
rect 46474 25304 46480 25316
rect 46532 25304 46538 25356
rect 48222 25344 48228 25356
rect 48183 25316 48228 25344
rect 48222 25304 48228 25316
rect 48280 25304 48286 25356
rect 35621 25279 35679 25285
rect 35621 25245 35633 25279
rect 35667 25245 35679 25279
rect 35621 25239 35679 25245
rect 35805 25279 35863 25285
rect 35805 25245 35817 25279
rect 35851 25245 35863 25279
rect 36354 25276 36360 25288
rect 36315 25248 36360 25276
rect 35805 25239 35863 25245
rect 20916 25180 22094 25208
rect 23385 25211 23443 25217
rect 18414 25140 18420 25152
rect 18375 25112 18420 25140
rect 18414 25100 18420 25112
rect 18472 25100 18478 25152
rect 18782 25100 18788 25152
rect 18840 25140 18846 25152
rect 20916 25140 20944 25180
rect 23385 25177 23397 25211
rect 23431 25208 23443 25211
rect 23658 25208 23664 25220
rect 23431 25180 23664 25208
rect 23431 25177 23443 25180
rect 23385 25171 23443 25177
rect 23658 25168 23664 25180
rect 23716 25168 23722 25220
rect 24578 25168 24584 25220
rect 24636 25208 24642 25220
rect 31386 25217 31392 25220
rect 24673 25211 24731 25217
rect 24673 25208 24685 25211
rect 24636 25180 24685 25208
rect 24636 25168 24642 25180
rect 24673 25177 24685 25180
rect 24719 25177 24731 25211
rect 24673 25171 24731 25177
rect 31380 25171 31392 25217
rect 31444 25208 31450 25220
rect 35820 25208 35848 25239
rect 36354 25236 36360 25248
rect 36412 25236 36418 25288
rect 36906 25276 36912 25288
rect 36867 25248 36912 25276
rect 36906 25236 36912 25248
rect 36964 25236 36970 25288
rect 37274 25236 37280 25288
rect 37332 25276 37338 25288
rect 37645 25279 37703 25285
rect 37645 25276 37657 25279
rect 37332 25248 37657 25276
rect 37332 25236 37338 25248
rect 37645 25245 37657 25248
rect 37691 25245 37703 25279
rect 37645 25239 37703 25245
rect 36446 25208 36452 25220
rect 31444 25180 31480 25208
rect 35820 25180 36452 25208
rect 31386 25168 31392 25171
rect 31444 25168 31450 25180
rect 36446 25168 36452 25180
rect 36504 25168 36510 25220
rect 36817 25211 36875 25217
rect 36817 25177 36829 25211
rect 36863 25177 36875 25211
rect 36817 25171 36875 25177
rect 37912 25211 37970 25217
rect 37912 25177 37924 25211
rect 37958 25208 37970 25211
rect 38010 25208 38016 25220
rect 37958 25180 38016 25208
rect 37958 25177 37970 25180
rect 37912 25171 37970 25177
rect 21634 25140 21640 25152
rect 18840 25112 20944 25140
rect 21595 25112 21640 25140
rect 18840 25100 18846 25112
rect 21634 25100 21640 25112
rect 21692 25100 21698 25152
rect 27890 25140 27896 25152
rect 27851 25112 27896 25140
rect 27890 25100 27896 25112
rect 27948 25140 27954 25152
rect 28718 25140 28724 25152
rect 27948 25112 28724 25140
rect 27948 25100 27954 25112
rect 28718 25100 28724 25112
rect 28776 25100 28782 25152
rect 29914 25140 29920 25152
rect 29875 25112 29920 25140
rect 29914 25100 29920 25112
rect 29972 25100 29978 25152
rect 34146 25100 34152 25152
rect 34204 25140 34210 25152
rect 36832 25140 36860 25171
rect 38010 25168 38016 25180
rect 38068 25168 38074 25220
rect 46661 25211 46719 25217
rect 46661 25177 46673 25211
rect 46707 25208 46719 25211
rect 47118 25208 47124 25220
rect 46707 25180 47124 25208
rect 46707 25177 46719 25180
rect 46661 25171 46719 25177
rect 47118 25168 47124 25180
rect 47176 25168 47182 25220
rect 34204 25112 36860 25140
rect 34204 25100 34210 25112
rect 38470 25100 38476 25152
rect 38528 25140 38534 25152
rect 39025 25143 39083 25149
rect 39025 25140 39037 25143
rect 38528 25112 39037 25140
rect 38528 25100 38534 25112
rect 39025 25109 39037 25112
rect 39071 25109 39083 25143
rect 39025 25103 39083 25109
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 12342 24936 12348 24948
rect 12303 24908 12348 24936
rect 12342 24896 12348 24908
rect 12400 24896 12406 24948
rect 17586 24896 17592 24948
rect 17644 24936 17650 24948
rect 17644 24908 19288 24936
rect 17644 24896 17650 24908
rect 18414 24877 18420 24880
rect 18408 24868 18420 24877
rect 16224 24840 16436 24868
rect 18375 24840 18420 24868
rect 1578 24760 1584 24812
rect 1636 24800 1642 24812
rect 2225 24803 2283 24809
rect 2225 24800 2237 24803
rect 1636 24772 2237 24800
rect 1636 24760 1642 24772
rect 2225 24769 2237 24772
rect 2271 24769 2283 24803
rect 12526 24800 12532 24812
rect 12487 24772 12532 24800
rect 2225 24763 2283 24769
rect 12526 24760 12532 24772
rect 12584 24760 12590 24812
rect 13814 24800 13820 24812
rect 13775 24772 13820 24800
rect 13814 24760 13820 24772
rect 13872 24760 13878 24812
rect 14084 24803 14142 24809
rect 14084 24769 14096 24803
rect 14130 24800 14142 24803
rect 14366 24800 14372 24812
rect 14130 24772 14372 24800
rect 14130 24769 14142 24772
rect 14084 24763 14142 24769
rect 14366 24760 14372 24772
rect 14424 24760 14430 24812
rect 15838 24800 15844 24812
rect 15799 24772 15844 24800
rect 15838 24760 15844 24772
rect 15896 24760 15902 24812
rect 16117 24803 16175 24809
rect 16117 24769 16129 24803
rect 16163 24800 16175 24803
rect 16224 24800 16252 24840
rect 16163 24772 16252 24800
rect 16301 24803 16359 24809
rect 16163 24769 16175 24772
rect 16117 24763 16175 24769
rect 16301 24769 16313 24803
rect 16347 24769 16359 24803
rect 16408 24800 16436 24840
rect 18408 24831 18420 24840
rect 18414 24828 18420 24831
rect 18472 24828 18478 24880
rect 19260 24868 19288 24908
rect 19334 24896 19340 24948
rect 19392 24936 19398 24948
rect 19521 24939 19579 24945
rect 19521 24936 19533 24939
rect 19392 24908 19533 24936
rect 19392 24896 19398 24908
rect 19521 24905 19533 24908
rect 19567 24905 19579 24939
rect 19521 24899 19579 24905
rect 21361 24939 21419 24945
rect 21361 24905 21373 24939
rect 21407 24936 21419 24939
rect 21634 24936 21640 24948
rect 21407 24908 21640 24936
rect 21407 24905 21419 24908
rect 21361 24899 21419 24905
rect 21634 24896 21640 24908
rect 21692 24896 21698 24948
rect 21744 24908 27660 24936
rect 21744 24868 21772 24908
rect 19260 24840 21772 24868
rect 23486 24871 23544 24877
rect 23486 24837 23498 24871
rect 23532 24837 23544 24871
rect 23486 24831 23544 24837
rect 24136 24840 24440 24868
rect 19978 24800 19984 24812
rect 16408 24772 19984 24800
rect 16301 24763 16359 24769
rect 12802 24732 12808 24744
rect 12763 24704 12808 24732
rect 12802 24692 12808 24704
rect 12860 24692 12866 24744
rect 16316 24732 16344 24763
rect 19978 24760 19984 24772
rect 20036 24760 20042 24812
rect 20254 24760 20260 24812
rect 20312 24800 20318 24812
rect 21177 24803 21235 24809
rect 21177 24800 21189 24803
rect 20312 24772 21189 24800
rect 20312 24760 20318 24772
rect 21177 24769 21189 24772
rect 21223 24769 21235 24803
rect 21177 24763 21235 24769
rect 21453 24803 21511 24809
rect 21453 24769 21465 24803
rect 21499 24800 21511 24803
rect 22094 24800 22100 24812
rect 21499 24772 22100 24800
rect 21499 24769 21511 24772
rect 21453 24763 21511 24769
rect 22094 24760 22100 24772
rect 22152 24760 22158 24812
rect 22189 24803 22247 24809
rect 22189 24769 22201 24803
rect 22235 24769 22247 24803
rect 22370 24800 22376 24812
rect 22331 24772 22376 24800
rect 22189 24763 22247 24769
rect 18138 24732 18144 24744
rect 15304 24704 16344 24732
rect 18099 24704 18144 24732
rect 15304 24676 15332 24704
rect 18138 24692 18144 24704
rect 18196 24692 18202 24744
rect 15197 24667 15255 24673
rect 15197 24633 15209 24667
rect 15243 24664 15255 24667
rect 15286 24664 15292 24676
rect 15243 24636 15292 24664
rect 15243 24633 15255 24636
rect 15197 24627 15255 24633
rect 15286 24624 15292 24636
rect 15344 24624 15350 24676
rect 17034 24664 17040 24676
rect 15488 24636 17040 24664
rect 12713 24599 12771 24605
rect 12713 24565 12725 24599
rect 12759 24596 12771 24599
rect 15488 24596 15516 24636
rect 17034 24624 17040 24636
rect 17092 24624 17098 24676
rect 21177 24667 21235 24673
rect 21177 24633 21189 24667
rect 21223 24664 21235 24667
rect 22204 24664 22232 24763
rect 22370 24760 22376 24772
rect 22428 24760 22434 24812
rect 23106 24800 23112 24812
rect 23067 24772 23112 24800
rect 23106 24760 23112 24772
rect 23164 24760 23170 24812
rect 23198 24760 23204 24812
rect 23256 24800 23262 24812
rect 23492 24800 23520 24831
rect 23750 24800 23756 24812
rect 23256 24772 23520 24800
rect 23711 24772 23756 24800
rect 23256 24760 23262 24772
rect 23750 24760 23756 24772
rect 23808 24760 23814 24812
rect 22462 24732 22468 24744
rect 22375 24704 22468 24732
rect 22462 24692 22468 24704
rect 22520 24732 22526 24744
rect 24136 24732 24164 24840
rect 24210 24760 24216 24812
rect 24268 24800 24274 24812
rect 24305 24803 24363 24809
rect 24305 24800 24317 24803
rect 24268 24772 24317 24800
rect 24268 24760 24274 24772
rect 24305 24769 24317 24772
rect 24351 24769 24363 24803
rect 24412 24800 24440 24840
rect 25332 24840 26280 24868
rect 25332 24800 25360 24840
rect 24412 24772 25360 24800
rect 25400 24803 25458 24809
rect 24305 24763 24363 24769
rect 25400 24769 25412 24803
rect 25446 24800 25458 24803
rect 25682 24800 25688 24812
rect 25446 24772 25688 24800
rect 25446 24769 25458 24772
rect 25400 24763 25458 24769
rect 25682 24760 25688 24772
rect 25740 24760 25746 24812
rect 25866 24760 25872 24812
rect 25924 24800 25930 24812
rect 25924 24772 26188 24800
rect 25924 24760 25930 24772
rect 24394 24732 24400 24744
rect 22520 24704 24164 24732
rect 24355 24704 24400 24732
rect 22520 24692 22526 24704
rect 24394 24692 24400 24704
rect 24452 24692 24458 24744
rect 25133 24735 25191 24741
rect 25133 24701 25145 24735
rect 25179 24701 25191 24735
rect 25133 24695 25191 24701
rect 24762 24664 24768 24676
rect 21223 24636 22232 24664
rect 24504 24636 24768 24664
rect 21223 24633 21235 24636
rect 21177 24627 21235 24633
rect 15654 24596 15660 24608
rect 12759 24568 15516 24596
rect 15615 24568 15660 24596
rect 12759 24565 12771 24568
rect 12713 24559 12771 24565
rect 15654 24556 15660 24568
rect 15712 24556 15718 24608
rect 22002 24596 22008 24608
rect 21963 24568 22008 24596
rect 22002 24556 22008 24568
rect 22060 24556 22066 24608
rect 23382 24556 23388 24608
rect 23440 24596 23446 24608
rect 24504 24605 24532 24636
rect 24762 24624 24768 24636
rect 24820 24624 24826 24676
rect 23477 24599 23535 24605
rect 23477 24596 23489 24599
rect 23440 24568 23489 24596
rect 23440 24556 23446 24568
rect 23477 24565 23489 24568
rect 23523 24565 23535 24599
rect 23477 24559 23535 24565
rect 24489 24599 24547 24605
rect 24489 24565 24501 24599
rect 24535 24565 24547 24599
rect 24670 24596 24676 24608
rect 24631 24568 24676 24596
rect 24489 24559 24547 24565
rect 24670 24556 24676 24568
rect 24728 24556 24734 24608
rect 25148 24596 25176 24695
rect 26160 24664 26188 24772
rect 26252 24732 26280 24840
rect 27632 24812 27660 24908
rect 29638 24896 29644 24948
rect 29696 24936 29702 24948
rect 31297 24939 31355 24945
rect 29696 24908 31248 24936
rect 29696 24896 29702 24908
rect 29724 24871 29782 24877
rect 29724 24837 29736 24871
rect 29770 24868 29782 24871
rect 29914 24868 29920 24880
rect 29770 24840 29920 24868
rect 29770 24837 29782 24840
rect 29724 24831 29782 24837
rect 29914 24828 29920 24840
rect 29972 24828 29978 24880
rect 27341 24803 27399 24809
rect 27341 24769 27353 24803
rect 27387 24800 27399 24803
rect 27522 24800 27528 24812
rect 27387 24772 27528 24800
rect 27387 24769 27399 24772
rect 27341 24763 27399 24769
rect 27522 24760 27528 24772
rect 27580 24760 27586 24812
rect 27614 24760 27620 24812
rect 27672 24800 27678 24812
rect 30650 24800 30656 24812
rect 27672 24772 27765 24800
rect 27816 24772 30656 24800
rect 27672 24760 27678 24772
rect 27816 24732 27844 24772
rect 30650 24760 30656 24772
rect 30708 24760 30714 24812
rect 29454 24732 29460 24744
rect 26252 24704 27844 24732
rect 29415 24704 29460 24732
rect 29454 24692 29460 24704
rect 29512 24692 29518 24744
rect 31220 24732 31248 24908
rect 31297 24905 31309 24939
rect 31343 24936 31355 24939
rect 31386 24936 31392 24948
rect 31343 24908 31392 24936
rect 31343 24905 31355 24908
rect 31297 24899 31355 24905
rect 31386 24896 31392 24908
rect 31444 24896 31450 24948
rect 32490 24896 32496 24948
rect 32548 24896 32554 24948
rect 38010 24936 38016 24948
rect 37971 24908 38016 24936
rect 38010 24896 38016 24908
rect 38068 24896 38074 24948
rect 32508 24868 32536 24896
rect 36173 24871 36231 24877
rect 32508 24840 32904 24868
rect 31481 24803 31539 24809
rect 31481 24769 31493 24803
rect 31527 24800 31539 24803
rect 32309 24803 32367 24809
rect 32309 24800 32321 24803
rect 31527 24772 32321 24800
rect 31527 24769 31539 24772
rect 31481 24763 31539 24769
rect 32309 24769 32321 24772
rect 32355 24769 32367 24803
rect 32309 24763 32367 24769
rect 32493 24803 32551 24809
rect 32493 24769 32505 24803
rect 32539 24769 32551 24803
rect 32766 24800 32772 24812
rect 32727 24772 32772 24800
rect 32493 24763 32551 24769
rect 31662 24732 31668 24744
rect 31220 24704 31668 24732
rect 31662 24692 31668 24704
rect 31720 24692 31726 24744
rect 31754 24692 31760 24744
rect 31812 24732 31818 24744
rect 32508 24732 32536 24763
rect 32766 24760 32772 24772
rect 32824 24760 32830 24812
rect 32876 24809 32904 24840
rect 33520 24840 33732 24868
rect 32870 24803 32928 24809
rect 32870 24769 32882 24803
rect 32916 24769 32928 24803
rect 32870 24763 32928 24769
rect 33134 24760 33140 24812
rect 33192 24800 33198 24812
rect 33520 24800 33548 24840
rect 33192 24772 33548 24800
rect 33597 24803 33655 24809
rect 33192 24760 33198 24772
rect 33597 24769 33609 24803
rect 33643 24769 33655 24803
rect 33704 24800 33732 24840
rect 36173 24837 36185 24871
rect 36219 24868 36231 24871
rect 36354 24868 36360 24880
rect 36219 24840 36360 24868
rect 36219 24837 36231 24840
rect 36173 24831 36231 24837
rect 36354 24828 36360 24840
rect 36412 24868 36418 24880
rect 37366 24868 37372 24880
rect 36412 24840 37372 24868
rect 36412 24828 36418 24840
rect 37366 24828 37372 24840
rect 37424 24828 37430 24880
rect 47394 24828 47400 24880
rect 47452 24868 47458 24880
rect 47762 24868 47768 24880
rect 47452 24840 47768 24868
rect 47452 24828 47458 24840
rect 47762 24828 47768 24840
rect 47820 24828 47826 24880
rect 33870 24800 33876 24812
rect 33704 24772 33876 24800
rect 33597 24763 33655 24769
rect 33612 24732 33640 24763
rect 33870 24760 33876 24772
rect 33928 24760 33934 24812
rect 34054 24800 34060 24812
rect 34015 24772 34060 24800
rect 34054 24760 34060 24772
rect 34112 24760 34118 24812
rect 35710 24760 35716 24812
rect 35768 24800 35774 24812
rect 35805 24803 35863 24809
rect 35805 24800 35817 24803
rect 35768 24772 35817 24800
rect 35768 24760 35774 24772
rect 35805 24769 35817 24772
rect 35851 24769 35863 24803
rect 35986 24800 35992 24812
rect 35947 24772 35992 24800
rect 35805 24763 35863 24769
rect 35986 24760 35992 24772
rect 36044 24760 36050 24812
rect 36265 24803 36323 24809
rect 36265 24769 36277 24803
rect 36311 24800 36323 24803
rect 36446 24800 36452 24812
rect 36311 24772 36452 24800
rect 36311 24769 36323 24772
rect 36265 24763 36323 24769
rect 36446 24760 36452 24772
rect 36504 24760 36510 24812
rect 36722 24800 36728 24812
rect 36683 24772 36728 24800
rect 36722 24760 36728 24772
rect 36780 24760 36786 24812
rect 36909 24803 36967 24809
rect 36909 24769 36921 24803
rect 36955 24769 36967 24803
rect 38194 24800 38200 24812
rect 38155 24772 38200 24800
rect 36909 24763 36967 24769
rect 33962 24732 33968 24744
rect 31812 24704 31857 24732
rect 32508 24704 33968 24732
rect 31812 24692 31818 24704
rect 33962 24692 33968 24704
rect 34020 24692 34026 24744
rect 36078 24692 36084 24744
rect 36136 24732 36142 24744
rect 36924 24732 36952 24763
rect 38194 24760 38200 24772
rect 38252 24760 38258 24812
rect 47026 24800 47032 24812
rect 46987 24772 47032 24800
rect 47026 24760 47032 24772
rect 47084 24760 47090 24812
rect 47118 24760 47124 24812
rect 47176 24800 47182 24812
rect 48133 24803 48191 24809
rect 47176 24772 47221 24800
rect 47176 24760 47182 24772
rect 48133 24769 48145 24803
rect 48179 24800 48191 24803
rect 48222 24800 48228 24812
rect 48179 24772 48228 24800
rect 48179 24769 48191 24772
rect 48133 24763 48191 24769
rect 48222 24760 48228 24772
rect 48280 24760 48286 24812
rect 38470 24732 38476 24744
rect 36136 24704 38476 24732
rect 36136 24692 36142 24704
rect 38470 24692 38476 24704
rect 38528 24692 38534 24744
rect 26513 24667 26571 24673
rect 26513 24664 26525 24667
rect 26160 24636 26525 24664
rect 26513 24633 26525 24636
rect 26559 24633 26571 24667
rect 46842 24664 46848 24676
rect 26513 24627 26571 24633
rect 30760 24636 46848 24664
rect 26234 24596 26240 24608
rect 25148 24568 26240 24596
rect 26234 24556 26240 24568
rect 26292 24556 26298 24608
rect 27154 24596 27160 24608
rect 27115 24568 27160 24596
rect 27154 24556 27160 24568
rect 27212 24556 27218 24608
rect 27525 24599 27583 24605
rect 27525 24565 27537 24599
rect 27571 24596 27583 24599
rect 29638 24596 29644 24608
rect 27571 24568 29644 24596
rect 27571 24565 27583 24568
rect 27525 24559 27583 24565
rect 29638 24556 29644 24568
rect 29696 24556 29702 24608
rect 29730 24556 29736 24608
rect 29788 24596 29794 24608
rect 30760 24596 30788 24636
rect 46842 24624 46848 24636
rect 46900 24624 46906 24676
rect 29788 24568 30788 24596
rect 29788 24556 29794 24568
rect 30834 24556 30840 24608
rect 30892 24596 30898 24608
rect 30892 24568 30937 24596
rect 30892 24556 30898 24568
rect 32766 24556 32772 24608
rect 32824 24596 32830 24608
rect 33413 24599 33471 24605
rect 33413 24596 33425 24599
rect 32824 24568 33425 24596
rect 32824 24556 32830 24568
rect 33413 24565 33425 24568
rect 33459 24565 33471 24599
rect 33413 24559 33471 24565
rect 36354 24556 36360 24608
rect 36412 24596 36418 24608
rect 36725 24599 36783 24605
rect 36725 24596 36737 24599
rect 36412 24568 36737 24596
rect 36412 24556 36418 24568
rect 36725 24565 36737 24568
rect 36771 24565 36783 24599
rect 38378 24596 38384 24608
rect 38339 24568 38384 24596
rect 36725 24559 36783 24565
rect 38378 24556 38384 24568
rect 38436 24596 38442 24608
rect 38838 24596 38844 24608
rect 38436 24568 38844 24596
rect 38436 24556 38442 24568
rect 38838 24556 38844 24568
rect 38896 24556 38902 24608
rect 46934 24556 46940 24608
rect 46992 24596 46998 24608
rect 48225 24599 48283 24605
rect 48225 24596 48237 24599
rect 46992 24568 48237 24596
rect 46992 24556 46998 24568
rect 48225 24565 48237 24568
rect 48271 24565 48283 24599
rect 48225 24559 48283 24565
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 14366 24392 14372 24404
rect 14327 24364 14372 24392
rect 14366 24352 14372 24364
rect 14424 24352 14430 24404
rect 15838 24352 15844 24404
rect 15896 24392 15902 24404
rect 23014 24392 23020 24404
rect 15896 24364 23020 24392
rect 15896 24352 15902 24364
rect 23014 24352 23020 24364
rect 23072 24352 23078 24404
rect 23198 24392 23204 24404
rect 23159 24364 23204 24392
rect 23198 24352 23204 24364
rect 23256 24352 23262 24404
rect 23658 24392 23664 24404
rect 23619 24364 23664 24392
rect 23658 24352 23664 24364
rect 23716 24352 23722 24404
rect 29825 24395 29883 24401
rect 24504 24364 25176 24392
rect 14737 24327 14795 24333
rect 14737 24293 14749 24327
rect 14783 24324 14795 24327
rect 17310 24324 17316 24336
rect 14783 24296 17316 24324
rect 14783 24293 14795 24296
rect 14737 24287 14795 24293
rect 17310 24284 17316 24296
rect 17368 24284 17374 24336
rect 23382 24284 23388 24336
rect 23440 24324 23446 24336
rect 24504 24324 24532 24364
rect 23440 24296 24532 24324
rect 24581 24327 24639 24333
rect 23440 24284 23446 24296
rect 24581 24293 24593 24327
rect 24627 24293 24639 24327
rect 24581 24287 24639 24293
rect 15654 24256 15660 24268
rect 14568 24228 15660 24256
rect 14568 24197 14596 24228
rect 15654 24216 15660 24228
rect 15712 24216 15718 24268
rect 22094 24216 22100 24268
rect 22152 24256 22158 24268
rect 24486 24256 24492 24268
rect 22152 24228 24492 24256
rect 22152 24216 22158 24228
rect 24486 24216 24492 24228
rect 24544 24216 24550 24268
rect 14553 24191 14611 24197
rect 14553 24157 14565 24191
rect 14599 24157 14611 24191
rect 14553 24151 14611 24157
rect 14829 24191 14887 24197
rect 14829 24157 14841 24191
rect 14875 24157 14887 24191
rect 14829 24151 14887 24157
rect 17129 24191 17187 24197
rect 17129 24157 17141 24191
rect 17175 24188 17187 24191
rect 17494 24188 17500 24200
rect 17175 24160 17500 24188
rect 17175 24157 17187 24160
rect 17129 24151 17187 24157
rect 12802 24080 12808 24132
rect 12860 24120 12866 24132
rect 14844 24120 14872 24151
rect 17494 24148 17500 24160
rect 17552 24148 17558 24200
rect 18141 24191 18199 24197
rect 18141 24157 18153 24191
rect 18187 24188 18199 24191
rect 19242 24188 19248 24200
rect 18187 24160 19248 24188
rect 18187 24157 18199 24160
rect 18141 24151 18199 24157
rect 19242 24148 19248 24160
rect 19300 24148 19306 24200
rect 20622 24188 20628 24200
rect 20583 24160 20628 24188
rect 20622 24148 20628 24160
rect 20680 24148 20686 24200
rect 20892 24191 20950 24197
rect 20892 24157 20904 24191
rect 20938 24188 20950 24191
rect 22002 24188 22008 24200
rect 20938 24160 22008 24188
rect 20938 24157 20950 24160
rect 20892 24151 20950 24157
rect 22002 24148 22008 24160
rect 22060 24148 22066 24200
rect 23106 24188 23112 24200
rect 23019 24160 23112 24188
rect 23106 24148 23112 24160
rect 23164 24148 23170 24200
rect 23382 24188 23388 24200
rect 23343 24160 23388 24188
rect 23382 24148 23388 24160
rect 23440 24148 23446 24200
rect 24596 24188 24624 24287
rect 25148 24265 25176 24364
rect 29825 24361 29837 24395
rect 29871 24392 29883 24395
rect 30098 24392 30104 24404
rect 29871 24364 30104 24392
rect 29871 24361 29883 24364
rect 29825 24355 29883 24361
rect 30098 24352 30104 24364
rect 30156 24352 30162 24404
rect 42886 24392 42892 24404
rect 31726 24364 42892 24392
rect 25590 24284 25596 24336
rect 25648 24324 25654 24336
rect 25777 24327 25835 24333
rect 25777 24324 25789 24327
rect 25648 24296 25789 24324
rect 25648 24284 25654 24296
rect 25777 24293 25789 24296
rect 25823 24293 25835 24327
rect 31726 24324 31754 24364
rect 42886 24352 42892 24364
rect 42944 24352 42950 24404
rect 25777 24287 25835 24293
rect 28092 24296 31754 24324
rect 33689 24327 33747 24333
rect 25133 24259 25191 24265
rect 25133 24225 25145 24259
rect 25179 24225 25191 24259
rect 25133 24219 25191 24225
rect 26234 24216 26240 24268
rect 26292 24256 26298 24268
rect 27065 24259 27123 24265
rect 27065 24256 27077 24259
rect 26292 24228 27077 24256
rect 26292 24216 26298 24228
rect 27065 24225 27077 24228
rect 27111 24225 27123 24259
rect 27065 24219 27123 24225
rect 26053 24191 26111 24197
rect 26053 24188 26065 24191
rect 24596 24160 26065 24188
rect 26053 24157 26065 24160
rect 26099 24157 26111 24191
rect 26053 24151 26111 24157
rect 27154 24148 27160 24200
rect 27212 24188 27218 24200
rect 27321 24191 27379 24197
rect 27321 24188 27333 24191
rect 27212 24160 27333 24188
rect 27212 24148 27218 24160
rect 27321 24157 27333 24160
rect 27367 24157 27379 24191
rect 27321 24151 27379 24157
rect 17402 24120 17408 24132
rect 12860 24092 17408 24120
rect 12860 24080 12866 24092
rect 17402 24080 17408 24092
rect 17460 24080 17466 24132
rect 18506 24120 18512 24132
rect 18419 24092 18512 24120
rect 18506 24080 18512 24092
rect 18564 24120 18570 24132
rect 20254 24120 20260 24132
rect 18564 24092 20260 24120
rect 18564 24080 18570 24092
rect 20254 24080 20260 24092
rect 20312 24080 20318 24132
rect 23124 24120 23152 24148
rect 23474 24120 23480 24132
rect 23124 24092 23480 24120
rect 23474 24080 23480 24092
rect 23532 24120 23538 24132
rect 24762 24120 24768 24132
rect 23532 24092 24768 24120
rect 23532 24080 23538 24092
rect 24762 24080 24768 24092
rect 24820 24120 24826 24132
rect 25774 24120 25780 24132
rect 24820 24092 25084 24120
rect 25735 24092 25780 24120
rect 24820 24080 24826 24092
rect 16942 24052 16948 24064
rect 16903 24024 16948 24052
rect 16942 24012 16948 24024
rect 17000 24012 17006 24064
rect 21358 24012 21364 24064
rect 21416 24052 21422 24064
rect 22005 24055 22063 24061
rect 22005 24052 22017 24055
rect 21416 24024 22017 24052
rect 21416 24012 21422 24024
rect 22005 24021 22017 24024
rect 22051 24021 22063 24055
rect 22005 24015 22063 24021
rect 24394 24012 24400 24064
rect 24452 24052 24458 24064
rect 25056 24061 25084 24092
rect 25774 24080 25780 24092
rect 25832 24080 25838 24132
rect 25866 24080 25872 24132
rect 25924 24120 25930 24132
rect 25961 24123 26019 24129
rect 25961 24120 25973 24123
rect 25924 24092 25973 24120
rect 25924 24080 25930 24092
rect 25961 24089 25973 24092
rect 26007 24089 26019 24123
rect 25961 24083 26019 24089
rect 24949 24055 25007 24061
rect 24949 24052 24961 24055
rect 24452 24024 24961 24052
rect 24452 24012 24458 24024
rect 24949 24021 24961 24024
rect 24995 24021 25007 24055
rect 24949 24015 25007 24021
rect 25041 24055 25099 24061
rect 25041 24021 25053 24055
rect 25087 24052 25099 24055
rect 28092 24052 28120 24296
rect 33689 24293 33701 24327
rect 33735 24324 33747 24327
rect 34054 24324 34060 24336
rect 33735 24296 34060 24324
rect 33735 24293 33747 24296
rect 33689 24287 33747 24293
rect 34054 24284 34060 24296
rect 34112 24324 34118 24336
rect 39758 24324 39764 24336
rect 34112 24296 39764 24324
rect 34112 24284 34118 24296
rect 39758 24284 39764 24296
rect 39816 24284 39822 24336
rect 31570 24256 31576 24268
rect 30300 24228 31576 24256
rect 30300 24200 30328 24228
rect 31570 24216 31576 24228
rect 31628 24216 31634 24268
rect 35986 24216 35992 24268
rect 36044 24256 36050 24268
rect 36044 24228 36492 24256
rect 36044 24216 36050 24228
rect 30009 24191 30067 24197
rect 30009 24157 30021 24191
rect 30055 24157 30067 24191
rect 30282 24188 30288 24200
rect 30243 24160 30288 24188
rect 30009 24151 30067 24157
rect 30024 24120 30052 24151
rect 30282 24148 30288 24160
rect 30340 24148 30346 24200
rect 30469 24191 30527 24197
rect 30469 24157 30481 24191
rect 30515 24188 30527 24191
rect 32309 24191 32367 24197
rect 30515 24160 30871 24188
rect 30515 24157 30527 24160
rect 30469 24151 30527 24157
rect 30742 24120 30748 24132
rect 30024 24092 30748 24120
rect 30742 24080 30748 24092
rect 30800 24080 30806 24132
rect 25087 24024 28120 24052
rect 25087 24021 25099 24024
rect 25041 24015 25099 24021
rect 28166 24012 28172 24064
rect 28224 24052 28230 24064
rect 28445 24055 28503 24061
rect 28445 24052 28457 24055
rect 28224 24024 28457 24052
rect 28224 24012 28230 24024
rect 28445 24021 28457 24024
rect 28491 24021 28503 24055
rect 28445 24015 28503 24021
rect 29822 24012 29828 24064
rect 29880 24052 29886 24064
rect 30843 24052 30871 24160
rect 32309 24157 32321 24191
rect 32355 24188 32367 24191
rect 33778 24188 33784 24200
rect 32355 24160 33784 24188
rect 32355 24157 32367 24160
rect 32309 24151 32367 24157
rect 33778 24148 33784 24160
rect 33836 24148 33842 24200
rect 33870 24148 33876 24200
rect 33928 24188 33934 24200
rect 34054 24188 34060 24200
rect 33928 24160 34060 24188
rect 33928 24148 33934 24160
rect 34054 24148 34060 24160
rect 34112 24148 34118 24200
rect 36354 24188 36360 24200
rect 36315 24160 36360 24188
rect 36354 24148 36360 24160
rect 36412 24148 36418 24200
rect 36464 24197 36492 24228
rect 37274 24216 37280 24268
rect 37332 24256 37338 24268
rect 40037 24259 40095 24265
rect 40037 24256 40049 24259
rect 37332 24228 40049 24256
rect 37332 24216 37338 24228
rect 40037 24225 40049 24228
rect 40083 24225 40095 24259
rect 40037 24219 40095 24225
rect 36449 24191 36507 24197
rect 36449 24157 36461 24191
rect 36495 24157 36507 24191
rect 36449 24151 36507 24157
rect 39390 24148 39396 24200
rect 39448 24188 39454 24200
rect 39485 24191 39543 24197
rect 39485 24188 39497 24191
rect 39448 24160 39497 24188
rect 39448 24148 39454 24160
rect 39485 24157 39497 24160
rect 39531 24157 39543 24191
rect 39485 24151 39543 24157
rect 32582 24129 32588 24132
rect 32576 24083 32588 24129
rect 32640 24120 32646 24132
rect 40282 24123 40340 24129
rect 40282 24120 40294 24123
rect 32640 24092 32676 24120
rect 39316 24092 40294 24120
rect 32582 24080 32588 24083
rect 32640 24080 32646 24092
rect 29880 24024 30871 24052
rect 36357 24055 36415 24061
rect 29880 24012 29886 24024
rect 36357 24021 36369 24055
rect 36403 24052 36415 24055
rect 36446 24052 36452 24064
rect 36403 24024 36452 24052
rect 36403 24021 36415 24024
rect 36357 24015 36415 24021
rect 36446 24012 36452 24024
rect 36504 24012 36510 24064
rect 39316 24061 39344 24092
rect 40282 24089 40294 24092
rect 40328 24089 40340 24123
rect 40282 24083 40340 24089
rect 39301 24055 39359 24061
rect 39301 24021 39313 24055
rect 39347 24021 39359 24055
rect 39301 24015 39359 24021
rect 40862 24012 40868 24064
rect 40920 24052 40926 24064
rect 41417 24055 41475 24061
rect 41417 24052 41429 24055
rect 40920 24024 41429 24052
rect 40920 24012 40926 24024
rect 41417 24021 41429 24024
rect 41463 24021 41475 24055
rect 41417 24015 41475 24021
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 17494 23848 17500 23860
rect 17455 23820 17500 23848
rect 17494 23808 17500 23820
rect 17552 23808 17558 23860
rect 25038 23848 25044 23860
rect 24999 23820 25044 23848
rect 25038 23808 25044 23820
rect 25096 23808 25102 23860
rect 25682 23848 25688 23860
rect 25643 23820 25688 23848
rect 25682 23808 25688 23820
rect 25740 23808 25746 23860
rect 27522 23848 27528 23860
rect 27483 23820 27528 23848
rect 27522 23808 27528 23820
rect 27580 23808 27586 23860
rect 27632 23820 30052 23848
rect 11882 23780 11888 23792
rect 11843 23752 11888 23780
rect 11882 23740 11888 23752
rect 11940 23740 11946 23792
rect 16850 23740 16856 23792
rect 16908 23780 16914 23792
rect 17037 23783 17095 23789
rect 17037 23780 17049 23783
rect 16908 23752 17049 23780
rect 16908 23740 16914 23752
rect 17037 23749 17049 23752
rect 17083 23780 17095 23783
rect 18506 23780 18512 23792
rect 17083 23752 18512 23780
rect 17083 23749 17095 23752
rect 17037 23743 17095 23749
rect 18506 23740 18512 23752
rect 18564 23740 18570 23792
rect 18785 23783 18843 23789
rect 18785 23749 18797 23783
rect 18831 23780 18843 23783
rect 19426 23780 19432 23792
rect 18831 23752 19432 23780
rect 18831 23749 18843 23752
rect 18785 23743 18843 23749
rect 19426 23740 19432 23752
rect 19484 23740 19490 23792
rect 19797 23783 19855 23789
rect 19797 23749 19809 23783
rect 19843 23780 19855 23783
rect 20162 23780 20168 23792
rect 19843 23752 20168 23780
rect 19843 23749 19855 23752
rect 19797 23743 19855 23749
rect 20162 23740 20168 23752
rect 20220 23740 20226 23792
rect 24394 23740 24400 23792
rect 24452 23780 24458 23792
rect 24673 23783 24731 23789
rect 24673 23780 24685 23783
rect 24452 23752 24685 23780
rect 24452 23740 24458 23752
rect 24673 23749 24685 23752
rect 24719 23749 24731 23783
rect 24673 23743 24731 23749
rect 24857 23783 24915 23789
rect 24857 23749 24869 23783
rect 24903 23780 24915 23783
rect 27632 23780 27660 23820
rect 29914 23780 29920 23792
rect 24903 23752 27660 23780
rect 27724 23752 29920 23780
rect 24903 23749 24915 23752
rect 24857 23743 24915 23749
rect 17954 23712 17960 23724
rect 17915 23684 17960 23712
rect 17954 23672 17960 23684
rect 18012 23672 18018 23724
rect 18874 23672 18880 23724
rect 18932 23712 18938 23724
rect 19981 23715 20039 23721
rect 19981 23712 19993 23715
rect 18932 23684 19993 23712
rect 18932 23672 18938 23684
rect 19981 23681 19993 23684
rect 20027 23681 20039 23715
rect 19981 23675 20039 23681
rect 21910 23672 21916 23724
rect 21968 23712 21974 23724
rect 22465 23715 22523 23721
rect 22465 23712 22477 23715
rect 21968 23684 22477 23712
rect 21968 23672 21974 23684
rect 22465 23681 22477 23684
rect 22511 23681 22523 23715
rect 22465 23675 22523 23681
rect 24121 23715 24179 23721
rect 24121 23681 24133 23715
rect 24167 23712 24179 23715
rect 24210 23712 24216 23724
rect 24167 23684 24216 23712
rect 24167 23681 24179 23684
rect 24121 23675 24179 23681
rect 24210 23672 24216 23684
rect 24268 23712 24274 23724
rect 24872 23712 24900 23743
rect 25590 23712 25596 23724
rect 24268 23684 24900 23712
rect 25551 23684 25596 23712
rect 24268 23672 24274 23684
rect 25590 23672 25596 23684
rect 25648 23672 25654 23724
rect 25774 23712 25780 23724
rect 25735 23684 25780 23712
rect 25774 23672 25780 23684
rect 25832 23672 25838 23724
rect 27724 23721 27752 23752
rect 29914 23740 29920 23752
rect 29972 23740 29978 23792
rect 30024 23780 30052 23820
rect 30742 23808 30748 23860
rect 30800 23848 30806 23860
rect 32398 23848 32404 23860
rect 30800 23820 32404 23848
rect 30800 23808 30806 23820
rect 32398 23808 32404 23820
rect 32456 23808 32462 23860
rect 32582 23848 32588 23860
rect 32543 23820 32588 23848
rect 32582 23808 32588 23820
rect 32640 23808 32646 23860
rect 39390 23848 39396 23860
rect 39351 23820 39396 23848
rect 39390 23808 39396 23820
rect 39448 23808 39454 23860
rect 39758 23848 39764 23860
rect 39719 23820 39764 23848
rect 39758 23808 39764 23820
rect 39816 23808 39822 23860
rect 39853 23851 39911 23857
rect 39853 23817 39865 23851
rect 39899 23848 39911 23851
rect 41141 23851 41199 23857
rect 41141 23848 41153 23851
rect 39899 23820 41153 23848
rect 39899 23817 39911 23820
rect 39853 23811 39911 23817
rect 41141 23817 41153 23820
rect 41187 23817 41199 23851
rect 41141 23811 41199 23817
rect 46934 23780 46940 23792
rect 30024 23752 46940 23780
rect 46934 23740 46940 23752
rect 46992 23740 46998 23792
rect 27709 23715 27767 23721
rect 27709 23712 27721 23715
rect 26528 23684 27721 23712
rect 26528 23644 26556 23684
rect 27709 23681 27721 23684
rect 27755 23681 27767 23715
rect 27709 23675 27767 23681
rect 27985 23715 28043 23721
rect 27985 23681 27997 23715
rect 28031 23681 28043 23715
rect 28166 23712 28172 23724
rect 28127 23684 28172 23712
rect 27985 23675 28043 23681
rect 22664 23616 26556 23644
rect 17405 23579 17463 23585
rect 17405 23545 17417 23579
rect 17451 23576 17463 23579
rect 18046 23576 18052 23588
rect 17451 23548 18052 23576
rect 17451 23545 17463 23548
rect 17405 23539 17463 23545
rect 18046 23536 18052 23548
rect 18104 23536 18110 23588
rect 4062 23468 4068 23520
rect 4120 23508 4126 23520
rect 11054 23508 11060 23520
rect 4120 23480 11060 23508
rect 4120 23468 4126 23480
rect 11054 23468 11060 23480
rect 11112 23468 11118 23520
rect 12161 23511 12219 23517
rect 12161 23477 12173 23511
rect 12207 23508 12219 23511
rect 13354 23508 13360 23520
rect 12207 23480 13360 23508
rect 12207 23477 12219 23480
rect 12161 23471 12219 23477
rect 13354 23468 13360 23480
rect 13412 23468 13418 23520
rect 20165 23511 20223 23517
rect 20165 23477 20177 23511
rect 20211 23508 20223 23511
rect 21450 23508 21456 23520
rect 20211 23480 21456 23508
rect 20211 23477 20223 23480
rect 20165 23471 20223 23477
rect 21450 23468 21456 23480
rect 21508 23468 21514 23520
rect 22278 23468 22284 23520
rect 22336 23508 22342 23520
rect 22664 23517 22692 23616
rect 26694 23604 26700 23656
rect 26752 23644 26758 23656
rect 28000 23644 28028 23675
rect 28166 23672 28172 23684
rect 28224 23672 28230 23724
rect 29546 23712 29552 23724
rect 29507 23684 29552 23712
rect 29546 23672 29552 23684
rect 29604 23672 29610 23724
rect 29638 23672 29644 23724
rect 29696 23712 29702 23724
rect 29733 23715 29791 23721
rect 29733 23712 29745 23715
rect 29696 23684 29745 23712
rect 29696 23672 29702 23684
rect 29733 23681 29745 23684
rect 29779 23681 29791 23715
rect 32766 23712 32772 23724
rect 32727 23684 32772 23712
rect 29733 23675 29791 23681
rect 32766 23672 32772 23684
rect 32824 23672 32830 23724
rect 33778 23712 33784 23724
rect 33739 23684 33784 23712
rect 33778 23672 33784 23684
rect 33836 23672 33842 23724
rect 33870 23672 33876 23724
rect 33928 23712 33934 23724
rect 34037 23715 34095 23721
rect 34037 23712 34049 23715
rect 33928 23684 34049 23712
rect 33928 23672 33934 23684
rect 34037 23681 34049 23684
rect 34083 23681 34095 23715
rect 36446 23712 36452 23724
rect 36407 23684 36452 23712
rect 34037 23675 34095 23681
rect 36446 23672 36452 23684
rect 36504 23672 36510 23724
rect 36633 23715 36691 23721
rect 36633 23681 36645 23715
rect 36679 23712 36691 23715
rect 37366 23712 37372 23724
rect 36679 23684 37372 23712
rect 36679 23681 36691 23684
rect 36633 23675 36691 23681
rect 37366 23672 37372 23684
rect 37424 23672 37430 23724
rect 40773 23715 40831 23721
rect 40773 23681 40785 23715
rect 40819 23712 40831 23715
rect 40862 23712 40868 23724
rect 40819 23684 40868 23712
rect 40819 23681 40831 23684
rect 40773 23675 40831 23681
rect 40862 23672 40868 23684
rect 40920 23672 40926 23724
rect 46290 23712 46296 23724
rect 46251 23684 46296 23712
rect 46290 23672 46296 23684
rect 46348 23672 46354 23724
rect 29822 23644 29828 23656
rect 26752 23616 28028 23644
rect 29783 23616 29828 23644
rect 26752 23604 26758 23616
rect 23014 23536 23020 23588
rect 23072 23576 23078 23588
rect 27890 23576 27896 23588
rect 23072 23548 27896 23576
rect 23072 23536 23078 23548
rect 27890 23536 27896 23548
rect 27948 23536 27954 23588
rect 28000 23576 28028 23616
rect 29822 23604 29828 23616
rect 29880 23604 29886 23656
rect 31846 23604 31852 23656
rect 31904 23644 31910 23656
rect 33045 23647 33103 23653
rect 33045 23644 33057 23647
rect 31904 23616 33057 23644
rect 31904 23604 31910 23616
rect 33045 23613 33057 23616
rect 33091 23613 33103 23647
rect 33045 23607 33103 23613
rect 39942 23604 39948 23656
rect 40000 23644 40006 23656
rect 40678 23644 40684 23656
rect 40000 23616 40045 23644
rect 40639 23616 40684 23644
rect 40000 23604 40006 23616
rect 40678 23604 40684 23616
rect 40736 23604 40742 23656
rect 30098 23576 30104 23588
rect 28000 23548 30104 23576
rect 30098 23536 30104 23548
rect 30156 23536 30162 23588
rect 31662 23536 31668 23588
rect 31720 23576 31726 23588
rect 32953 23579 33011 23585
rect 32953 23576 32965 23579
rect 31720 23548 32965 23576
rect 31720 23536 31726 23548
rect 32953 23545 32965 23548
rect 32999 23576 33011 23579
rect 33134 23576 33140 23588
rect 32999 23548 33140 23576
rect 32999 23545 33011 23548
rect 32953 23539 33011 23545
rect 33134 23536 33140 23548
rect 33192 23536 33198 23588
rect 22649 23511 22707 23517
rect 22649 23508 22661 23511
rect 22336 23480 22661 23508
rect 22336 23468 22342 23480
rect 22649 23477 22661 23480
rect 22695 23477 22707 23511
rect 22649 23471 22707 23477
rect 23382 23468 23388 23520
rect 23440 23508 23446 23520
rect 23937 23511 23995 23517
rect 23937 23508 23949 23511
rect 23440 23480 23949 23508
rect 23440 23468 23446 23480
rect 23937 23477 23949 23480
rect 23983 23477 23995 23511
rect 23937 23471 23995 23477
rect 24762 23468 24768 23520
rect 24820 23508 24826 23520
rect 24857 23511 24915 23517
rect 24857 23508 24869 23511
rect 24820 23480 24869 23508
rect 24820 23468 24826 23480
rect 24857 23477 24869 23480
rect 24903 23477 24915 23511
rect 24857 23471 24915 23477
rect 25774 23468 25780 23520
rect 25832 23508 25838 23520
rect 28258 23508 28264 23520
rect 25832 23480 28264 23508
rect 25832 23468 25838 23480
rect 28258 23468 28264 23480
rect 28316 23468 28322 23520
rect 29365 23511 29423 23517
rect 29365 23477 29377 23511
rect 29411 23508 29423 23511
rect 29454 23508 29460 23520
rect 29411 23480 29460 23508
rect 29411 23477 29423 23480
rect 29365 23471 29423 23477
rect 29454 23468 29460 23480
rect 29512 23468 29518 23520
rect 31478 23468 31484 23520
rect 31536 23508 31542 23520
rect 34054 23508 34060 23520
rect 31536 23480 34060 23508
rect 31536 23468 31542 23480
rect 34054 23468 34060 23480
rect 34112 23468 34118 23520
rect 35161 23511 35219 23517
rect 35161 23477 35173 23511
rect 35207 23508 35219 23511
rect 35342 23508 35348 23520
rect 35207 23480 35348 23508
rect 35207 23477 35219 23480
rect 35161 23471 35219 23477
rect 35342 23468 35348 23480
rect 35400 23468 35406 23520
rect 36538 23508 36544 23520
rect 36499 23480 36544 23508
rect 36538 23468 36544 23480
rect 36596 23468 36602 23520
rect 46382 23508 46388 23520
rect 46343 23480 46388 23508
rect 46382 23468 46388 23480
rect 46440 23468 46446 23520
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 12986 23264 12992 23316
rect 13044 23304 13050 23316
rect 17681 23307 17739 23313
rect 17681 23304 17693 23307
rect 13044 23276 17693 23304
rect 13044 23264 13050 23276
rect 17681 23273 17693 23276
rect 17727 23273 17739 23307
rect 18046 23304 18052 23316
rect 18007 23276 18052 23304
rect 17681 23267 17739 23273
rect 11054 23168 11060 23180
rect 11015 23140 11060 23168
rect 11054 23128 11060 23140
rect 11112 23128 11118 23180
rect 13906 23128 13912 23180
rect 13964 23168 13970 23180
rect 14277 23171 14335 23177
rect 14277 23168 14289 23171
rect 13964 23140 14289 23168
rect 13964 23128 13970 23140
rect 14277 23137 14289 23140
rect 14323 23137 14335 23171
rect 17696 23168 17724 23267
rect 18046 23264 18052 23276
rect 18104 23264 18110 23316
rect 22741 23307 22799 23313
rect 22741 23273 22753 23307
rect 22787 23304 22799 23307
rect 23474 23304 23480 23316
rect 22787 23276 23480 23304
rect 22787 23273 22799 23276
rect 22741 23267 22799 23273
rect 23474 23264 23480 23276
rect 23532 23264 23538 23316
rect 24578 23264 24584 23316
rect 24636 23304 24642 23316
rect 24857 23307 24915 23313
rect 24857 23304 24869 23307
rect 24636 23276 24869 23304
rect 24636 23264 24642 23276
rect 24857 23273 24869 23276
rect 24903 23273 24915 23307
rect 24857 23267 24915 23273
rect 29546 23264 29552 23316
rect 29604 23304 29610 23316
rect 29733 23307 29791 23313
rect 29733 23304 29745 23307
rect 29604 23276 29745 23304
rect 29604 23264 29610 23276
rect 29733 23273 29745 23276
rect 29779 23273 29791 23307
rect 29733 23267 29791 23273
rect 40313 23307 40371 23313
rect 40313 23273 40325 23307
rect 40359 23304 40371 23307
rect 40678 23304 40684 23316
rect 40359 23276 40684 23304
rect 40359 23273 40371 23276
rect 40313 23267 40371 23273
rect 40678 23264 40684 23276
rect 40736 23264 40742 23316
rect 27617 23239 27675 23245
rect 27617 23205 27629 23239
rect 27663 23205 27675 23239
rect 27617 23199 27675 23205
rect 17696 23140 18276 23168
rect 14277 23131 14335 23137
rect 10134 23100 10140 23112
rect 10095 23072 10140 23100
rect 10134 23060 10140 23072
rect 10192 23060 10198 23112
rect 14550 23100 14556 23112
rect 14511 23072 14556 23100
rect 14550 23060 14556 23072
rect 14608 23060 14614 23112
rect 16025 23103 16083 23109
rect 16025 23069 16037 23103
rect 16071 23100 16083 23103
rect 18138 23100 18144 23112
rect 16071 23072 18144 23100
rect 16071 23069 16083 23072
rect 16025 23063 16083 23069
rect 18138 23060 18144 23072
rect 18196 23060 18202 23112
rect 18248 23100 18276 23140
rect 18414 23128 18420 23180
rect 18472 23168 18478 23180
rect 18601 23171 18659 23177
rect 18601 23168 18613 23171
rect 18472 23140 18613 23168
rect 18472 23128 18478 23140
rect 18601 23137 18613 23140
rect 18647 23137 18659 23171
rect 19426 23168 19432 23180
rect 19387 23140 19432 23168
rect 18601 23131 18659 23137
rect 19426 23128 19432 23140
rect 19484 23128 19490 23180
rect 27632 23168 27660 23199
rect 39209 23171 39267 23177
rect 20456 23140 31754 23168
rect 18506 23100 18512 23112
rect 18248 23072 18512 23100
rect 18506 23060 18512 23072
rect 18564 23060 18570 23112
rect 18874 23060 18880 23112
rect 18932 23100 18938 23112
rect 20456 23100 20484 23140
rect 21450 23100 21456 23112
rect 18932 23072 20484 23100
rect 21411 23072 21456 23100
rect 18932 23060 18938 23072
rect 21450 23060 21456 23072
rect 21508 23060 21514 23112
rect 24670 23100 24676 23112
rect 24631 23072 24676 23100
rect 24670 23060 24676 23072
rect 24728 23060 24734 23112
rect 26234 23060 26240 23112
rect 26292 23100 26298 23112
rect 27433 23103 27491 23109
rect 27433 23100 27445 23103
rect 26292 23072 27445 23100
rect 26292 23060 26298 23072
rect 27433 23069 27445 23072
rect 27479 23100 27491 23103
rect 27706 23100 27712 23112
rect 27479 23072 27712 23100
rect 27479 23069 27491 23072
rect 27433 23063 27491 23069
rect 27706 23060 27712 23072
rect 27764 23060 27770 23112
rect 29914 23100 29920 23112
rect 29875 23072 29920 23100
rect 29914 23060 29920 23072
rect 29972 23060 29978 23112
rect 30098 23060 30104 23112
rect 30156 23100 30162 23112
rect 30193 23103 30251 23109
rect 30193 23100 30205 23103
rect 30156 23072 30205 23100
rect 30156 23060 30162 23072
rect 30193 23069 30205 23072
rect 30239 23069 30251 23103
rect 30193 23063 30251 23069
rect 30377 23103 30435 23109
rect 30377 23069 30389 23103
rect 30423 23100 30435 23103
rect 30558 23100 30564 23112
rect 30423 23072 30564 23100
rect 30423 23069 30435 23072
rect 30377 23063 30435 23069
rect 10321 23035 10379 23041
rect 10321 23001 10333 23035
rect 10367 23032 10379 23035
rect 10502 23032 10508 23044
rect 10367 23004 10508 23032
rect 10367 23001 10379 23004
rect 10321 22995 10379 23001
rect 10502 22992 10508 23004
rect 10560 22992 10566 23044
rect 16292 23035 16350 23041
rect 16292 23001 16304 23035
rect 16338 23032 16350 23035
rect 16942 23032 16948 23044
rect 16338 23004 16948 23032
rect 16338 23001 16350 23004
rect 16292 22995 16350 23001
rect 16942 22992 16948 23004
rect 17000 22992 17006 23044
rect 18417 23035 18475 23041
rect 18417 23032 18429 23035
rect 17420 23004 18429 23032
rect 17310 22924 17316 22976
rect 17368 22964 17374 22976
rect 17420 22973 17448 23004
rect 18417 23001 18429 23004
rect 18463 23001 18475 23035
rect 18417 22995 18475 23001
rect 19696 23035 19754 23041
rect 19696 23001 19708 23035
rect 19742 23032 19754 23035
rect 22557 23035 22615 23041
rect 19742 23004 21312 23032
rect 19742 23001 19754 23004
rect 19696 22995 19754 23001
rect 17405 22967 17463 22973
rect 17405 22964 17417 22967
rect 17368 22936 17417 22964
rect 17368 22924 17374 22936
rect 17405 22933 17417 22936
rect 17451 22933 17463 22967
rect 17405 22927 17463 22933
rect 20530 22924 20536 22976
rect 20588 22964 20594 22976
rect 21284 22973 21312 23004
rect 22557 23001 22569 23035
rect 22603 23032 22615 23035
rect 22646 23032 22652 23044
rect 22603 23004 22652 23032
rect 22603 23001 22615 23004
rect 22557 22995 22615 23001
rect 22646 22992 22652 23004
rect 22704 22992 22710 23044
rect 22773 23035 22831 23041
rect 22773 23001 22785 23035
rect 22819 23032 22831 23035
rect 23382 23032 23388 23044
rect 22819 23004 23388 23032
rect 22819 23001 22831 23004
rect 22773 22995 22831 23001
rect 23382 22992 23388 23004
rect 23440 22992 23446 23044
rect 30208 23032 30236 23063
rect 30558 23060 30564 23072
rect 30616 23060 30622 23112
rect 31726 23100 31754 23140
rect 39209 23137 39221 23171
rect 39255 23168 39267 23171
rect 40034 23168 40040 23180
rect 39255 23140 40040 23168
rect 39255 23137 39267 23140
rect 39209 23131 39267 23137
rect 40034 23128 40040 23140
rect 40092 23128 40098 23180
rect 47578 23168 47584 23180
rect 47539 23140 47584 23168
rect 47578 23128 47584 23140
rect 47636 23128 47642 23180
rect 33873 23103 33931 23109
rect 33873 23100 33885 23103
rect 31726 23072 33885 23100
rect 33873 23069 33885 23072
rect 33919 23100 33931 23103
rect 33962 23100 33968 23112
rect 33919 23072 33968 23100
rect 33919 23069 33931 23072
rect 33873 23063 33931 23069
rect 33962 23060 33968 23072
rect 34020 23060 34026 23112
rect 34054 23060 34060 23112
rect 34112 23100 34118 23112
rect 34149 23103 34207 23109
rect 34149 23100 34161 23103
rect 34112 23072 34161 23100
rect 34112 23060 34118 23072
rect 34149 23069 34161 23072
rect 34195 23069 34207 23103
rect 34149 23063 34207 23069
rect 34333 23103 34391 23109
rect 34333 23069 34345 23103
rect 34379 23100 34391 23103
rect 35342 23100 35348 23112
rect 34379 23072 35348 23100
rect 34379 23069 34391 23072
rect 34333 23063 34391 23069
rect 35342 23060 35348 23072
rect 35400 23060 35406 23112
rect 36262 23060 36268 23112
rect 36320 23100 36326 23112
rect 36357 23103 36415 23109
rect 36357 23100 36369 23103
rect 36320 23072 36369 23100
rect 36320 23060 36326 23072
rect 36357 23069 36369 23072
rect 36403 23069 36415 23103
rect 36538 23100 36544 23112
rect 36499 23072 36544 23100
rect 36357 23063 36415 23069
rect 36538 23060 36544 23072
rect 36596 23060 36602 23112
rect 36633 23103 36691 23109
rect 36633 23069 36645 23103
rect 36679 23100 36691 23103
rect 37461 23103 37519 23109
rect 37461 23100 37473 23103
rect 36679 23072 37473 23100
rect 36679 23069 36691 23072
rect 36633 23063 36691 23069
rect 37461 23069 37473 23072
rect 37507 23069 37519 23103
rect 39114 23100 39120 23112
rect 39075 23072 39120 23100
rect 37461 23063 37519 23069
rect 39114 23060 39120 23072
rect 39172 23060 39178 23112
rect 39301 23103 39359 23109
rect 39301 23069 39313 23103
rect 39347 23069 39359 23103
rect 39301 23063 39359 23069
rect 31478 23032 31484 23044
rect 30208 23004 31484 23032
rect 31478 22992 31484 23004
rect 31536 22992 31542 23044
rect 36446 22992 36452 23044
rect 36504 23032 36510 23044
rect 37093 23035 37151 23041
rect 37093 23032 37105 23035
rect 36504 23004 37105 23032
rect 36504 22992 36510 23004
rect 37093 23001 37105 23004
rect 37139 23001 37151 23035
rect 37093 22995 37151 23001
rect 37277 23035 37335 23041
rect 37277 23001 37289 23035
rect 37323 23001 37335 23035
rect 39316 23032 39344 23063
rect 39390 23060 39396 23112
rect 39448 23100 39454 23112
rect 40221 23103 40279 23109
rect 39448 23072 39493 23100
rect 39448 23060 39454 23072
rect 40221 23069 40233 23103
rect 40267 23100 40279 23103
rect 40310 23100 40316 23112
rect 40267 23072 40316 23100
rect 40267 23069 40279 23072
rect 40221 23063 40279 23069
rect 40310 23060 40316 23072
rect 40368 23060 40374 23112
rect 40405 23103 40463 23109
rect 40405 23069 40417 23103
rect 40451 23100 40463 23103
rect 40586 23100 40592 23112
rect 40451 23072 40592 23100
rect 40451 23069 40463 23072
rect 40405 23063 40463 23069
rect 39574 23032 39580 23044
rect 39316 23004 39580 23032
rect 37277 22995 37335 23001
rect 20809 22967 20867 22973
rect 20809 22964 20821 22967
rect 20588 22936 20821 22964
rect 20588 22924 20594 22936
rect 20809 22933 20821 22936
rect 20855 22933 20867 22967
rect 20809 22927 20867 22933
rect 21269 22967 21327 22973
rect 21269 22933 21281 22967
rect 21315 22933 21327 22967
rect 22922 22964 22928 22976
rect 22883 22936 22928 22964
rect 21269 22927 21327 22933
rect 22922 22924 22928 22936
rect 22980 22924 22986 22976
rect 27706 22924 27712 22976
rect 27764 22964 27770 22976
rect 31846 22964 31852 22976
rect 27764 22936 31852 22964
rect 27764 22924 27770 22936
rect 31846 22924 31852 22936
rect 31904 22924 31910 22976
rect 33686 22964 33692 22976
rect 33647 22936 33692 22964
rect 33686 22924 33692 22936
rect 33744 22924 33750 22976
rect 35802 22924 35808 22976
rect 35860 22964 35866 22976
rect 36173 22967 36231 22973
rect 36173 22964 36185 22967
rect 35860 22936 36185 22964
rect 35860 22924 35866 22936
rect 36173 22933 36185 22936
rect 36219 22933 36231 22967
rect 37292 22964 37320 22995
rect 39574 22992 39580 23004
rect 39632 23032 39638 23044
rect 40420 23032 40448 23063
rect 40586 23060 40592 23072
rect 40644 23060 40650 23112
rect 45922 23100 45928 23112
rect 45883 23072 45928 23100
rect 45922 23060 45928 23072
rect 45980 23060 45986 23112
rect 46106 23032 46112 23044
rect 39632 23004 40448 23032
rect 46067 23004 46112 23032
rect 39632 22992 39638 23004
rect 46106 22992 46112 23004
rect 46164 22992 46170 23044
rect 37366 22964 37372 22976
rect 37279 22936 37372 22964
rect 36173 22927 36231 22933
rect 37366 22924 37372 22936
rect 37424 22964 37430 22976
rect 38933 22967 38991 22973
rect 38933 22964 38945 22967
rect 37424 22936 38945 22964
rect 37424 22924 37430 22936
rect 38933 22933 38945 22936
rect 38979 22933 38991 22967
rect 38933 22927 38991 22933
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 10502 22760 10508 22772
rect 10463 22732 10508 22760
rect 10502 22720 10508 22732
rect 10560 22720 10566 22772
rect 18233 22763 18291 22769
rect 18233 22729 18245 22763
rect 18279 22760 18291 22763
rect 18966 22760 18972 22772
rect 18279 22732 18972 22760
rect 18279 22729 18291 22732
rect 18233 22723 18291 22729
rect 18966 22720 18972 22732
rect 19024 22720 19030 22772
rect 20162 22760 20168 22772
rect 20123 22732 20168 22760
rect 20162 22720 20168 22732
rect 20220 22720 20226 22772
rect 20530 22760 20536 22772
rect 20491 22732 20536 22760
rect 20530 22720 20536 22732
rect 20588 22720 20594 22772
rect 20625 22763 20683 22769
rect 20625 22729 20637 22763
rect 20671 22760 20683 22763
rect 27706 22760 27712 22772
rect 20671 22732 27712 22760
rect 20671 22729 20683 22732
rect 20625 22723 20683 22729
rect 27706 22720 27712 22732
rect 27764 22720 27770 22772
rect 31754 22760 31760 22772
rect 27816 22732 31760 22760
rect 14550 22692 14556 22704
rect 12268 22664 14556 22692
rect 10410 22624 10416 22636
rect 10371 22596 10416 22624
rect 10410 22584 10416 22596
rect 10468 22584 10474 22636
rect 12158 22516 12164 22568
rect 12216 22556 12222 22568
rect 12268 22565 12296 22664
rect 12526 22633 12532 22636
rect 12520 22587 12532 22633
rect 12584 22624 12590 22636
rect 14200 22633 14228 22664
rect 14550 22652 14556 22664
rect 14608 22652 14614 22704
rect 16850 22692 16856 22704
rect 16811 22664 16856 22692
rect 16850 22652 16856 22664
rect 16908 22652 16914 22704
rect 14185 22627 14243 22633
rect 12584 22596 12620 22624
rect 12526 22584 12532 22587
rect 12584 22584 12590 22596
rect 14185 22593 14197 22627
rect 14231 22593 14243 22627
rect 14185 22587 14243 22593
rect 14274 22584 14280 22636
rect 14332 22624 14338 22636
rect 14441 22627 14499 22633
rect 14441 22624 14453 22627
rect 14332 22596 14453 22624
rect 14332 22584 14338 22596
rect 14441 22593 14453 22596
rect 14487 22593 14499 22627
rect 14441 22587 14499 22593
rect 18141 22627 18199 22633
rect 18141 22593 18153 22627
rect 18187 22624 18199 22627
rect 18782 22624 18788 22636
rect 18187 22596 18788 22624
rect 18187 22593 18199 22596
rect 18141 22587 18199 22593
rect 18782 22584 18788 22596
rect 18840 22584 18846 22636
rect 18984 22624 19012 22720
rect 22189 22695 22247 22701
rect 22189 22661 22201 22695
rect 22235 22692 22247 22695
rect 22922 22692 22928 22704
rect 22235 22664 22928 22692
rect 22235 22661 22247 22664
rect 22189 22655 22247 22661
rect 22922 22652 22928 22664
rect 22980 22652 22986 22704
rect 27816 22692 27844 22732
rect 31754 22720 31760 22732
rect 31812 22720 31818 22772
rect 33597 22763 33655 22769
rect 33597 22729 33609 22763
rect 33643 22760 33655 22763
rect 33870 22760 33876 22772
rect 33643 22732 33876 22760
rect 33643 22729 33655 22732
rect 33597 22723 33655 22729
rect 33870 22720 33876 22732
rect 33928 22720 33934 22772
rect 38746 22760 38752 22772
rect 34072 22732 38752 22760
rect 29362 22692 29368 22704
rect 23400 22664 27844 22692
rect 29196 22664 29368 22692
rect 23400 22624 23428 22664
rect 18984 22596 23428 22624
rect 23474 22584 23480 22636
rect 23532 22624 23538 22636
rect 24489 22627 24547 22633
rect 24489 22624 24501 22627
rect 23532 22596 23577 22624
rect 23768 22596 24501 22624
rect 23532 22584 23538 22596
rect 12253 22559 12311 22565
rect 12253 22556 12265 22559
rect 12216 22528 12265 22556
rect 12216 22516 12222 22528
rect 12253 22525 12265 22528
rect 12299 22525 12311 22559
rect 18414 22556 18420 22568
rect 18375 22528 18420 22556
rect 12253 22519 12311 22525
rect 18414 22516 18420 22528
rect 18472 22556 18478 22568
rect 19334 22556 19340 22568
rect 18472 22528 19340 22556
rect 18472 22516 18478 22528
rect 19334 22516 19340 22528
rect 19392 22556 19398 22568
rect 20717 22559 20775 22565
rect 20717 22556 20729 22559
rect 19392 22528 20729 22556
rect 19392 22516 19398 22528
rect 20717 22525 20729 22528
rect 20763 22556 20775 22559
rect 21726 22556 21732 22568
rect 20763 22528 21732 22556
rect 20763 22525 20775 22528
rect 20717 22519 20775 22525
rect 21726 22516 21732 22528
rect 21784 22516 21790 22568
rect 22646 22516 22652 22568
rect 22704 22556 22710 22568
rect 23198 22556 23204 22568
rect 22704 22528 23204 22556
rect 22704 22516 22710 22528
rect 23198 22516 23204 22528
rect 23256 22556 23262 22568
rect 23768 22565 23796 22596
rect 24489 22593 24501 22596
rect 24535 22593 24547 22627
rect 24489 22587 24547 22593
rect 28994 22584 29000 22636
rect 29052 22624 29058 22636
rect 29196 22633 29224 22664
rect 29362 22652 29368 22664
rect 29420 22652 29426 22704
rect 30834 22652 30840 22704
rect 30892 22692 30898 22704
rect 32493 22695 32551 22701
rect 32493 22692 32505 22695
rect 30892 22664 32505 22692
rect 30892 22652 30898 22664
rect 29454 22633 29460 22636
rect 29181 22627 29239 22633
rect 29181 22624 29193 22627
rect 29052 22596 29193 22624
rect 29052 22584 29058 22596
rect 29181 22593 29193 22596
rect 29227 22593 29239 22627
rect 29448 22624 29460 22633
rect 29415 22596 29460 22624
rect 29181 22587 29239 22593
rect 29448 22587 29460 22596
rect 29454 22584 29460 22587
rect 29512 22584 29518 22636
rect 31772 22633 31800 22664
rect 32493 22661 32505 22664
rect 32539 22661 32551 22695
rect 32493 22655 32551 22661
rect 33502 22652 33508 22704
rect 33560 22692 33566 22704
rect 34072 22692 34100 22732
rect 38746 22720 38752 22732
rect 38804 22760 38810 22772
rect 39666 22760 39672 22772
rect 38804 22732 39672 22760
rect 38804 22720 38810 22732
rect 39666 22720 39672 22732
rect 39724 22720 39730 22772
rect 40034 22720 40040 22772
rect 40092 22760 40098 22772
rect 40497 22763 40555 22769
rect 40497 22760 40509 22763
rect 40092 22732 40509 22760
rect 40092 22720 40098 22732
rect 40497 22729 40509 22732
rect 40543 22760 40555 22763
rect 40862 22760 40868 22772
rect 40543 22732 40868 22760
rect 40543 22729 40555 22732
rect 40497 22723 40555 22729
rect 40862 22720 40868 22732
rect 40920 22720 40926 22772
rect 46106 22760 46112 22772
rect 46067 22732 46112 22760
rect 46106 22720 46112 22732
rect 46164 22720 46170 22772
rect 33560 22664 34100 22692
rect 33560 22652 33566 22664
rect 31573 22627 31631 22633
rect 31573 22593 31585 22627
rect 31619 22593 31631 22627
rect 31573 22587 31631 22593
rect 31757 22627 31815 22633
rect 31757 22593 31769 22627
rect 31803 22624 31815 22627
rect 32309 22627 32367 22633
rect 31803 22596 31837 22624
rect 31803 22593 31815 22596
rect 31757 22587 31815 22593
rect 32309 22593 32321 22627
rect 32355 22593 32367 22627
rect 32309 22587 32367 22593
rect 23753 22559 23811 22565
rect 23753 22556 23765 22559
rect 23256 22528 23765 22556
rect 23256 22516 23262 22528
rect 23753 22525 23765 22528
rect 23799 22525 23811 22559
rect 31588 22556 31616 22587
rect 31846 22556 31852 22568
rect 31588 22528 31852 22556
rect 23753 22519 23811 22525
rect 31846 22516 31852 22528
rect 31904 22556 31910 22568
rect 32324 22556 32352 22587
rect 33686 22584 33692 22636
rect 33744 22624 33750 22636
rect 34072 22633 34100 22664
rect 35342 22652 35348 22704
rect 35400 22692 35406 22704
rect 38841 22695 38899 22701
rect 35400 22664 36400 22692
rect 35400 22652 35406 22664
rect 33781 22627 33839 22633
rect 33781 22624 33793 22627
rect 33744 22596 33793 22624
rect 33744 22584 33750 22596
rect 33781 22593 33793 22596
rect 33827 22593 33839 22627
rect 33781 22587 33839 22593
rect 34057 22627 34115 22633
rect 34057 22593 34069 22627
rect 34103 22593 34115 22627
rect 35802 22624 35808 22636
rect 35763 22596 35808 22624
rect 34057 22587 34115 22593
rect 35802 22584 35808 22596
rect 35860 22584 35866 22636
rect 35894 22584 35900 22636
rect 35952 22624 35958 22636
rect 36372 22633 36400 22664
rect 38841 22661 38853 22695
rect 38887 22692 38899 22695
rect 39114 22692 39120 22704
rect 38887 22664 39120 22692
rect 38887 22661 38899 22664
rect 38841 22655 38899 22661
rect 39114 22652 39120 22664
rect 39172 22692 39178 22704
rect 39485 22695 39543 22701
rect 39485 22692 39497 22695
rect 39172 22664 39497 22692
rect 39172 22652 39178 22664
rect 39485 22661 39497 22664
rect 39531 22692 39543 22695
rect 40405 22695 40463 22701
rect 40405 22692 40417 22695
rect 39531 22664 40417 22692
rect 39531 22661 39543 22664
rect 39485 22655 39543 22661
rect 40405 22661 40417 22664
rect 40451 22661 40463 22695
rect 40405 22655 40463 22661
rect 35989 22627 36047 22633
rect 35989 22624 36001 22627
rect 35952 22596 36001 22624
rect 35952 22584 35958 22596
rect 35989 22593 36001 22596
rect 36035 22593 36047 22627
rect 35989 22587 36047 22593
rect 36357 22627 36415 22633
rect 36357 22593 36369 22627
rect 36403 22593 36415 22627
rect 38470 22624 38476 22636
rect 38431 22596 38476 22624
rect 36357 22587 36415 22593
rect 38470 22584 38476 22596
rect 38528 22584 38534 22636
rect 38657 22627 38715 22633
rect 38657 22593 38669 22627
rect 38703 22624 38715 22627
rect 38930 22624 38936 22636
rect 38703 22596 38936 22624
rect 38703 22593 38715 22596
rect 38657 22587 38715 22593
rect 38930 22584 38936 22596
rect 38988 22584 38994 22636
rect 39298 22624 39304 22636
rect 39259 22596 39304 22624
rect 39298 22584 39304 22596
rect 39356 22584 39362 22636
rect 39574 22624 39580 22636
rect 39535 22596 39580 22624
rect 39574 22584 39580 22596
rect 39632 22584 39638 22636
rect 39669 22627 39727 22633
rect 39669 22593 39681 22627
rect 39715 22624 39727 22627
rect 40034 22624 40040 22636
rect 39715 22596 40040 22624
rect 39715 22593 39727 22596
rect 39669 22587 39727 22593
rect 40034 22584 40040 22596
rect 40092 22584 40098 22636
rect 40313 22627 40371 22633
rect 40313 22593 40325 22627
rect 40359 22593 40371 22627
rect 40313 22587 40371 22593
rect 31904 22528 32352 22556
rect 31904 22516 31910 22528
rect 33134 22516 33140 22568
rect 33192 22556 33198 22568
rect 33965 22559 34023 22565
rect 33965 22556 33977 22559
rect 33192 22528 33977 22556
rect 33192 22516 33198 22528
rect 33965 22525 33977 22528
rect 34011 22525 34023 22559
rect 36078 22556 36084 22568
rect 36039 22528 36084 22556
rect 33965 22519 34023 22525
rect 36078 22516 36084 22528
rect 36136 22516 36142 22568
rect 36170 22516 36176 22568
rect 36228 22556 36234 22568
rect 38948 22556 38976 22584
rect 39206 22556 39212 22568
rect 36228 22528 36273 22556
rect 38948 22528 39212 22556
rect 36228 22516 36234 22528
rect 39206 22516 39212 22528
rect 39264 22516 39270 22568
rect 39316 22556 39344 22584
rect 40328 22556 40356 22587
rect 40586 22584 40592 22636
rect 40644 22624 40650 22636
rect 40681 22627 40739 22633
rect 40681 22624 40693 22627
rect 40644 22596 40693 22624
rect 40644 22584 40650 22596
rect 40681 22593 40693 22596
rect 40727 22593 40739 22627
rect 43070 22624 43076 22636
rect 43031 22596 43076 22624
rect 40681 22587 40739 22593
rect 43070 22584 43076 22596
rect 43128 22584 43134 22636
rect 43806 22584 43812 22636
rect 43864 22624 43870 22636
rect 43973 22627 44031 22633
rect 43973 22624 43985 22627
rect 43864 22596 43985 22624
rect 43864 22584 43870 22596
rect 43973 22593 43985 22596
rect 44019 22593 44031 22627
rect 43973 22587 44031 22593
rect 46017 22627 46075 22633
rect 46017 22593 46029 22627
rect 46063 22624 46075 22627
rect 46290 22624 46296 22636
rect 46063 22596 46296 22624
rect 46063 22593 46075 22596
rect 46017 22587 46075 22593
rect 46290 22584 46296 22596
rect 46348 22624 46354 22636
rect 46842 22624 46848 22636
rect 46348 22596 46848 22624
rect 46348 22584 46354 22596
rect 46842 22584 46848 22596
rect 46900 22584 46906 22636
rect 42886 22556 42892 22568
rect 39316 22528 40356 22556
rect 42847 22528 42892 22556
rect 42886 22516 42892 22528
rect 42944 22516 42950 22568
rect 43717 22559 43775 22565
rect 43717 22525 43729 22559
rect 43763 22525 43775 22559
rect 43717 22519 43775 22525
rect 17221 22491 17279 22497
rect 17221 22457 17233 22491
rect 17267 22488 17279 22491
rect 17773 22491 17831 22497
rect 17773 22488 17785 22491
rect 17267 22460 17785 22488
rect 17267 22457 17279 22460
rect 17221 22451 17279 22457
rect 17773 22457 17785 22460
rect 17819 22457 17831 22491
rect 24210 22488 24216 22500
rect 17773 22451 17831 22457
rect 23584 22460 24216 22488
rect 13170 22380 13176 22432
rect 13228 22420 13234 22432
rect 13633 22423 13691 22429
rect 13633 22420 13645 22423
rect 13228 22392 13645 22420
rect 13228 22380 13234 22392
rect 13633 22389 13645 22392
rect 13679 22389 13691 22423
rect 15562 22420 15568 22432
rect 15523 22392 15568 22420
rect 13633 22383 13691 22389
rect 15562 22380 15568 22392
rect 15620 22380 15626 22432
rect 17313 22423 17371 22429
rect 17313 22389 17325 22423
rect 17359 22420 17371 22423
rect 18046 22420 18052 22432
rect 17359 22392 18052 22420
rect 17359 22389 17371 22392
rect 17313 22383 17371 22389
rect 18046 22380 18052 22392
rect 18104 22380 18110 22432
rect 21726 22380 21732 22432
rect 21784 22420 21790 22432
rect 23584 22429 23612 22460
rect 24210 22448 24216 22460
rect 24268 22448 24274 22500
rect 31665 22491 31723 22497
rect 31665 22457 31677 22491
rect 31711 22488 31723 22491
rect 32858 22488 32864 22500
rect 31711 22460 32864 22488
rect 31711 22457 31723 22460
rect 31665 22451 31723 22457
rect 32858 22448 32864 22460
rect 32916 22448 32922 22500
rect 39853 22491 39911 22497
rect 39853 22457 39865 22491
rect 39899 22488 39911 22491
rect 40218 22488 40224 22500
rect 39899 22460 40224 22488
rect 39899 22457 39911 22460
rect 39853 22451 39911 22457
rect 40218 22448 40224 22460
rect 40276 22448 40282 22500
rect 22281 22423 22339 22429
rect 22281 22420 22293 22423
rect 21784 22392 22293 22420
rect 21784 22380 21790 22392
rect 22281 22389 22293 22392
rect 22327 22389 22339 22423
rect 22281 22383 22339 22389
rect 23569 22423 23627 22429
rect 23569 22389 23581 22423
rect 23615 22389 23627 22423
rect 23569 22383 23627 22389
rect 23658 22380 23664 22432
rect 23716 22420 23722 22432
rect 24029 22423 24087 22429
rect 24029 22420 24041 22423
rect 23716 22392 24041 22420
rect 23716 22380 23722 22392
rect 24029 22389 24041 22392
rect 24075 22389 24087 22423
rect 24029 22383 24087 22389
rect 24394 22380 24400 22432
rect 24452 22420 24458 22432
rect 24581 22423 24639 22429
rect 24581 22420 24593 22423
rect 24452 22392 24593 22420
rect 24452 22380 24458 22392
rect 24581 22389 24593 22392
rect 24627 22389 24639 22423
rect 30558 22420 30564 22432
rect 30471 22392 30564 22420
rect 24581 22383 24639 22389
rect 30558 22380 30564 22392
rect 30616 22420 30622 22432
rect 31386 22420 31392 22432
rect 30616 22392 31392 22420
rect 30616 22380 30622 22392
rect 31386 22380 31392 22392
rect 31444 22380 31450 22432
rect 32674 22420 32680 22432
rect 32635 22392 32680 22420
rect 32674 22380 32680 22392
rect 32732 22380 32738 22432
rect 36538 22420 36544 22432
rect 36499 22392 36544 22420
rect 36538 22380 36544 22392
rect 36596 22380 36602 22432
rect 40034 22380 40040 22432
rect 40092 22420 40098 22432
rect 40405 22423 40463 22429
rect 40405 22420 40417 22423
rect 40092 22392 40417 22420
rect 40092 22380 40098 22392
rect 40405 22389 40417 22392
rect 40451 22389 40463 22423
rect 41506 22420 41512 22432
rect 41467 22392 41512 22420
rect 40405 22383 40463 22389
rect 41506 22380 41512 22392
rect 41564 22380 41570 22432
rect 43257 22423 43315 22429
rect 43257 22389 43269 22423
rect 43303 22420 43315 22423
rect 43622 22420 43628 22432
rect 43303 22392 43628 22420
rect 43303 22389 43315 22392
rect 43257 22383 43315 22389
rect 43622 22380 43628 22392
rect 43680 22380 43686 22432
rect 43732 22420 43760 22519
rect 44358 22420 44364 22432
rect 43732 22392 44364 22420
rect 44358 22380 44364 22392
rect 44416 22380 44422 22432
rect 45097 22423 45155 22429
rect 45097 22389 45109 22423
rect 45143 22420 45155 22423
rect 45462 22420 45468 22432
rect 45143 22392 45468 22420
rect 45143 22389 45155 22392
rect 45097 22383 45155 22389
rect 45462 22380 45468 22392
rect 45520 22380 45526 22432
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 12345 22219 12403 22225
rect 12345 22185 12357 22219
rect 12391 22216 12403 22219
rect 12526 22216 12532 22228
rect 12391 22188 12532 22216
rect 12391 22185 12403 22188
rect 12345 22179 12403 22185
rect 12526 22176 12532 22188
rect 12584 22176 12590 22228
rect 14274 22216 14280 22228
rect 14235 22188 14280 22216
rect 14274 22176 14280 22188
rect 14332 22176 14338 22228
rect 18506 22176 18512 22228
rect 18564 22216 18570 22228
rect 29822 22216 29828 22228
rect 18564 22188 29828 22216
rect 18564 22176 18570 22188
rect 29822 22176 29828 22188
rect 29880 22176 29886 22228
rect 32769 22219 32827 22225
rect 32769 22185 32781 22219
rect 32815 22216 32827 22219
rect 33962 22216 33968 22228
rect 32815 22188 33968 22216
rect 32815 22185 32827 22188
rect 32769 22179 32827 22185
rect 33962 22176 33968 22188
rect 34020 22176 34026 22228
rect 38565 22219 38623 22225
rect 38565 22185 38577 22219
rect 38611 22216 38623 22219
rect 39298 22216 39304 22228
rect 38611 22188 39304 22216
rect 38611 22185 38623 22188
rect 38565 22179 38623 22185
rect 39298 22176 39304 22188
rect 39356 22176 39362 22228
rect 39390 22176 39396 22228
rect 39448 22216 39454 22228
rect 39485 22219 39543 22225
rect 39485 22216 39497 22219
rect 39448 22188 39497 22216
rect 39448 22176 39454 22188
rect 39485 22185 39497 22188
rect 39531 22185 39543 22219
rect 39485 22179 39543 22185
rect 40126 22176 40132 22228
rect 40184 22216 40190 22228
rect 40221 22219 40279 22225
rect 40221 22216 40233 22219
rect 40184 22188 40233 22216
rect 40184 22176 40190 22188
rect 40221 22185 40233 22188
rect 40267 22185 40279 22219
rect 40221 22179 40279 22185
rect 40494 22176 40500 22228
rect 40552 22176 40558 22228
rect 4614 22108 4620 22160
rect 4672 22148 4678 22160
rect 5258 22148 5264 22160
rect 4672 22120 5264 22148
rect 4672 22108 4678 22120
rect 5258 22108 5264 22120
rect 5316 22148 5322 22160
rect 11514 22148 11520 22160
rect 5316 22120 11520 22148
rect 5316 22108 5322 22120
rect 11514 22108 11520 22120
rect 11572 22108 11578 22160
rect 13541 22151 13599 22157
rect 13541 22117 13553 22151
rect 13587 22148 13599 22151
rect 14918 22148 14924 22160
rect 13587 22120 14924 22148
rect 13587 22117 13599 22120
rect 13541 22111 13599 22117
rect 14918 22108 14924 22120
rect 14976 22108 14982 22160
rect 20625 22151 20683 22157
rect 20625 22117 20637 22151
rect 20671 22148 20683 22151
rect 21177 22151 21235 22157
rect 21177 22148 21189 22151
rect 20671 22120 21189 22148
rect 20671 22117 20683 22120
rect 20625 22111 20683 22117
rect 21177 22117 21189 22120
rect 21223 22117 21235 22151
rect 21177 22111 21235 22117
rect 23106 22108 23112 22160
rect 23164 22148 23170 22160
rect 23566 22148 23572 22160
rect 23164 22120 23572 22148
rect 23164 22108 23170 22120
rect 23566 22108 23572 22120
rect 23624 22108 23630 22160
rect 33134 22148 33140 22160
rect 33095 22120 33140 22148
rect 33134 22108 33140 22120
rect 33192 22108 33198 22160
rect 37182 22108 37188 22160
rect 37240 22148 37246 22160
rect 40512 22148 40540 22176
rect 37240 22120 40540 22148
rect 37240 22108 37246 22120
rect 42886 22108 42892 22160
rect 42944 22148 42950 22160
rect 44082 22148 44088 22160
rect 42944 22120 44088 22148
rect 42944 22108 42950 22120
rect 44082 22108 44088 22120
rect 44140 22108 44146 22160
rect 46566 22148 46572 22160
rect 44192 22120 46572 22148
rect 13262 22080 13268 22092
rect 13223 22052 13268 22080
rect 13262 22040 13268 22052
rect 13320 22040 13326 22092
rect 15562 22040 15568 22092
rect 15620 22080 15626 22092
rect 15749 22083 15807 22089
rect 15749 22080 15761 22083
rect 15620 22052 15761 22080
rect 15620 22040 15626 22052
rect 15749 22049 15761 22052
rect 15795 22049 15807 22083
rect 15749 22043 15807 22049
rect 15838 22040 15844 22092
rect 15896 22080 15902 22092
rect 20717 22083 20775 22089
rect 15896 22052 15941 22080
rect 15896 22040 15902 22052
rect 20717 22049 20729 22083
rect 20763 22049 20775 22083
rect 21726 22080 21732 22092
rect 21687 22052 21732 22080
rect 20717 22043 20775 22049
rect 2038 21972 2044 22024
rect 2096 22012 2102 22024
rect 2225 22015 2283 22021
rect 2225 22012 2237 22015
rect 2096 21984 2237 22012
rect 2096 21972 2102 21984
rect 2225 21981 2237 21984
rect 2271 21981 2283 22015
rect 2225 21975 2283 21981
rect 12529 22015 12587 22021
rect 12529 21981 12541 22015
rect 12575 22012 12587 22015
rect 12802 22012 12808 22024
rect 12575 21984 12808 22012
rect 12575 21981 12587 21984
rect 12529 21975 12587 21981
rect 12802 21972 12808 21984
rect 12860 21972 12866 22024
rect 13170 22012 13176 22024
rect 13131 21984 13176 22012
rect 13170 21972 13176 21984
rect 13228 21972 13234 22024
rect 13906 21972 13912 22024
rect 13964 22012 13970 22024
rect 14461 22015 14519 22021
rect 14461 22012 14473 22015
rect 13964 21984 14473 22012
rect 13964 21972 13970 21984
rect 14461 21981 14473 21984
rect 14507 21981 14519 22015
rect 14461 21975 14519 21981
rect 15657 22015 15715 22021
rect 15657 21981 15669 22015
rect 15703 22012 15715 22015
rect 17310 22012 17316 22024
rect 15703 21984 17316 22012
rect 15703 21981 15715 21984
rect 15657 21975 15715 21981
rect 17310 21972 17316 21984
rect 17368 21972 17374 22024
rect 17405 22015 17463 22021
rect 17405 21981 17417 22015
rect 17451 22012 17463 22015
rect 18138 22012 18144 22024
rect 17451 21984 18144 22012
rect 17451 21981 17463 21984
rect 17405 21975 17463 21981
rect 18138 21972 18144 21984
rect 18196 21972 18202 22024
rect 20732 22012 20760 22043
rect 21726 22040 21732 22052
rect 21784 22040 21790 22092
rect 22922 22040 22928 22092
rect 22980 22080 22986 22092
rect 30466 22080 30472 22092
rect 22980 22052 30472 22080
rect 22980 22040 22986 22052
rect 22557 22015 22615 22021
rect 22557 22012 22569 22015
rect 20732 21984 22569 22012
rect 22557 21981 22569 21984
rect 22603 21981 22615 22015
rect 23106 22012 23112 22024
rect 23067 21984 23112 22012
rect 22557 21975 22615 21981
rect 23106 21972 23112 21984
rect 23164 21972 23170 22024
rect 23198 21972 23204 22024
rect 23256 22012 23262 22024
rect 23293 22015 23351 22021
rect 23293 22012 23305 22015
rect 23256 21984 23305 22012
rect 23256 21972 23262 21984
rect 23293 21981 23305 21984
rect 23339 21981 23351 22015
rect 23293 21975 23351 21981
rect 24486 21972 24492 22024
rect 24544 22012 24550 22024
rect 24765 22015 24823 22021
rect 24765 22012 24777 22015
rect 24544 21984 24777 22012
rect 24544 21972 24550 21984
rect 24765 21981 24777 21984
rect 24811 21981 24823 22015
rect 25038 22012 25044 22024
rect 24999 21984 25044 22012
rect 24765 21975 24823 21981
rect 17672 21947 17730 21953
rect 17672 21913 17684 21947
rect 17718 21944 17730 21947
rect 17770 21944 17776 21956
rect 17718 21916 17776 21944
rect 17718 21913 17730 21916
rect 17672 21907 17730 21913
rect 17770 21904 17776 21916
rect 17828 21904 17834 21956
rect 20254 21944 20260 21956
rect 20167 21916 20260 21944
rect 20254 21904 20260 21916
rect 20312 21944 20318 21956
rect 24504 21944 24532 21972
rect 20312 21916 24532 21944
rect 24780 21944 24808 21975
rect 25038 21972 25044 21984
rect 25096 21972 25102 22024
rect 25225 22015 25283 22021
rect 25225 21981 25237 22015
rect 25271 22012 25283 22015
rect 26694 22012 26700 22024
rect 25271 21984 26700 22012
rect 25271 21981 25283 21984
rect 25225 21975 25283 21981
rect 26694 21972 26700 21984
rect 26752 21972 26758 22024
rect 26804 22021 26832 22052
rect 30466 22040 30472 22052
rect 30524 22040 30530 22092
rect 33689 22083 33747 22089
rect 33689 22080 33701 22083
rect 32968 22052 33701 22080
rect 26789 22015 26847 22021
rect 26789 21981 26801 22015
rect 26835 21981 26847 22015
rect 26789 21975 26847 21981
rect 27065 22015 27123 22021
rect 27065 21981 27077 22015
rect 27111 21981 27123 22015
rect 27065 21975 27123 21981
rect 27249 22015 27307 22021
rect 27249 21981 27261 22015
rect 27295 22012 27307 22015
rect 27614 22012 27620 22024
rect 27295 21984 27620 22012
rect 27295 21981 27307 21984
rect 27249 21975 27307 21981
rect 25590 21944 25596 21956
rect 24780 21916 25596 21944
rect 20312 21904 20318 21916
rect 25590 21904 25596 21916
rect 25648 21904 25654 21956
rect 25685 21947 25743 21953
rect 25685 21913 25697 21947
rect 25731 21913 25743 21947
rect 25866 21944 25872 21956
rect 25827 21916 25872 21944
rect 25685 21907 25743 21913
rect 15289 21879 15347 21885
rect 15289 21845 15301 21879
rect 15335 21876 15347 21879
rect 15930 21876 15936 21888
rect 15335 21848 15936 21876
rect 15335 21845 15347 21848
rect 15289 21839 15347 21845
rect 15930 21836 15936 21848
rect 15988 21836 15994 21888
rect 18782 21876 18788 21888
rect 18743 21848 18788 21876
rect 18782 21836 18788 21848
rect 18840 21836 18846 21888
rect 21450 21836 21456 21888
rect 21508 21876 21514 21888
rect 21545 21879 21603 21885
rect 21545 21876 21557 21879
rect 21508 21848 21557 21876
rect 21508 21836 21514 21848
rect 21545 21845 21557 21848
rect 21591 21845 21603 21879
rect 21545 21839 21603 21845
rect 21634 21836 21640 21888
rect 21692 21876 21698 21888
rect 22370 21876 22376 21888
rect 21692 21848 21737 21876
rect 22331 21848 22376 21876
rect 21692 21836 21698 21848
rect 22370 21836 22376 21848
rect 22428 21836 22434 21888
rect 23474 21876 23480 21888
rect 23435 21848 23480 21876
rect 23474 21836 23480 21848
rect 23532 21836 23538 21888
rect 24578 21876 24584 21888
rect 24539 21848 24584 21876
rect 24578 21836 24584 21848
rect 24636 21836 24642 21888
rect 25700 21876 25728 21907
rect 25866 21904 25872 21916
rect 25924 21904 25930 21956
rect 26234 21944 26240 21956
rect 25976 21916 26240 21944
rect 25976 21876 26004 21916
rect 26234 21904 26240 21916
rect 26292 21904 26298 21956
rect 27080 21944 27108 21975
rect 27614 21972 27620 21984
rect 27672 21972 27678 22024
rect 30561 22015 30619 22021
rect 30561 21981 30573 22015
rect 30607 22012 30619 22015
rect 30650 22012 30656 22024
rect 30607 21984 30656 22012
rect 30607 21981 30619 21984
rect 30561 21975 30619 21981
rect 30650 21972 30656 21984
rect 30708 21972 30714 22024
rect 31202 21972 31208 22024
rect 31260 22012 31266 22024
rect 32968 22021 32996 22052
rect 33689 22049 33701 22052
rect 33735 22049 33747 22083
rect 33689 22043 33747 22049
rect 34238 22040 34244 22092
rect 34296 22080 34302 22092
rect 35894 22080 35900 22092
rect 34296 22052 35900 22080
rect 34296 22040 34302 22052
rect 35894 22040 35900 22052
rect 35952 22040 35958 22092
rect 40126 22040 40132 22092
rect 40184 22080 40190 22092
rect 40954 22080 40960 22092
rect 40184 22052 40960 22080
rect 40184 22040 40190 22052
rect 40954 22040 40960 22052
rect 41012 22040 41018 22092
rect 41325 22083 41383 22089
rect 41325 22049 41337 22083
rect 41371 22080 41383 22083
rect 41506 22080 41512 22092
rect 41371 22052 41512 22080
rect 41371 22049 41383 22052
rect 41325 22043 41383 22049
rect 41506 22040 41512 22052
rect 41564 22040 41570 22092
rect 32953 22015 33011 22021
rect 31260 21984 31754 22012
rect 31260 21972 31266 21984
rect 27154 21944 27160 21956
rect 27067 21916 27160 21944
rect 27154 21904 27160 21916
rect 27212 21944 27218 21956
rect 30282 21944 30288 21956
rect 27212 21916 30288 21944
rect 27212 21904 27218 21916
rect 30282 21904 30288 21916
rect 30340 21904 30346 21956
rect 30828 21947 30886 21953
rect 30828 21913 30840 21947
rect 30874 21944 30886 21947
rect 31570 21944 31576 21956
rect 30874 21916 31576 21944
rect 30874 21913 30886 21916
rect 30828 21907 30886 21913
rect 31570 21904 31576 21916
rect 31628 21904 31634 21956
rect 31726 21944 31754 21984
rect 32953 21981 32965 22015
rect 32999 21981 33011 22015
rect 32953 21975 33011 21981
rect 33229 22015 33287 22021
rect 33229 21981 33241 22015
rect 33275 22012 33287 22015
rect 33410 22012 33416 22024
rect 33275 21984 33416 22012
rect 33275 21981 33287 21984
rect 33229 21975 33287 21981
rect 33244 21944 33272 21975
rect 33410 21972 33416 21984
rect 33468 21972 33474 22024
rect 33870 22012 33876 22024
rect 33831 21984 33876 22012
rect 33870 21972 33876 21984
rect 33928 21972 33934 22024
rect 34054 21972 34060 22024
rect 34112 22012 34118 22024
rect 34149 22015 34207 22021
rect 34149 22012 34161 22015
rect 34112 21984 34161 22012
rect 34112 21972 34118 21984
rect 34149 21981 34161 21984
rect 34195 21981 34207 22015
rect 34149 21975 34207 21981
rect 34333 22015 34391 22021
rect 34333 21981 34345 22015
rect 34379 22012 34391 22015
rect 35066 22012 35072 22024
rect 34379 21984 35072 22012
rect 34379 21981 34391 21984
rect 34333 21975 34391 21981
rect 35066 21972 35072 21984
rect 35124 21972 35130 22024
rect 36173 22015 36231 22021
rect 36173 21981 36185 22015
rect 36219 22012 36231 22015
rect 37274 22012 37280 22024
rect 36219 21984 37280 22012
rect 36219 21981 36231 21984
rect 36173 21975 36231 21981
rect 37274 21972 37280 21984
rect 37332 21972 37338 22024
rect 38470 22012 38476 22024
rect 38383 21984 38476 22012
rect 38470 21972 38476 21984
rect 38528 21972 38534 22024
rect 38657 22015 38715 22021
rect 38657 21981 38669 22015
rect 38703 22012 38715 22015
rect 39206 22012 39212 22024
rect 38703 21984 39212 22012
rect 38703 21981 38715 21984
rect 38657 21975 38715 21981
rect 39206 21972 39212 21984
rect 39264 21972 39270 22024
rect 39301 22015 39359 22021
rect 39301 21981 39313 22015
rect 39347 22012 39359 22015
rect 39758 22012 39764 22024
rect 39347 21984 39764 22012
rect 39347 21981 39359 21984
rect 39301 21975 39359 21981
rect 31726 21916 33272 21944
rect 36440 21947 36498 21953
rect 36440 21913 36452 21947
rect 36486 21944 36498 21947
rect 36538 21944 36544 21956
rect 36486 21916 36544 21944
rect 36486 21913 36498 21916
rect 36440 21907 36498 21913
rect 36538 21904 36544 21916
rect 36596 21904 36602 21956
rect 38488 21944 38516 21972
rect 39316 21944 39344 21975
rect 39758 21972 39764 21984
rect 39816 22012 39822 22024
rect 41046 22012 41052 22024
rect 39816 21984 41052 22012
rect 39816 21972 39822 21984
rect 41046 21972 41052 21984
rect 41104 21972 41110 22024
rect 43165 22015 43223 22021
rect 43165 21981 43177 22015
rect 43211 22012 43223 22015
rect 44192 22012 44220 22120
rect 46566 22108 46572 22120
rect 46624 22108 46630 22160
rect 44269 22083 44327 22089
rect 44269 22049 44281 22083
rect 44315 22080 44327 22083
rect 45922 22080 45928 22092
rect 44315 22052 45928 22080
rect 44315 22049 44327 22052
rect 44269 22043 44327 22049
rect 45922 22040 45928 22052
rect 45980 22040 45986 22092
rect 46382 22080 46388 22092
rect 46343 22052 46388 22080
rect 46382 22040 46388 22052
rect 46440 22040 46446 22092
rect 46658 22080 46664 22092
rect 46619 22052 46664 22080
rect 46658 22040 46664 22052
rect 46716 22040 46722 22092
rect 43211 21984 44220 22012
rect 45373 22015 45431 22021
rect 43211 21981 43223 21984
rect 43165 21975 43223 21981
rect 45373 21981 45385 22015
rect 45419 21981 45431 22015
rect 45373 21975 45431 21981
rect 40034 21944 40040 21956
rect 38488 21916 39344 21944
rect 39995 21916 40040 21944
rect 40034 21904 40040 21916
rect 40092 21904 40098 21956
rect 40218 21904 40224 21956
rect 40276 21953 40282 21956
rect 40276 21947 40295 21953
rect 40283 21913 40295 21947
rect 40276 21907 40295 21913
rect 40276 21904 40282 21907
rect 40862 21904 40868 21956
rect 40920 21944 40926 21956
rect 41509 21947 41567 21953
rect 41509 21944 41521 21947
rect 40920 21916 41521 21944
rect 40920 21904 40926 21916
rect 41509 21913 41521 21916
rect 41555 21913 41567 21947
rect 45388 21944 45416 21975
rect 45462 21972 45468 22024
rect 45520 22012 45526 22024
rect 46201 22015 46259 22021
rect 46201 22012 46213 22015
rect 45520 21984 46213 22012
rect 45520 21972 45526 21984
rect 46201 21981 46213 21984
rect 46247 21981 46259 22015
rect 46201 21975 46259 21981
rect 41509 21907 41567 21913
rect 43640 21916 45416 21944
rect 25700 21848 26004 21876
rect 26053 21879 26111 21885
rect 26053 21845 26065 21879
rect 26099 21876 26111 21879
rect 26142 21876 26148 21888
rect 26099 21848 26148 21876
rect 26099 21845 26111 21848
rect 26053 21839 26111 21845
rect 26142 21836 26148 21848
rect 26200 21836 26206 21888
rect 26605 21879 26663 21885
rect 26605 21845 26617 21879
rect 26651 21876 26663 21879
rect 27338 21876 27344 21888
rect 26651 21848 27344 21876
rect 26651 21845 26663 21848
rect 26605 21839 26663 21845
rect 27338 21836 27344 21848
rect 27396 21836 27402 21888
rect 31110 21836 31116 21888
rect 31168 21876 31174 21888
rect 31846 21876 31852 21888
rect 31168 21848 31852 21876
rect 31168 21836 31174 21848
rect 31846 21836 31852 21848
rect 31904 21876 31910 21888
rect 31941 21879 31999 21885
rect 31941 21876 31953 21879
rect 31904 21848 31953 21876
rect 31904 21836 31910 21848
rect 31941 21845 31953 21848
rect 31987 21845 31999 21879
rect 31941 21839 31999 21845
rect 36078 21836 36084 21888
rect 36136 21876 36142 21888
rect 36722 21876 36728 21888
rect 36136 21848 36728 21876
rect 36136 21836 36142 21848
rect 36722 21836 36728 21848
rect 36780 21876 36786 21888
rect 37553 21879 37611 21885
rect 37553 21876 37565 21879
rect 36780 21848 37565 21876
rect 36780 21836 36786 21848
rect 37553 21845 37565 21848
rect 37599 21845 37611 21879
rect 37553 21839 37611 21845
rect 39482 21836 39488 21888
rect 39540 21876 39546 21888
rect 43640 21885 43668 21916
rect 40405 21879 40463 21885
rect 40405 21876 40417 21879
rect 39540 21848 40417 21876
rect 39540 21836 39546 21848
rect 40405 21845 40417 21848
rect 40451 21845 40463 21879
rect 40405 21839 40463 21845
rect 43625 21879 43683 21885
rect 43625 21845 43637 21879
rect 43671 21845 43683 21879
rect 43990 21876 43996 21888
rect 43951 21848 43996 21876
rect 43625 21839 43683 21845
rect 43990 21836 43996 21848
rect 44048 21836 44054 21888
rect 44082 21836 44088 21888
rect 44140 21876 44146 21888
rect 45186 21876 45192 21888
rect 44140 21848 44185 21876
rect 45147 21848 45192 21876
rect 44140 21836 44146 21848
rect 45186 21836 45192 21848
rect 45244 21836 45250 21888
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 13262 21672 13268 21684
rect 13223 21644 13268 21672
rect 13262 21632 13268 21644
rect 13320 21632 13326 21684
rect 13906 21672 13912 21684
rect 13867 21644 13912 21672
rect 13906 21632 13912 21644
rect 13964 21632 13970 21684
rect 17770 21672 17776 21684
rect 17731 21644 17776 21672
rect 17770 21632 17776 21644
rect 17828 21632 17834 21684
rect 21450 21672 21456 21684
rect 19904 21644 21456 21672
rect 13170 21564 13176 21616
rect 13228 21604 13234 21616
rect 14369 21607 14427 21613
rect 14369 21604 14381 21607
rect 13228 21576 14381 21604
rect 13228 21564 13234 21576
rect 14369 21573 14381 21576
rect 14415 21573 14427 21607
rect 14369 21567 14427 21573
rect 15933 21607 15991 21613
rect 15933 21573 15945 21607
rect 15979 21604 15991 21607
rect 19904 21604 19932 21644
rect 21450 21632 21456 21644
rect 21508 21632 21514 21684
rect 21634 21632 21640 21684
rect 21692 21672 21698 21684
rect 25225 21675 25283 21681
rect 21692 21644 25176 21672
rect 21692 21632 21698 21644
rect 20622 21604 20628 21616
rect 15979 21576 19932 21604
rect 20088 21576 20628 21604
rect 15979 21573 15991 21576
rect 15933 21567 15991 21573
rect 2038 21536 2044 21548
rect 1999 21508 2044 21536
rect 2038 21496 2044 21508
rect 2096 21496 2102 21548
rect 9582 21536 9588 21548
rect 9543 21508 9588 21536
rect 9582 21496 9588 21508
rect 9640 21496 9646 21548
rect 10410 21536 10416 21548
rect 10371 21508 10416 21536
rect 10410 21496 10416 21508
rect 10468 21496 10474 21548
rect 12152 21539 12210 21545
rect 12152 21505 12164 21539
rect 12198 21536 12210 21539
rect 12434 21536 12440 21548
rect 12198 21508 12440 21536
rect 12198 21505 12210 21508
rect 12152 21499 12210 21505
rect 12434 21496 12440 21508
rect 12492 21496 12498 21548
rect 14277 21539 14335 21545
rect 14277 21505 14289 21539
rect 14323 21536 14335 21539
rect 17957 21539 18015 21545
rect 14323 21508 16574 21536
rect 14323 21505 14335 21508
rect 14277 21499 14335 21505
rect 2225 21471 2283 21477
rect 2225 21437 2237 21471
rect 2271 21468 2283 21471
rect 2314 21468 2320 21480
rect 2271 21440 2320 21468
rect 2271 21437 2283 21440
rect 2225 21431 2283 21437
rect 2314 21428 2320 21440
rect 2372 21428 2378 21480
rect 2774 21468 2780 21480
rect 2735 21440 2780 21468
rect 2774 21428 2780 21440
rect 2832 21428 2838 21480
rect 9677 21471 9735 21477
rect 9677 21437 9689 21471
rect 9723 21468 9735 21471
rect 10318 21468 10324 21480
rect 9723 21440 10324 21468
rect 9723 21437 9735 21440
rect 9677 21431 9735 21437
rect 10318 21428 10324 21440
rect 10376 21428 10382 21480
rect 11885 21471 11943 21477
rect 11885 21437 11897 21471
rect 11931 21437 11943 21471
rect 11885 21431 11943 21437
rect 9953 21403 10011 21409
rect 9953 21369 9965 21403
rect 9999 21400 10011 21403
rect 10042 21400 10048 21412
rect 9999 21372 10048 21400
rect 9999 21369 10011 21372
rect 9953 21363 10011 21369
rect 10042 21360 10048 21372
rect 10100 21360 10106 21412
rect 10226 21292 10232 21344
rect 10284 21332 10290 21344
rect 10505 21335 10563 21341
rect 10505 21332 10517 21335
rect 10284 21304 10517 21332
rect 10284 21292 10290 21304
rect 10505 21301 10517 21304
rect 10551 21301 10563 21335
rect 11900 21332 11928 21431
rect 13354 21428 13360 21480
rect 13412 21468 13418 21480
rect 14461 21471 14519 21477
rect 14461 21468 14473 21471
rect 13412 21440 14473 21468
rect 13412 21428 13418 21440
rect 14461 21437 14473 21440
rect 14507 21468 14519 21471
rect 15838 21468 15844 21480
rect 14507 21440 15844 21468
rect 14507 21437 14519 21440
rect 14461 21431 14519 21437
rect 15838 21428 15844 21440
rect 15896 21428 15902 21480
rect 16022 21468 16028 21480
rect 15983 21440 16028 21468
rect 16022 21428 16028 21440
rect 16080 21428 16086 21480
rect 16117 21471 16175 21477
rect 16117 21437 16129 21471
rect 16163 21437 16175 21471
rect 16546 21468 16574 21508
rect 17957 21505 17969 21539
rect 18003 21536 18015 21539
rect 18046 21536 18052 21548
rect 18003 21508 18052 21536
rect 18003 21505 18015 21508
rect 17957 21499 18015 21505
rect 18046 21496 18052 21508
rect 18104 21496 18110 21548
rect 20088 21545 20116 21576
rect 20622 21564 20628 21576
rect 20680 21604 20686 21616
rect 24112 21607 24170 21613
rect 20680 21576 23888 21604
rect 20680 21564 20686 21576
rect 23860 21548 23888 21576
rect 24112 21573 24124 21607
rect 24158 21604 24170 21607
rect 24578 21604 24584 21616
rect 24158 21576 24584 21604
rect 24158 21573 24170 21576
rect 24112 21567 24170 21573
rect 24578 21564 24584 21576
rect 24636 21564 24642 21616
rect 25148 21604 25176 21644
rect 25225 21641 25237 21675
rect 25271 21672 25283 21675
rect 25866 21672 25872 21684
rect 25271 21644 25872 21672
rect 25271 21641 25283 21644
rect 25225 21635 25283 21641
rect 25866 21632 25872 21644
rect 25924 21632 25930 21684
rect 31202 21672 31208 21684
rect 25976 21644 31208 21672
rect 25976 21604 26004 21644
rect 31202 21632 31208 21644
rect 31260 21632 31266 21684
rect 31570 21672 31576 21684
rect 31531 21644 31576 21672
rect 31570 21632 31576 21644
rect 31628 21632 31634 21684
rect 35618 21632 35624 21684
rect 35676 21672 35682 21684
rect 40862 21672 40868 21684
rect 35676 21644 40540 21672
rect 40823 21644 40868 21672
rect 35676 21632 35682 21644
rect 25148 21576 26004 21604
rect 27172 21576 28994 21604
rect 20073 21539 20131 21545
rect 20073 21505 20085 21539
rect 20119 21505 20131 21539
rect 20073 21499 20131 21505
rect 20340 21539 20398 21545
rect 20340 21505 20352 21539
rect 20386 21536 20398 21539
rect 22370 21536 22376 21548
rect 20386 21508 22376 21536
rect 20386 21505 20398 21508
rect 20340 21499 20398 21505
rect 22370 21496 22376 21508
rect 22428 21496 22434 21548
rect 23109 21539 23167 21545
rect 23109 21505 23121 21539
rect 23155 21536 23167 21539
rect 23658 21536 23664 21548
rect 23155 21508 23664 21536
rect 23155 21505 23167 21508
rect 23109 21499 23167 21505
rect 23658 21496 23664 21508
rect 23716 21496 23722 21548
rect 23842 21536 23848 21548
rect 23755 21508 23848 21536
rect 23842 21496 23848 21508
rect 23900 21496 23906 21548
rect 25866 21536 25872 21548
rect 25827 21508 25872 21536
rect 25866 21496 25872 21508
rect 25924 21496 25930 21548
rect 26234 21536 26240 21548
rect 26195 21508 26240 21536
rect 26234 21496 26240 21508
rect 26292 21496 26298 21548
rect 27172 21545 27200 21576
rect 28966 21548 28994 21576
rect 30650 21564 30656 21616
rect 30708 21604 30714 21616
rect 33778 21604 33784 21616
rect 30708 21576 33784 21604
rect 30708 21564 30714 21576
rect 27157 21539 27215 21545
rect 27157 21505 27169 21539
rect 27203 21505 27215 21539
rect 27157 21499 27215 21505
rect 27246 21496 27252 21548
rect 27304 21536 27310 21548
rect 27413 21539 27471 21545
rect 27413 21536 27425 21539
rect 27304 21508 27425 21536
rect 27304 21496 27310 21508
rect 27413 21505 27425 21508
rect 27459 21505 27471 21539
rect 27413 21499 27471 21505
rect 28166 21496 28172 21548
rect 28224 21536 28230 21548
rect 28718 21536 28724 21548
rect 28224 21508 28724 21536
rect 28224 21496 28230 21508
rect 28718 21496 28724 21508
rect 28776 21496 28782 21548
rect 28966 21506 29000 21548
rect 29052 21545 29058 21548
rect 29270 21545 29276 21548
rect 28994 21496 29000 21506
rect 29052 21536 29062 21545
rect 29253 21539 29276 21545
rect 29052 21508 29145 21536
rect 29052 21499 29062 21508
rect 29253 21505 29265 21539
rect 29253 21499 29276 21505
rect 29052 21496 29058 21499
rect 29270 21496 29276 21499
rect 29328 21496 29334 21548
rect 30837 21539 30895 21545
rect 30837 21505 30849 21539
rect 30883 21505 30895 21539
rect 31018 21536 31024 21548
rect 30979 21508 31024 21536
rect 30837 21499 30895 21505
rect 18782 21468 18788 21480
rect 16546 21440 18788 21468
rect 16117 21431 16175 21437
rect 15856 21400 15884 21428
rect 16132 21400 16160 21431
rect 18782 21428 18788 21440
rect 18840 21428 18846 21480
rect 25222 21428 25228 21480
rect 25280 21468 25286 21480
rect 26421 21471 26479 21477
rect 26421 21468 26433 21471
rect 25280 21440 26433 21468
rect 25280 21428 25286 21440
rect 26421 21437 26433 21440
rect 26467 21468 26479 21471
rect 26467 21440 27200 21468
rect 26467 21437 26479 21440
rect 26421 21431 26479 21437
rect 15856 21372 16160 21400
rect 12158 21332 12164 21344
rect 11900 21304 12164 21332
rect 10505 21295 10563 21301
rect 12158 21292 12164 21304
rect 12216 21292 12222 21344
rect 13814 21292 13820 21344
rect 13872 21332 13878 21344
rect 15565 21335 15623 21341
rect 15565 21332 15577 21335
rect 13872 21304 15577 21332
rect 13872 21292 13878 21304
rect 15565 21301 15577 21304
rect 15611 21301 15623 21335
rect 15565 21295 15623 21301
rect 23106 21292 23112 21344
rect 23164 21332 23170 21344
rect 23293 21335 23351 21341
rect 23293 21332 23305 21335
rect 23164 21304 23305 21332
rect 23164 21292 23170 21304
rect 23293 21301 23305 21304
rect 23339 21301 23351 21335
rect 27172 21332 27200 21440
rect 28184 21440 28994 21468
rect 28184 21332 28212 21440
rect 28966 21412 28994 21440
rect 28966 21372 29000 21412
rect 28994 21360 29000 21372
rect 29052 21360 29058 21412
rect 30852 21400 30880 21499
rect 31018 21496 31024 21508
rect 31076 21496 31082 21548
rect 31110 21496 31116 21548
rect 31168 21536 31174 21548
rect 31386 21536 31392 21548
rect 31168 21508 31213 21536
rect 31347 21508 31392 21536
rect 31168 21496 31174 21508
rect 31386 21496 31392 21508
rect 31444 21496 31450 21548
rect 32950 21536 32956 21548
rect 32911 21508 32956 21536
rect 32950 21496 32956 21508
rect 33008 21496 33014 21548
rect 33134 21536 33140 21548
rect 33095 21508 33140 21536
rect 33134 21496 33140 21508
rect 33192 21496 33198 21548
rect 33226 21496 33232 21548
rect 33284 21536 33290 21548
rect 33704 21545 33732 21576
rect 33778 21564 33784 21576
rect 33836 21564 33842 21616
rect 33962 21613 33968 21616
rect 33956 21604 33968 21613
rect 33923 21576 33968 21604
rect 33956 21567 33968 21576
rect 33962 21564 33968 21567
rect 34020 21564 34026 21616
rect 39850 21604 39856 21616
rect 39811 21576 39856 21604
rect 39850 21564 39856 21576
rect 39908 21564 39914 21616
rect 40512 21604 40540 21644
rect 40862 21632 40868 21644
rect 40920 21632 40926 21684
rect 42797 21675 42855 21681
rect 42797 21641 42809 21675
rect 42843 21672 42855 21675
rect 43070 21672 43076 21684
rect 42843 21644 43076 21672
rect 42843 21641 42855 21644
rect 42797 21635 42855 21641
rect 43070 21632 43076 21644
rect 43128 21632 43134 21684
rect 43717 21675 43775 21681
rect 43717 21641 43729 21675
rect 43763 21672 43775 21675
rect 43806 21672 43812 21684
rect 43763 21644 43812 21672
rect 43763 21641 43775 21644
rect 43717 21635 43775 21641
rect 43806 21632 43812 21644
rect 43864 21632 43870 21684
rect 45741 21675 45799 21681
rect 45741 21641 45753 21675
rect 45787 21672 45799 21675
rect 45922 21672 45928 21684
rect 45787 21644 45928 21672
rect 45787 21641 45799 21644
rect 45741 21635 45799 21641
rect 45922 21632 45928 21644
rect 45980 21632 45986 21684
rect 44628 21607 44686 21613
rect 40512 21576 44588 21604
rect 33689 21539 33747 21545
rect 33284 21508 33329 21536
rect 33284 21496 33290 21508
rect 33689 21505 33701 21539
rect 33735 21505 33747 21539
rect 36170 21536 36176 21548
rect 33689 21499 33747 21505
rect 33796 21508 36176 21536
rect 31202 21468 31208 21480
rect 31163 21440 31208 21468
rect 31202 21428 31208 21440
rect 31260 21468 31266 21480
rect 33796 21468 33824 21508
rect 36170 21496 36176 21508
rect 36228 21536 36234 21548
rect 37182 21536 37188 21548
rect 36228 21508 37188 21536
rect 36228 21496 36234 21508
rect 37182 21496 37188 21508
rect 37240 21496 37246 21548
rect 39482 21496 39488 21548
rect 39540 21536 39546 21548
rect 39758 21545 39764 21546
rect 39584 21539 39642 21545
rect 39584 21536 39596 21539
rect 39540 21508 39596 21536
rect 39540 21496 39546 21508
rect 39584 21505 39596 21508
rect 39630 21505 39642 21539
rect 39584 21499 39642 21505
rect 39725 21539 39764 21545
rect 39725 21505 39737 21539
rect 39725 21499 39764 21505
rect 39758 21494 39764 21499
rect 39816 21494 39822 21546
rect 39945 21539 40003 21545
rect 39945 21505 39957 21539
rect 39991 21505 40003 21539
rect 39945 21499 40003 21505
rect 40083 21539 40141 21545
rect 40083 21505 40095 21539
rect 40129 21536 40141 21539
rect 40586 21536 40592 21548
rect 40129 21508 40592 21536
rect 40129 21505 40141 21508
rect 40083 21499 40141 21505
rect 31260 21440 33824 21468
rect 31260 21428 31266 21440
rect 32769 21403 32827 21409
rect 32769 21400 32781 21403
rect 30852 21372 32781 21400
rect 32769 21369 32781 21372
rect 32815 21369 32827 21403
rect 35066 21400 35072 21412
rect 34979 21372 35072 21400
rect 32769 21363 32827 21369
rect 35066 21360 35072 21372
rect 35124 21400 35130 21412
rect 39960 21400 39988 21499
rect 40586 21496 40592 21508
rect 40644 21496 40650 21548
rect 40770 21496 40776 21548
rect 40828 21536 40834 21548
rect 42981 21539 43039 21545
rect 40828 21508 40873 21536
rect 40828 21496 40834 21508
rect 42981 21505 42993 21539
rect 43027 21536 43039 21539
rect 43070 21536 43076 21548
rect 43027 21508 43076 21536
rect 43027 21505 43039 21508
rect 42981 21499 43039 21505
rect 43070 21496 43076 21508
rect 43128 21496 43134 21548
rect 43165 21539 43223 21545
rect 43165 21505 43177 21539
rect 43211 21505 43223 21539
rect 43165 21499 43223 21505
rect 43257 21539 43315 21545
rect 43257 21505 43269 21539
rect 43303 21536 43315 21539
rect 43346 21536 43352 21548
rect 43303 21508 43352 21536
rect 43303 21505 43315 21508
rect 43257 21499 43315 21505
rect 42794 21468 42800 21480
rect 40880 21440 42800 21468
rect 35124 21372 39988 21400
rect 35124 21360 35130 21372
rect 40586 21360 40592 21412
rect 40644 21400 40650 21412
rect 40880 21400 40908 21440
rect 42794 21428 42800 21440
rect 42852 21428 42858 21480
rect 40644 21372 40908 21400
rect 40644 21360 40650 21372
rect 40954 21360 40960 21412
rect 41012 21400 41018 21412
rect 43180 21400 43208 21499
rect 43346 21496 43352 21508
rect 43404 21496 43410 21548
rect 43622 21496 43628 21548
rect 43680 21536 43686 21548
rect 43901 21539 43959 21545
rect 43901 21536 43913 21539
rect 43680 21508 43913 21536
rect 43680 21496 43686 21508
rect 43901 21505 43913 21508
rect 43947 21505 43959 21539
rect 44358 21536 44364 21548
rect 44319 21508 44364 21536
rect 43901 21499 43959 21505
rect 44358 21496 44364 21508
rect 44416 21496 44422 21548
rect 44560 21536 44588 21576
rect 44628 21573 44640 21607
rect 44674 21604 44686 21607
rect 45186 21604 45192 21616
rect 44674 21576 45192 21604
rect 44674 21573 44686 21576
rect 44628 21567 44686 21573
rect 45186 21564 45192 21576
rect 45244 21564 45250 21616
rect 47026 21536 47032 21548
rect 44560 21508 47032 21536
rect 47026 21496 47032 21508
rect 47084 21496 47090 21548
rect 43438 21400 43444 21412
rect 41012 21372 43444 21400
rect 41012 21360 41018 21372
rect 43438 21360 43444 21372
rect 43496 21360 43502 21412
rect 28534 21332 28540 21344
rect 27172 21304 28212 21332
rect 28495 21304 28540 21332
rect 23293 21295 23351 21301
rect 28534 21292 28540 21304
rect 28592 21292 28598 21344
rect 28902 21292 28908 21344
rect 28960 21332 28966 21344
rect 30377 21335 30435 21341
rect 30377 21332 30389 21335
rect 28960 21304 30389 21332
rect 28960 21292 28966 21304
rect 30377 21301 30389 21304
rect 30423 21301 30435 21335
rect 30377 21295 30435 21301
rect 32950 21292 32956 21344
rect 33008 21332 33014 21344
rect 36262 21332 36268 21344
rect 33008 21304 36268 21332
rect 33008 21292 33014 21304
rect 36262 21292 36268 21304
rect 36320 21292 36326 21344
rect 38102 21292 38108 21344
rect 38160 21332 38166 21344
rect 38562 21332 38568 21344
rect 38160 21304 38568 21332
rect 38160 21292 38166 21304
rect 38562 21292 38568 21304
rect 38620 21332 38626 21344
rect 38930 21332 38936 21344
rect 38620 21304 38936 21332
rect 38620 21292 38626 21304
rect 38930 21292 38936 21304
rect 38988 21292 38994 21344
rect 40221 21335 40279 21341
rect 40221 21301 40233 21335
rect 40267 21332 40279 21335
rect 40310 21332 40316 21344
rect 40267 21304 40316 21332
rect 40267 21301 40279 21304
rect 40221 21295 40279 21301
rect 40310 21292 40316 21304
rect 40368 21292 40374 21344
rect 46658 21292 46664 21344
rect 46716 21332 46722 21344
rect 47121 21335 47179 21341
rect 47121 21332 47133 21335
rect 46716 21304 47133 21332
rect 46716 21292 46722 21304
rect 47121 21301 47133 21304
rect 47167 21301 47179 21335
rect 47946 21332 47952 21344
rect 47907 21304 47952 21332
rect 47121 21295 47179 21301
rect 47946 21292 47952 21304
rect 48004 21292 48010 21344
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 2314 21128 2320 21140
rect 2275 21100 2320 21128
rect 2314 21088 2320 21100
rect 2372 21088 2378 21140
rect 12802 21128 12808 21140
rect 12763 21100 12808 21128
rect 12802 21088 12808 21100
rect 12860 21088 12866 21140
rect 16022 21088 16028 21140
rect 16080 21128 16086 21140
rect 16669 21131 16727 21137
rect 16669 21128 16681 21131
rect 16080 21100 16681 21128
rect 16080 21088 16086 21100
rect 16669 21097 16681 21100
rect 16715 21097 16727 21131
rect 16669 21091 16727 21097
rect 24581 21131 24639 21137
rect 24581 21097 24593 21131
rect 24627 21128 24639 21131
rect 25038 21128 25044 21140
rect 24627 21100 25044 21128
rect 24627 21097 24639 21100
rect 24581 21091 24639 21097
rect 25038 21088 25044 21100
rect 25096 21088 25102 21140
rect 27154 21128 27160 21140
rect 27115 21100 27160 21128
rect 27154 21088 27160 21100
rect 27212 21088 27218 21140
rect 28905 21131 28963 21137
rect 28905 21097 28917 21131
rect 28951 21128 28963 21131
rect 29270 21128 29276 21140
rect 28951 21100 29276 21128
rect 28951 21097 28963 21100
rect 28905 21091 28963 21097
rect 29270 21088 29276 21100
rect 29328 21088 29334 21140
rect 33226 21088 33232 21140
rect 33284 21128 33290 21140
rect 34057 21131 34115 21137
rect 34057 21128 34069 21131
rect 33284 21100 34069 21128
rect 33284 21088 33290 21100
rect 34057 21097 34069 21100
rect 34103 21097 34115 21131
rect 34057 21091 34115 21097
rect 38304 21100 41000 21128
rect 6886 21032 10548 21060
rect 2225 20927 2283 20933
rect 2225 20893 2237 20927
rect 2271 20924 2283 20927
rect 2314 20924 2320 20936
rect 2271 20896 2320 20924
rect 2271 20893 2283 20896
rect 2225 20887 2283 20893
rect 2314 20884 2320 20896
rect 2372 20884 2378 20936
rect 4154 20884 4160 20936
rect 4212 20924 4218 20936
rect 4525 20927 4583 20933
rect 4525 20924 4537 20927
rect 4212 20896 4537 20924
rect 4212 20884 4218 20896
rect 4525 20893 4537 20896
rect 4571 20893 4583 20927
rect 4525 20887 4583 20893
rect 3510 20816 3516 20868
rect 3568 20856 3574 20868
rect 6886 20856 6914 21032
rect 10226 20992 10232 21004
rect 10187 20964 10232 20992
rect 10226 20952 10232 20964
rect 10284 20952 10290 21004
rect 10520 21001 10548 21032
rect 23474 21020 23480 21072
rect 23532 21060 23538 21072
rect 23532 21032 25084 21060
rect 23532 21020 23538 21032
rect 10505 20995 10563 21001
rect 10505 20961 10517 20995
rect 10551 20961 10563 20995
rect 13262 20992 13268 21004
rect 13223 20964 13268 20992
rect 10505 20955 10563 20961
rect 13262 20952 13268 20964
rect 13320 20952 13326 21004
rect 13354 20952 13360 21004
rect 13412 20992 13418 21004
rect 23842 20992 23848 21004
rect 13412 20964 13457 20992
rect 23803 20964 23848 20992
rect 13412 20952 13418 20964
rect 23842 20952 23848 20964
rect 23900 20952 23906 21004
rect 24320 20964 24992 20992
rect 10042 20924 10048 20936
rect 10003 20896 10048 20924
rect 10042 20884 10048 20896
rect 10100 20884 10106 20936
rect 12158 20884 12164 20936
rect 12216 20924 12222 20936
rect 15289 20927 15347 20933
rect 15289 20924 15301 20927
rect 12216 20896 15301 20924
rect 12216 20884 12222 20896
rect 15289 20893 15301 20896
rect 15335 20893 15347 20927
rect 19978 20924 19984 20936
rect 19939 20896 19984 20924
rect 15289 20887 15347 20893
rect 19978 20884 19984 20896
rect 20036 20884 20042 20936
rect 23382 20884 23388 20936
rect 23440 20924 23446 20936
rect 24320 20924 24348 20964
rect 23440 20896 24348 20924
rect 23440 20884 23446 20896
rect 24394 20884 24400 20936
rect 24452 20924 24458 20936
rect 24964 20933 24992 20964
rect 25056 20933 25084 21032
rect 28350 21020 28356 21072
rect 28408 21060 28414 21072
rect 31018 21060 31024 21072
rect 28408 21032 31024 21060
rect 28408 21020 28414 21032
rect 31018 21020 31024 21032
rect 31076 21060 31082 21072
rect 34238 21060 34244 21072
rect 31076 21032 34244 21060
rect 31076 21020 31082 21032
rect 34238 21020 34244 21032
rect 34296 21020 34302 21072
rect 30374 20992 30380 21004
rect 26068 20964 30380 20992
rect 24857 20927 24915 20933
rect 24857 20924 24869 20927
rect 24452 20896 24869 20924
rect 24452 20884 24458 20896
rect 24857 20893 24869 20896
rect 24903 20893 24915 20927
rect 24857 20887 24915 20893
rect 24949 20927 25007 20933
rect 24949 20893 24961 20927
rect 24995 20893 25007 20927
rect 24949 20887 25007 20893
rect 25041 20927 25099 20933
rect 25041 20893 25053 20927
rect 25087 20893 25099 20927
rect 25041 20887 25099 20893
rect 25225 20927 25283 20933
rect 25225 20893 25237 20927
rect 25271 20924 25283 20927
rect 25866 20924 25872 20936
rect 25271 20896 25872 20924
rect 25271 20893 25283 20896
rect 25225 20887 25283 20893
rect 25866 20884 25872 20896
rect 25924 20884 25930 20936
rect 3568 20828 6914 20856
rect 3568 20816 3574 20828
rect 15194 20816 15200 20868
rect 15252 20856 15258 20868
rect 15534 20859 15592 20865
rect 15534 20856 15546 20859
rect 15252 20828 15546 20856
rect 15252 20816 15258 20828
rect 15534 20825 15546 20828
rect 15580 20825 15592 20859
rect 15534 20819 15592 20825
rect 22094 20816 22100 20868
rect 22152 20856 22158 20868
rect 23109 20859 23167 20865
rect 23109 20856 23121 20859
rect 22152 20828 23121 20856
rect 22152 20816 22158 20828
rect 23109 20825 23121 20828
rect 23155 20856 23167 20859
rect 26068 20856 26096 20964
rect 30374 20952 30380 20964
rect 30432 20952 30438 21004
rect 31386 20952 31392 21004
rect 31444 20992 31450 21004
rect 38304 20992 38332 21100
rect 40972 21060 41000 21100
rect 41046 21088 41052 21140
rect 41104 21128 41110 21140
rect 41417 21131 41475 21137
rect 41417 21128 41429 21131
rect 41104 21100 41429 21128
rect 41104 21088 41110 21100
rect 41417 21097 41429 21100
rect 41463 21097 41475 21131
rect 41417 21091 41475 21097
rect 42797 21131 42855 21137
rect 42797 21097 42809 21131
rect 42843 21128 42855 21131
rect 42886 21128 42892 21140
rect 42843 21100 42892 21128
rect 42843 21097 42855 21100
rect 42797 21091 42855 21097
rect 42886 21088 42892 21100
rect 42944 21088 42950 21140
rect 43438 21128 43444 21140
rect 43399 21100 43444 21128
rect 43438 21088 43444 21100
rect 43496 21088 43502 21140
rect 43625 21131 43683 21137
rect 43625 21097 43637 21131
rect 43671 21128 43683 21131
rect 43990 21128 43996 21140
rect 43671 21100 43996 21128
rect 43671 21097 43683 21100
rect 43625 21091 43683 21097
rect 43990 21088 43996 21100
rect 44048 21088 44054 21140
rect 48038 21128 48044 21140
rect 44744 21100 48044 21128
rect 44744 21060 44772 21100
rect 48038 21088 48044 21100
rect 48096 21088 48102 21140
rect 47946 21060 47952 21072
rect 40972 21032 44772 21060
rect 46492 21032 47952 21060
rect 31444 20964 38332 20992
rect 31444 20952 31450 20964
rect 26142 20884 26148 20936
rect 26200 20924 26206 20936
rect 28166 20924 28172 20936
rect 26200 20896 26245 20924
rect 28127 20896 28172 20924
rect 26200 20884 26206 20896
rect 28166 20884 28172 20896
rect 28224 20884 28230 20936
rect 28350 20924 28356 20936
rect 28311 20896 28356 20924
rect 28350 20884 28356 20896
rect 28408 20884 28414 20936
rect 28445 20927 28503 20933
rect 28445 20893 28457 20927
rect 28491 20893 28503 20927
rect 28445 20887 28503 20893
rect 28537 20927 28595 20933
rect 28537 20893 28549 20927
rect 28583 20924 28595 20927
rect 28626 20924 28632 20936
rect 28583 20896 28632 20924
rect 28583 20893 28595 20896
rect 28537 20887 28595 20893
rect 27065 20859 27123 20865
rect 27065 20856 27077 20859
rect 23155 20828 26096 20856
rect 26160 20828 27077 20856
rect 23155 20825 23167 20828
rect 23109 20819 23167 20825
rect 13170 20788 13176 20800
rect 13131 20760 13176 20788
rect 13170 20748 13176 20760
rect 13228 20748 13234 20800
rect 19426 20748 19432 20800
rect 19484 20788 19490 20800
rect 19797 20791 19855 20797
rect 19797 20788 19809 20791
rect 19484 20760 19809 20788
rect 19484 20748 19490 20760
rect 19797 20757 19809 20760
rect 19843 20757 19855 20791
rect 19797 20751 19855 20757
rect 23198 20748 23204 20800
rect 23256 20788 23262 20800
rect 26160 20788 26188 20828
rect 27065 20825 27077 20828
rect 27111 20825 27123 20859
rect 27065 20819 27123 20825
rect 28460 20800 28488 20887
rect 28626 20884 28632 20896
rect 28684 20884 28690 20936
rect 28718 20884 28724 20936
rect 28776 20924 28782 20936
rect 28776 20896 28821 20924
rect 28776 20884 28782 20896
rect 30392 20856 30420 20952
rect 32674 20924 32680 20936
rect 32635 20896 32680 20924
rect 32674 20884 32680 20896
rect 32732 20884 32738 20936
rect 32858 20924 32864 20936
rect 32819 20896 32864 20924
rect 32858 20884 32864 20896
rect 32916 20884 32922 20936
rect 33686 20924 33692 20936
rect 33599 20896 33692 20924
rect 33686 20884 33692 20896
rect 33744 20924 33750 20936
rect 34146 20924 34152 20936
rect 33744 20896 34152 20924
rect 33744 20884 33750 20896
rect 34146 20884 34152 20896
rect 34204 20884 34210 20936
rect 37829 20927 37887 20933
rect 37829 20893 37841 20927
rect 37875 20893 37887 20927
rect 38102 20924 38108 20936
rect 38063 20896 38108 20924
rect 37829 20887 37887 20893
rect 31938 20856 31944 20868
rect 30392 20828 31944 20856
rect 31938 20816 31944 20828
rect 31996 20816 32002 20868
rect 32769 20859 32827 20865
rect 32769 20825 32781 20859
rect 32815 20856 32827 20859
rect 33870 20856 33876 20868
rect 32815 20828 33876 20856
rect 32815 20825 32827 20828
rect 32769 20819 32827 20825
rect 33870 20816 33876 20828
rect 33928 20816 33934 20868
rect 37844 20856 37872 20887
rect 38102 20884 38108 20896
rect 38160 20884 38166 20936
rect 38304 20933 38332 20964
rect 42613 20995 42671 21001
rect 42613 20961 42625 20995
rect 42659 20992 42671 20995
rect 42702 20992 42708 21004
rect 42659 20964 42708 20992
rect 42659 20961 42671 20964
rect 42613 20955 42671 20961
rect 42702 20952 42708 20964
rect 42760 20952 42766 21004
rect 44177 20995 44235 21001
rect 44177 20961 44189 20995
rect 44223 20992 44235 20995
rect 45462 20992 45468 21004
rect 44223 20964 45468 20992
rect 44223 20961 44235 20964
rect 44177 20955 44235 20961
rect 38289 20927 38347 20933
rect 38289 20893 38301 20927
rect 38335 20893 38347 20927
rect 40034 20924 40040 20936
rect 39995 20896 40040 20924
rect 38289 20887 38347 20893
rect 40034 20884 40040 20896
rect 40092 20884 40098 20936
rect 40310 20933 40316 20936
rect 40304 20924 40316 20933
rect 40271 20896 40316 20924
rect 40304 20887 40316 20896
rect 40310 20884 40316 20887
rect 40368 20884 40374 20936
rect 42429 20927 42487 20933
rect 42429 20893 42441 20927
rect 42475 20893 42487 20927
rect 42794 20924 42800 20936
rect 42707 20896 42800 20924
rect 42429 20887 42487 20893
rect 38746 20856 38752 20868
rect 37844 20828 38752 20856
rect 38304 20800 38332 20828
rect 38746 20816 38752 20828
rect 38804 20816 38810 20868
rect 23256 20760 26188 20788
rect 26421 20791 26479 20797
rect 23256 20748 23262 20760
rect 26421 20757 26433 20791
rect 26467 20788 26479 20791
rect 26694 20788 26700 20800
rect 26467 20760 26700 20788
rect 26467 20757 26479 20760
rect 26421 20751 26479 20757
rect 26694 20748 26700 20760
rect 26752 20748 26758 20800
rect 28442 20748 28448 20800
rect 28500 20748 28506 20800
rect 28626 20748 28632 20800
rect 28684 20788 28690 20800
rect 31202 20788 31208 20800
rect 28684 20760 31208 20788
rect 28684 20748 28690 20760
rect 31202 20748 31208 20760
rect 31260 20748 31266 20800
rect 37645 20791 37703 20797
rect 37645 20757 37657 20791
rect 37691 20788 37703 20791
rect 37918 20788 37924 20800
rect 37691 20760 37924 20788
rect 37691 20757 37703 20760
rect 37645 20751 37703 20757
rect 37918 20748 37924 20760
rect 37976 20748 37982 20800
rect 38286 20748 38292 20800
rect 38344 20748 38350 20800
rect 42444 20788 42472 20887
rect 42794 20884 42800 20896
rect 42852 20924 42858 20936
rect 42978 20924 42984 20936
rect 42852 20896 42984 20924
rect 42852 20884 42858 20896
rect 42978 20884 42984 20896
rect 43036 20884 43042 20936
rect 42521 20859 42579 20865
rect 42521 20825 42533 20859
rect 42567 20856 42579 20859
rect 43070 20856 43076 20868
rect 42567 20828 43076 20856
rect 42567 20825 42579 20828
rect 42521 20819 42579 20825
rect 43070 20816 43076 20828
rect 43128 20856 43134 20868
rect 43257 20859 43315 20865
rect 43257 20856 43269 20859
rect 43128 20828 43269 20856
rect 43128 20816 43134 20828
rect 43257 20825 43269 20828
rect 43303 20856 43315 20859
rect 44192 20856 44220 20955
rect 45462 20952 45468 20964
rect 45520 20952 45526 21004
rect 46492 21001 46520 21032
rect 47946 21020 47952 21032
rect 48004 21020 48010 21072
rect 46477 20995 46535 21001
rect 46477 20961 46489 20995
rect 46523 20961 46535 20995
rect 46658 20992 46664 21004
rect 46619 20964 46664 20992
rect 46477 20955 46535 20961
rect 46658 20952 46664 20964
rect 46716 20952 46722 21004
rect 48222 20992 48228 21004
rect 48183 20964 48228 20992
rect 48222 20952 48228 20964
rect 48280 20952 48286 21004
rect 44361 20927 44419 20933
rect 44361 20893 44373 20927
rect 44407 20924 44419 20927
rect 45922 20924 45928 20936
rect 44407 20896 45928 20924
rect 44407 20893 44419 20896
rect 44361 20887 44419 20893
rect 45922 20884 45928 20896
rect 45980 20884 45986 20936
rect 43303 20828 44220 20856
rect 43303 20825 43315 20828
rect 43257 20819 43315 20825
rect 43346 20788 43352 20800
rect 42444 20760 43352 20788
rect 43346 20748 43352 20760
rect 43404 20788 43410 20800
rect 43457 20791 43515 20797
rect 43457 20788 43469 20791
rect 43404 20760 43469 20788
rect 43404 20748 43410 20760
rect 43457 20757 43469 20760
rect 43503 20757 43515 20791
rect 43457 20751 43515 20757
rect 44266 20748 44272 20800
rect 44324 20788 44330 20800
rect 44545 20791 44603 20797
rect 44545 20788 44557 20791
rect 44324 20760 44557 20788
rect 44324 20748 44330 20760
rect 44545 20757 44557 20760
rect 44591 20757 44603 20791
rect 44545 20751 44603 20757
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 5074 20544 5080 20596
rect 5132 20584 5138 20596
rect 9582 20584 9588 20596
rect 5132 20556 9588 20584
rect 5132 20544 5138 20556
rect 9582 20544 9588 20556
rect 9640 20544 9646 20596
rect 12434 20584 12440 20596
rect 12395 20556 12440 20584
rect 12434 20544 12440 20556
rect 12492 20544 12498 20596
rect 15289 20587 15347 20593
rect 15289 20553 15301 20587
rect 15335 20584 15347 20587
rect 17862 20584 17868 20596
rect 15335 20556 17868 20584
rect 15335 20553 15347 20556
rect 15289 20547 15347 20553
rect 17862 20544 17868 20556
rect 17920 20544 17926 20596
rect 17954 20544 17960 20596
rect 18012 20584 18018 20596
rect 22094 20584 22100 20596
rect 18012 20556 22100 20584
rect 18012 20544 18018 20556
rect 22094 20544 22100 20556
rect 22152 20544 22158 20596
rect 23382 20544 23388 20596
rect 23440 20584 23446 20596
rect 24597 20587 24655 20593
rect 24597 20584 24609 20587
rect 23440 20556 24609 20584
rect 23440 20544 23446 20556
rect 24597 20553 24609 20556
rect 24643 20553 24655 20587
rect 24597 20547 24655 20553
rect 24765 20587 24823 20593
rect 24765 20553 24777 20587
rect 24811 20553 24823 20587
rect 24765 20547 24823 20553
rect 27157 20587 27215 20593
rect 27157 20553 27169 20587
rect 27203 20584 27215 20587
rect 27246 20584 27252 20596
rect 27203 20556 27252 20584
rect 27203 20553 27215 20556
rect 27157 20547 27215 20553
rect 13170 20476 13176 20528
rect 13228 20516 13234 20528
rect 13228 20488 19334 20516
rect 13228 20476 13234 20488
rect 4154 20448 4160 20460
rect 4115 20420 4160 20448
rect 4154 20408 4160 20420
rect 4212 20408 4218 20460
rect 10045 20451 10103 20457
rect 10045 20417 10057 20451
rect 10091 20448 10103 20451
rect 12526 20448 12532 20460
rect 10091 20420 12532 20448
rect 10091 20417 10103 20420
rect 10045 20411 10103 20417
rect 12526 20408 12532 20420
rect 12584 20408 12590 20460
rect 12621 20451 12679 20457
rect 12621 20417 12633 20451
rect 12667 20448 12679 20451
rect 13814 20448 13820 20460
rect 12667 20420 13820 20448
rect 12667 20417 12679 20420
rect 12621 20411 12679 20417
rect 13814 20408 13820 20420
rect 13872 20408 13878 20460
rect 18417 20451 18475 20457
rect 18417 20417 18429 20451
rect 18463 20448 18475 20451
rect 19058 20448 19064 20460
rect 18463 20420 19064 20448
rect 18463 20417 18475 20420
rect 18417 20411 18475 20417
rect 19058 20408 19064 20420
rect 19116 20408 19122 20460
rect 19306 20448 19334 20488
rect 19426 20476 19432 20528
rect 19484 20516 19490 20528
rect 19582 20519 19640 20525
rect 19582 20516 19594 20519
rect 19484 20488 19594 20516
rect 19484 20476 19490 20488
rect 19582 20485 19594 20488
rect 19628 20485 19640 20519
rect 24394 20516 24400 20528
rect 24355 20488 24400 20516
rect 19582 20479 19640 20485
rect 24394 20476 24400 20488
rect 24452 20476 24458 20528
rect 24780 20516 24808 20547
rect 27246 20544 27252 20556
rect 27304 20544 27310 20596
rect 29178 20584 29184 20596
rect 29091 20556 29184 20584
rect 29178 20544 29184 20556
rect 29236 20584 29242 20596
rect 29236 20556 29868 20584
rect 29236 20544 29242 20556
rect 25317 20519 25375 20525
rect 25317 20516 25329 20519
rect 24780 20488 25329 20516
rect 25317 20485 25329 20488
rect 25363 20485 25375 20519
rect 28353 20519 28411 20525
rect 28353 20516 28365 20519
rect 25317 20479 25375 20485
rect 27632 20488 28365 20516
rect 23382 20448 23388 20460
rect 19306 20420 20392 20448
rect 23343 20420 23388 20448
rect 4341 20383 4399 20389
rect 4341 20349 4353 20383
rect 4387 20380 4399 20383
rect 4890 20380 4896 20392
rect 4387 20352 4896 20380
rect 4387 20349 4399 20352
rect 4341 20343 4399 20349
rect 4890 20340 4896 20352
rect 4948 20340 4954 20392
rect 4985 20383 5043 20389
rect 4985 20349 4997 20383
rect 5031 20349 5043 20383
rect 10134 20380 10140 20392
rect 10095 20352 10140 20380
rect 4985 20343 5043 20349
rect 2958 20272 2964 20324
rect 3016 20312 3022 20324
rect 5000 20312 5028 20343
rect 10134 20340 10140 20352
rect 10192 20340 10198 20392
rect 10318 20340 10324 20392
rect 10376 20380 10382 20392
rect 10413 20383 10471 20389
rect 10413 20380 10425 20383
rect 10376 20352 10425 20380
rect 10376 20340 10382 20352
rect 10413 20349 10425 20352
rect 10459 20349 10471 20383
rect 10413 20343 10471 20349
rect 15286 20340 15292 20392
rect 15344 20380 15350 20392
rect 15381 20383 15439 20389
rect 15381 20380 15393 20383
rect 15344 20352 15393 20380
rect 15344 20340 15350 20352
rect 15381 20349 15393 20352
rect 15427 20349 15439 20383
rect 15381 20343 15439 20349
rect 15565 20383 15623 20389
rect 15565 20349 15577 20383
rect 15611 20380 15623 20383
rect 15838 20380 15844 20392
rect 15611 20352 15844 20380
rect 15611 20349 15623 20352
rect 15565 20343 15623 20349
rect 15838 20340 15844 20352
rect 15896 20340 15902 20392
rect 18138 20340 18144 20392
rect 18196 20380 18202 20392
rect 19337 20383 19395 20389
rect 19337 20380 19349 20383
rect 18196 20352 19349 20380
rect 18196 20340 18202 20352
rect 19337 20349 19349 20352
rect 19383 20349 19395 20383
rect 19337 20343 19395 20349
rect 3016 20284 5028 20312
rect 10152 20312 10180 20340
rect 20364 20312 20392 20420
rect 23382 20408 23388 20420
rect 23440 20408 23446 20460
rect 23474 20408 23480 20460
rect 23532 20448 23538 20460
rect 23661 20451 23719 20457
rect 23661 20448 23673 20451
rect 23532 20420 23673 20448
rect 23532 20408 23538 20420
rect 23661 20417 23673 20420
rect 23707 20417 23719 20451
rect 27338 20448 27344 20460
rect 27299 20420 27344 20448
rect 23661 20411 23719 20417
rect 27338 20408 27344 20420
rect 27396 20408 27402 20460
rect 27632 20457 27660 20488
rect 28353 20485 28365 20488
rect 28399 20516 28411 20519
rect 28534 20516 28540 20528
rect 28399 20488 28540 20516
rect 28399 20485 28411 20488
rect 28353 20479 28411 20485
rect 28534 20476 28540 20488
rect 28592 20516 28598 20528
rect 28592 20488 29224 20516
rect 28592 20476 28598 20488
rect 27617 20451 27675 20457
rect 27617 20417 27629 20451
rect 27663 20417 27675 20451
rect 27617 20411 27675 20417
rect 28169 20451 28227 20457
rect 28169 20417 28181 20451
rect 28215 20448 28227 20451
rect 28442 20448 28448 20460
rect 28215 20420 28448 20448
rect 28215 20417 28227 20420
rect 28169 20411 28227 20417
rect 28442 20408 28448 20420
rect 28500 20448 28506 20460
rect 28902 20448 28908 20460
rect 28500 20420 28908 20448
rect 28500 20408 28506 20420
rect 28902 20408 28908 20420
rect 28960 20448 28966 20460
rect 29196 20457 29224 20488
rect 29840 20457 29868 20556
rect 33134 20544 33140 20596
rect 33192 20584 33198 20596
rect 33781 20587 33839 20593
rect 33781 20584 33793 20587
rect 33192 20556 33793 20584
rect 33192 20544 33198 20556
rect 33781 20553 33793 20556
rect 33827 20553 33839 20587
rect 33781 20547 33839 20553
rect 35618 20544 35624 20596
rect 35676 20584 35682 20596
rect 41874 20584 41880 20596
rect 35676 20556 41880 20584
rect 35676 20544 35682 20556
rect 41874 20544 41880 20556
rect 41932 20544 41938 20596
rect 40034 20516 40040 20528
rect 37476 20488 40040 20516
rect 28997 20451 29055 20457
rect 28997 20448 29009 20451
rect 28960 20420 29009 20448
rect 28960 20408 28966 20420
rect 28997 20417 29009 20420
rect 29043 20417 29055 20451
rect 28997 20411 29055 20417
rect 29181 20451 29239 20457
rect 29181 20417 29193 20451
rect 29227 20417 29239 20451
rect 29181 20411 29239 20417
rect 29641 20451 29699 20457
rect 29641 20417 29653 20451
rect 29687 20417 29699 20451
rect 29641 20411 29699 20417
rect 29825 20451 29883 20457
rect 29825 20417 29837 20451
rect 29871 20417 29883 20451
rect 31018 20448 31024 20460
rect 30979 20420 31024 20448
rect 29825 20411 29883 20417
rect 23750 20380 23756 20392
rect 23711 20352 23756 20380
rect 23750 20340 23756 20352
rect 23808 20340 23814 20392
rect 28537 20383 28595 20389
rect 28537 20349 28549 20383
rect 28583 20380 28595 20383
rect 29656 20380 29684 20411
rect 31018 20408 31024 20420
rect 31076 20408 31082 20460
rect 31202 20408 31208 20460
rect 31260 20448 31266 20460
rect 31662 20448 31668 20460
rect 31260 20420 31668 20448
rect 31260 20408 31266 20420
rect 31662 20408 31668 20420
rect 31720 20408 31726 20460
rect 33686 20448 33692 20460
rect 33647 20420 33692 20448
rect 33686 20408 33692 20420
rect 33744 20408 33750 20460
rect 33870 20448 33876 20460
rect 33831 20420 33876 20448
rect 33870 20408 33876 20420
rect 33928 20408 33934 20460
rect 34333 20451 34391 20457
rect 34333 20417 34345 20451
rect 34379 20417 34391 20451
rect 34514 20448 34520 20460
rect 34475 20420 34520 20448
rect 34333 20411 34391 20417
rect 31294 20380 31300 20392
rect 28583 20352 29684 20380
rect 31255 20352 31300 20380
rect 28583 20349 28595 20352
rect 28537 20343 28595 20349
rect 31294 20340 31300 20352
rect 31352 20340 31358 20392
rect 34348 20380 34376 20411
rect 34514 20408 34520 20420
rect 34572 20408 34578 20460
rect 37476 20457 37504 20488
rect 40034 20476 40040 20488
rect 40092 20516 40098 20528
rect 40402 20516 40408 20528
rect 40092 20488 40408 20516
rect 40092 20476 40098 20488
rect 40402 20476 40408 20488
rect 40460 20476 40466 20528
rect 40494 20476 40500 20528
rect 40552 20516 40558 20528
rect 42702 20516 42708 20528
rect 40552 20488 42708 20516
rect 40552 20476 40558 20488
rect 42702 20476 42708 20488
rect 42760 20476 42766 20528
rect 37734 20457 37740 20460
rect 37461 20451 37519 20457
rect 37461 20417 37473 20451
rect 37507 20417 37519 20451
rect 37461 20411 37519 20417
rect 37728 20411 37740 20457
rect 37792 20448 37798 20460
rect 40310 20448 40316 20460
rect 37792 20420 37828 20448
rect 40271 20420 40316 20448
rect 37734 20408 37740 20411
rect 37792 20408 37798 20420
rect 40310 20408 40316 20420
rect 40368 20448 40374 20460
rect 40512 20448 40540 20476
rect 40368 20420 40540 20448
rect 40368 20408 40374 20420
rect 40586 20408 40592 20460
rect 40644 20448 40650 20460
rect 40773 20451 40831 20457
rect 40773 20448 40785 20451
rect 40644 20420 40785 20448
rect 40644 20408 40650 20420
rect 40773 20417 40785 20420
rect 40819 20417 40831 20451
rect 40773 20411 40831 20417
rect 46566 20408 46572 20460
rect 46624 20448 46630 20460
rect 46753 20451 46811 20457
rect 46753 20448 46765 20451
rect 46624 20420 46765 20448
rect 46624 20408 46630 20420
rect 46753 20417 46765 20420
rect 46799 20448 46811 20451
rect 46842 20448 46848 20460
rect 46799 20420 46848 20448
rect 46799 20417 46811 20420
rect 46753 20411 46811 20417
rect 46842 20408 46848 20420
rect 46900 20408 46906 20460
rect 34790 20380 34796 20392
rect 34348 20352 34796 20380
rect 34790 20340 34796 20352
rect 34848 20340 34854 20392
rect 39850 20340 39856 20392
rect 39908 20380 39914 20392
rect 40862 20380 40868 20392
rect 39908 20352 40868 20380
rect 39908 20340 39914 20352
rect 40862 20340 40868 20352
rect 40920 20340 40926 20392
rect 20622 20312 20628 20324
rect 10152 20284 19380 20312
rect 20364 20284 20628 20312
rect 3016 20272 3022 20284
rect 14921 20247 14979 20253
rect 14921 20213 14933 20247
rect 14967 20244 14979 20247
rect 15378 20244 15384 20256
rect 14967 20216 15384 20244
rect 14967 20213 14979 20216
rect 14921 20207 14979 20213
rect 15378 20204 15384 20216
rect 15436 20204 15442 20256
rect 18230 20244 18236 20256
rect 18191 20216 18236 20244
rect 18230 20204 18236 20216
rect 18288 20204 18294 20256
rect 19352 20244 19380 20284
rect 20622 20272 20628 20284
rect 20680 20312 20686 20324
rect 20717 20315 20775 20321
rect 20717 20312 20729 20315
rect 20680 20284 20729 20312
rect 20680 20272 20686 20284
rect 20717 20281 20729 20284
rect 20763 20281 20775 20315
rect 35618 20312 35624 20324
rect 20717 20275 20775 20281
rect 20824 20284 35624 20312
rect 20824 20244 20852 20284
rect 35618 20272 35624 20284
rect 35676 20272 35682 20324
rect 19352 20216 20852 20244
rect 23566 20204 23572 20256
rect 23624 20244 23630 20256
rect 24581 20247 24639 20253
rect 24581 20244 24593 20247
rect 23624 20216 24593 20244
rect 23624 20204 23630 20216
rect 24581 20213 24593 20216
rect 24627 20213 24639 20247
rect 24581 20207 24639 20213
rect 24854 20204 24860 20256
rect 24912 20244 24918 20256
rect 25409 20247 25467 20253
rect 25409 20244 25421 20247
rect 24912 20216 25421 20244
rect 24912 20204 24918 20216
rect 25409 20213 25421 20216
rect 25455 20213 25467 20247
rect 25409 20207 25467 20213
rect 26234 20204 26240 20256
rect 26292 20244 26298 20256
rect 27525 20247 27583 20253
rect 27525 20244 27537 20247
rect 26292 20216 27537 20244
rect 26292 20204 26298 20216
rect 27525 20213 27537 20216
rect 27571 20244 27583 20247
rect 28994 20244 29000 20256
rect 27571 20216 29000 20244
rect 27571 20213 27583 20216
rect 27525 20207 27583 20213
rect 28994 20204 29000 20216
rect 29052 20204 29058 20256
rect 29362 20204 29368 20256
rect 29420 20244 29426 20256
rect 29733 20247 29791 20253
rect 29733 20244 29745 20247
rect 29420 20216 29745 20244
rect 29420 20204 29426 20216
rect 29733 20213 29745 20216
rect 29779 20213 29791 20247
rect 29733 20207 29791 20213
rect 30837 20247 30895 20253
rect 30837 20213 30849 20247
rect 30883 20244 30895 20247
rect 30926 20244 30932 20256
rect 30883 20216 30932 20244
rect 30883 20213 30895 20216
rect 30837 20207 30895 20213
rect 30926 20204 30932 20216
rect 30984 20204 30990 20256
rect 33870 20204 33876 20256
rect 33928 20244 33934 20256
rect 34425 20247 34483 20253
rect 34425 20244 34437 20247
rect 33928 20216 34437 20244
rect 33928 20204 33934 20216
rect 34425 20213 34437 20216
rect 34471 20213 34483 20247
rect 34425 20207 34483 20213
rect 38194 20204 38200 20256
rect 38252 20244 38258 20256
rect 38841 20247 38899 20253
rect 38841 20244 38853 20247
rect 38252 20216 38853 20244
rect 38252 20204 38258 20216
rect 38841 20213 38853 20216
rect 38887 20213 38899 20247
rect 38841 20207 38899 20213
rect 46658 20204 46664 20256
rect 46716 20244 46722 20256
rect 46845 20247 46903 20253
rect 46845 20244 46857 20247
rect 46716 20216 46857 20244
rect 46716 20204 46722 20216
rect 46845 20213 46857 20216
rect 46891 20213 46903 20247
rect 47946 20244 47952 20256
rect 47907 20216 47952 20244
rect 46845 20207 46903 20213
rect 47946 20204 47952 20216
rect 48004 20204 48010 20256
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 4890 20040 4896 20052
rect 4851 20012 4896 20040
rect 4890 20000 4896 20012
rect 4948 20000 4954 20052
rect 15194 20040 15200 20052
rect 15155 20012 15200 20040
rect 15194 20000 15200 20012
rect 15252 20000 15258 20052
rect 17862 20000 17868 20052
rect 17920 20040 17926 20052
rect 20530 20040 20536 20052
rect 17920 20012 20536 20040
rect 17920 20000 17926 20012
rect 20530 20000 20536 20012
rect 20588 20000 20594 20052
rect 22557 20043 22615 20049
rect 22557 20009 22569 20043
rect 22603 20040 22615 20043
rect 23566 20040 23572 20052
rect 22603 20012 23572 20040
rect 22603 20009 22615 20012
rect 22557 20003 22615 20009
rect 23566 20000 23572 20012
rect 23624 20000 23630 20052
rect 28166 20000 28172 20052
rect 28224 20040 28230 20052
rect 28261 20043 28319 20049
rect 28261 20040 28273 20043
rect 28224 20012 28273 20040
rect 28224 20000 28230 20012
rect 28261 20009 28273 20012
rect 28307 20009 28319 20043
rect 28261 20003 28319 20009
rect 28994 20000 29000 20052
rect 29052 20040 29058 20052
rect 30098 20040 30104 20052
rect 29052 20012 30104 20040
rect 29052 20000 29058 20012
rect 30098 20000 30104 20012
rect 30156 20040 30162 20052
rect 32674 20040 32680 20052
rect 30156 20012 32680 20040
rect 30156 20000 30162 20012
rect 32674 20000 32680 20012
rect 32732 20000 32738 20052
rect 33686 20000 33692 20052
rect 33744 20040 33750 20052
rect 34146 20040 34152 20052
rect 33744 20012 34152 20040
rect 33744 20000 33750 20012
rect 34146 20000 34152 20012
rect 34204 20000 34210 20052
rect 34238 20000 34244 20052
rect 34296 20040 34302 20052
rect 35434 20040 35440 20052
rect 34296 20012 35440 20040
rect 34296 20000 34302 20012
rect 35434 20000 35440 20012
rect 35492 20040 35498 20052
rect 37734 20040 37740 20052
rect 35492 20012 36860 20040
rect 37695 20012 37740 20040
rect 35492 20000 35498 20012
rect 23382 19932 23388 19984
rect 23440 19932 23446 19984
rect 33962 19932 33968 19984
rect 34020 19932 34026 19984
rect 36832 19972 36860 20012
rect 37734 20000 37740 20012
rect 37792 20000 37798 20052
rect 40218 20000 40224 20052
rect 40276 20040 40282 20052
rect 40405 20043 40463 20049
rect 40405 20040 40417 20043
rect 40276 20012 40417 20040
rect 40276 20000 40282 20012
rect 40405 20009 40417 20012
rect 40451 20040 40463 20043
rect 40678 20040 40684 20052
rect 40451 20012 40684 20040
rect 40451 20009 40463 20012
rect 40405 20003 40463 20009
rect 40678 20000 40684 20012
rect 40736 20000 40742 20052
rect 39942 19972 39948 19984
rect 36832 19944 39948 19972
rect 39942 19932 39948 19944
rect 40000 19932 40006 19984
rect 47946 19972 47952 19984
rect 46492 19944 47952 19972
rect 10689 19907 10747 19913
rect 10689 19904 10701 19907
rect 6886 19876 10701 19904
rect 4798 19836 4804 19848
rect 4759 19808 4804 19836
rect 4798 19796 4804 19808
rect 4856 19836 4862 19848
rect 5534 19836 5540 19848
rect 4856 19808 5540 19836
rect 4856 19796 4862 19808
rect 5534 19796 5540 19808
rect 5592 19796 5598 19848
rect 198 19728 204 19780
rect 256 19768 262 19780
rect 6886 19768 6914 19876
rect 10689 19873 10701 19876
rect 10735 19873 10747 19907
rect 10689 19867 10747 19873
rect 18138 19864 18144 19916
rect 18196 19904 18202 19916
rect 18693 19907 18751 19913
rect 18693 19904 18705 19907
rect 18196 19876 18705 19904
rect 18196 19864 18202 19876
rect 18693 19873 18705 19876
rect 18739 19873 18751 19907
rect 18693 19867 18751 19873
rect 19334 19864 19340 19916
rect 19392 19904 19398 19916
rect 20809 19907 20867 19913
rect 20809 19904 20821 19907
rect 19392 19876 20821 19904
rect 19392 19864 19398 19876
rect 20809 19873 20821 19876
rect 20855 19873 20867 19907
rect 23400 19904 23428 19932
rect 30650 19904 30656 19916
rect 23400 19876 23612 19904
rect 30611 19876 30656 19904
rect 20809 19867 20867 19873
rect 9582 19836 9588 19848
rect 9543 19808 9588 19836
rect 9582 19796 9588 19808
rect 9640 19796 9646 19848
rect 10226 19836 10232 19848
rect 10187 19808 10232 19836
rect 10226 19796 10232 19808
rect 10284 19796 10290 19848
rect 15378 19836 15384 19848
rect 15339 19808 15384 19836
rect 15378 19796 15384 19808
rect 15436 19796 15442 19848
rect 15930 19796 15936 19848
rect 15988 19836 15994 19848
rect 16025 19839 16083 19845
rect 16025 19836 16037 19839
rect 15988 19808 16037 19836
rect 15988 19796 15994 19808
rect 16025 19805 16037 19808
rect 16071 19805 16083 19839
rect 17954 19836 17960 19848
rect 17915 19808 17960 19836
rect 16025 19799 16083 19805
rect 17954 19796 17960 19808
rect 18012 19796 18018 19848
rect 20622 19836 20628 19848
rect 20583 19808 20628 19836
rect 20622 19796 20628 19808
rect 20680 19796 20686 19848
rect 22370 19836 22376 19848
rect 22331 19808 22376 19836
rect 22370 19796 22376 19808
rect 22428 19796 22434 19848
rect 22646 19796 22652 19848
rect 22704 19836 22710 19848
rect 23385 19839 23443 19845
rect 22704 19808 22749 19836
rect 22704 19796 22710 19808
rect 23385 19805 23397 19839
rect 23431 19836 23443 19839
rect 23474 19836 23480 19848
rect 23431 19808 23480 19836
rect 23431 19805 23443 19808
rect 23385 19799 23443 19805
rect 23474 19796 23480 19808
rect 23532 19796 23538 19848
rect 23584 19845 23612 19876
rect 30650 19864 30656 19876
rect 30708 19864 30714 19916
rect 32950 19904 32956 19916
rect 31726 19876 32956 19904
rect 23569 19839 23627 19845
rect 23569 19805 23581 19839
rect 23615 19805 23627 19839
rect 27982 19836 27988 19848
rect 23569 19799 23627 19805
rect 23676 19808 27988 19836
rect 256 19740 6914 19768
rect 9677 19771 9735 19777
rect 256 19728 262 19740
rect 9677 19737 9689 19771
rect 9723 19768 9735 19771
rect 10413 19771 10471 19777
rect 10413 19768 10425 19771
rect 9723 19740 10425 19768
rect 9723 19737 9735 19740
rect 9677 19731 9735 19737
rect 10413 19737 10425 19740
rect 10459 19737 10471 19771
rect 10413 19731 10471 19737
rect 20717 19771 20775 19777
rect 20717 19737 20729 19771
rect 20763 19768 20775 19771
rect 23676 19768 23704 19808
rect 27982 19796 27988 19808
rect 28040 19796 28046 19848
rect 28442 19836 28448 19848
rect 28403 19808 28448 19836
rect 28442 19796 28448 19808
rect 28500 19796 28506 19848
rect 28718 19836 28724 19848
rect 28679 19808 28724 19836
rect 28718 19796 28724 19808
rect 28776 19796 28782 19848
rect 30926 19845 30932 19848
rect 30920 19836 30932 19845
rect 30887 19808 30932 19836
rect 30920 19799 30932 19808
rect 30926 19796 30932 19799
rect 30984 19796 30990 19848
rect 20763 19740 23704 19768
rect 23753 19771 23811 19777
rect 20763 19737 20775 19740
rect 20717 19731 20775 19737
rect 23753 19737 23765 19771
rect 23799 19768 23811 19771
rect 24673 19771 24731 19777
rect 24673 19768 24685 19771
rect 23799 19740 24685 19768
rect 23799 19737 23811 19740
rect 23753 19731 23811 19737
rect 24673 19737 24685 19740
rect 24719 19737 24731 19771
rect 24673 19731 24731 19737
rect 24857 19771 24915 19777
rect 24857 19737 24869 19771
rect 24903 19768 24915 19771
rect 25130 19768 25136 19780
rect 24903 19740 25136 19768
rect 24903 19737 24915 19740
rect 24857 19731 24915 19737
rect 25130 19728 25136 19740
rect 25188 19728 25194 19780
rect 28460 19768 28488 19796
rect 31726 19768 31754 19876
rect 32950 19864 32956 19876
rect 33008 19864 33014 19916
rect 33980 19904 34008 19932
rect 34241 19907 34299 19913
rect 34241 19904 34253 19907
rect 33980 19876 34253 19904
rect 34241 19873 34253 19876
rect 34287 19873 34299 19907
rect 34241 19867 34299 19873
rect 35161 19907 35219 19913
rect 35161 19873 35173 19907
rect 35207 19904 35219 19907
rect 35434 19904 35440 19916
rect 35207 19876 35440 19904
rect 35207 19873 35219 19876
rect 35161 19867 35219 19873
rect 35434 19864 35440 19876
rect 35492 19864 35498 19916
rect 38194 19904 38200 19916
rect 38155 19876 38200 19904
rect 38194 19864 38200 19876
rect 38252 19864 38258 19916
rect 32490 19836 32496 19848
rect 32403 19808 32496 19836
rect 32490 19796 32496 19808
rect 32548 19836 32554 19848
rect 32548 19808 32812 19836
rect 32548 19796 32554 19808
rect 28460 19740 31754 19768
rect 32677 19771 32735 19777
rect 32677 19737 32689 19771
rect 32723 19737 32735 19771
rect 32784 19768 32812 19808
rect 32858 19796 32864 19848
rect 32916 19836 32922 19848
rect 33965 19839 34023 19845
rect 33965 19836 33977 19839
rect 32916 19808 33977 19836
rect 32916 19796 32922 19808
rect 33965 19805 33977 19808
rect 34011 19836 34023 19839
rect 34514 19836 34520 19848
rect 34011 19808 34520 19836
rect 34011 19805 34023 19808
rect 33965 19799 34023 19805
rect 34514 19796 34520 19808
rect 34572 19796 34578 19848
rect 35069 19839 35127 19845
rect 35069 19805 35081 19839
rect 35115 19805 35127 19839
rect 35069 19799 35127 19805
rect 35897 19839 35955 19845
rect 35897 19805 35909 19839
rect 35943 19836 35955 19839
rect 37274 19836 37280 19848
rect 35943 19808 37280 19836
rect 35943 19805 35955 19808
rect 35897 19799 35955 19805
rect 33781 19771 33839 19777
rect 32784 19740 33732 19768
rect 32677 19731 32735 19737
rect 15470 19660 15476 19712
rect 15528 19700 15534 19712
rect 15841 19703 15899 19709
rect 15841 19700 15853 19703
rect 15528 19672 15853 19700
rect 15528 19660 15534 19672
rect 15841 19669 15853 19672
rect 15887 19669 15899 19703
rect 15841 19663 15899 19669
rect 20070 19660 20076 19712
rect 20128 19700 20134 19712
rect 20257 19703 20315 19709
rect 20257 19700 20269 19703
rect 20128 19672 20269 19700
rect 20128 19660 20134 19672
rect 20257 19669 20269 19672
rect 20303 19669 20315 19703
rect 22186 19700 22192 19712
rect 22147 19672 22192 19700
rect 20257 19663 20315 19669
rect 22186 19660 22192 19672
rect 22244 19660 22250 19712
rect 28629 19703 28687 19709
rect 28629 19669 28641 19703
rect 28675 19700 28687 19703
rect 29454 19700 29460 19712
rect 28675 19672 29460 19700
rect 28675 19669 28687 19672
rect 28629 19663 28687 19669
rect 29454 19660 29460 19672
rect 29512 19660 29518 19712
rect 32030 19700 32036 19712
rect 31943 19672 32036 19700
rect 32030 19660 32036 19672
rect 32088 19700 32094 19712
rect 32692 19700 32720 19731
rect 32858 19700 32864 19712
rect 32088 19672 32720 19700
rect 32819 19672 32864 19700
rect 32088 19660 32094 19672
rect 32858 19660 32864 19672
rect 32916 19660 32922 19712
rect 33704 19700 33732 19740
rect 33781 19737 33793 19771
rect 33827 19768 33839 19771
rect 35084 19768 35112 19799
rect 37274 19796 37280 19808
rect 37332 19796 37338 19848
rect 37918 19836 37924 19848
rect 37879 19808 37924 19836
rect 37918 19796 37924 19808
rect 37976 19796 37982 19848
rect 38105 19839 38163 19845
rect 38105 19805 38117 19839
rect 38151 19805 38163 19839
rect 39960 19836 39988 19932
rect 40402 19864 40408 19916
rect 40460 19904 40466 19916
rect 41877 19907 41935 19913
rect 41877 19904 41889 19907
rect 40460 19876 41889 19904
rect 40460 19864 40466 19876
rect 41877 19873 41889 19876
rect 41923 19873 41935 19907
rect 41877 19867 41935 19873
rect 44177 19907 44235 19913
rect 44177 19873 44189 19907
rect 44223 19904 44235 19907
rect 44450 19904 44456 19916
rect 44223 19876 44456 19904
rect 44223 19873 44235 19876
rect 44177 19867 44235 19873
rect 44450 19864 44456 19876
rect 44508 19864 44514 19916
rect 46492 19913 46520 19944
rect 47946 19932 47952 19944
rect 48004 19932 48010 19984
rect 46477 19907 46535 19913
rect 46477 19873 46489 19907
rect 46523 19873 46535 19907
rect 46658 19904 46664 19916
rect 46619 19876 46664 19904
rect 46477 19867 46535 19873
rect 46658 19864 46664 19876
rect 46716 19864 46722 19916
rect 48222 19904 48228 19916
rect 48183 19876 48228 19904
rect 48222 19864 48228 19876
rect 48280 19864 48286 19916
rect 40129 19839 40187 19845
rect 40129 19836 40141 19839
rect 39960 19808 40141 19836
rect 38105 19799 38163 19805
rect 40129 19805 40141 19808
rect 40175 19805 40187 19839
rect 42150 19836 42156 19848
rect 42111 19808 42156 19836
rect 40129 19799 40187 19805
rect 35618 19768 35624 19780
rect 33827 19740 35624 19768
rect 33827 19737 33839 19740
rect 33781 19731 33839 19737
rect 35618 19728 35624 19740
rect 35676 19728 35682 19780
rect 35986 19728 35992 19780
rect 36044 19768 36050 19780
rect 36142 19771 36200 19777
rect 36142 19768 36154 19771
rect 36044 19740 36154 19768
rect 36044 19728 36050 19740
rect 36142 19737 36154 19740
rect 36188 19737 36200 19771
rect 38120 19768 38148 19799
rect 42150 19796 42156 19808
rect 42208 19796 42214 19848
rect 43993 19839 44051 19845
rect 43993 19805 44005 19839
rect 44039 19836 44051 19839
rect 44266 19836 44272 19848
rect 44039 19808 44272 19836
rect 44039 19805 44051 19808
rect 43993 19799 44051 19805
rect 44266 19796 44272 19808
rect 44324 19796 44330 19848
rect 44361 19839 44419 19845
rect 44361 19805 44373 19839
rect 44407 19836 44419 19839
rect 44542 19836 44548 19848
rect 44407 19808 44548 19836
rect 44407 19805 44419 19808
rect 44361 19799 44419 19805
rect 44542 19796 44548 19808
rect 44600 19796 44606 19848
rect 38378 19768 38384 19780
rect 36142 19731 36200 19737
rect 37200 19740 38384 19768
rect 34238 19700 34244 19712
rect 33704 19672 34244 19700
rect 34238 19660 34244 19672
rect 34296 19660 34302 19712
rect 35342 19660 35348 19712
rect 35400 19700 35406 19712
rect 35437 19703 35495 19709
rect 35437 19700 35449 19703
rect 35400 19672 35449 19700
rect 35400 19660 35406 19672
rect 35437 19669 35449 19672
rect 35483 19669 35495 19703
rect 35437 19663 35495 19669
rect 35710 19660 35716 19712
rect 35768 19700 35774 19712
rect 37200 19700 37228 19740
rect 38378 19728 38384 19740
rect 38436 19768 38442 19780
rect 39022 19768 39028 19780
rect 38436 19740 39028 19768
rect 38436 19728 38442 19740
rect 39022 19728 39028 19740
rect 39080 19728 39086 19780
rect 43438 19728 43444 19780
rect 43496 19768 43502 19780
rect 44085 19771 44143 19777
rect 44085 19768 44097 19771
rect 43496 19740 44097 19768
rect 43496 19728 43502 19740
rect 44085 19737 44097 19740
rect 44131 19737 44143 19771
rect 44085 19731 44143 19737
rect 35768 19672 37228 19700
rect 37277 19703 37335 19709
rect 35768 19660 35774 19672
rect 37277 19669 37289 19703
rect 37323 19700 37335 19703
rect 37458 19700 37464 19712
rect 37323 19672 37464 19700
rect 37323 19669 37335 19672
rect 37277 19663 37335 19669
rect 37458 19660 37464 19672
rect 37516 19660 37522 19712
rect 41874 19660 41880 19712
rect 41932 19700 41938 19712
rect 43257 19703 43315 19709
rect 43257 19700 43269 19703
rect 41932 19672 43269 19700
rect 41932 19660 41938 19672
rect 43257 19669 43269 19672
rect 43303 19700 43315 19703
rect 43346 19700 43352 19712
rect 43303 19672 43352 19700
rect 43303 19669 43315 19672
rect 43257 19663 43315 19669
rect 43346 19660 43352 19672
rect 43404 19660 43410 19712
rect 44174 19660 44180 19712
rect 44232 19700 44238 19712
rect 44269 19703 44327 19709
rect 44269 19700 44281 19703
rect 44232 19672 44281 19700
rect 44232 19660 44238 19672
rect 44269 19669 44281 19672
rect 44315 19669 44327 19703
rect 44269 19663 44327 19669
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 12526 19456 12532 19508
rect 12584 19496 12590 19508
rect 13081 19499 13139 19505
rect 13081 19496 13093 19499
rect 12584 19468 13093 19496
rect 12584 19456 12590 19468
rect 13081 19465 13093 19468
rect 13127 19465 13139 19499
rect 13081 19459 13139 19465
rect 18233 19499 18291 19505
rect 18233 19465 18245 19499
rect 18279 19496 18291 19499
rect 19058 19496 19064 19508
rect 18279 19468 18736 19496
rect 19019 19468 19064 19496
rect 18279 19465 18291 19468
rect 18233 19459 18291 19465
rect 18708 19437 18736 19468
rect 19058 19456 19064 19468
rect 19116 19456 19122 19508
rect 19978 19456 19984 19508
rect 20036 19496 20042 19508
rect 20165 19499 20223 19505
rect 20165 19496 20177 19499
rect 20036 19468 20177 19496
rect 20036 19456 20042 19468
rect 20165 19465 20177 19468
rect 20211 19465 20223 19499
rect 20165 19459 20223 19465
rect 26418 19456 26424 19508
rect 26476 19496 26482 19508
rect 28077 19499 28135 19505
rect 28077 19496 28089 19499
rect 26476 19468 28089 19496
rect 26476 19456 26482 19468
rect 28077 19465 28089 19468
rect 28123 19465 28135 19499
rect 28077 19459 28135 19465
rect 28718 19456 28724 19508
rect 28776 19496 28782 19508
rect 28905 19499 28963 19505
rect 28905 19496 28917 19499
rect 28776 19468 28917 19496
rect 28776 19456 28782 19468
rect 28905 19465 28917 19468
rect 28951 19465 28963 19499
rect 29454 19496 29460 19508
rect 29415 19468 29460 19496
rect 28905 19459 28963 19465
rect 29454 19456 29460 19468
rect 29512 19456 29518 19508
rect 31018 19496 31024 19508
rect 30979 19468 31024 19496
rect 31018 19456 31024 19468
rect 31076 19456 31082 19508
rect 32674 19456 32680 19508
rect 32732 19496 32738 19508
rect 35710 19496 35716 19508
rect 32732 19468 35716 19496
rect 32732 19456 32738 19468
rect 35710 19456 35716 19468
rect 35768 19456 35774 19508
rect 35897 19499 35955 19505
rect 35897 19465 35909 19499
rect 35943 19496 35955 19499
rect 35986 19496 35992 19508
rect 35943 19468 35992 19496
rect 35943 19465 35955 19468
rect 35897 19459 35955 19465
rect 35986 19456 35992 19468
rect 36044 19456 36050 19508
rect 36541 19499 36599 19505
rect 36541 19496 36553 19499
rect 36096 19468 36553 19496
rect 17773 19431 17831 19437
rect 17773 19428 17785 19431
rect 17604 19400 17785 19428
rect 9950 19360 9956 19372
rect 9911 19332 9956 19360
rect 9950 19320 9956 19332
rect 10008 19320 10014 19372
rect 11514 19320 11520 19372
rect 11572 19360 11578 19372
rect 11701 19363 11759 19369
rect 11701 19360 11713 19363
rect 11572 19332 11713 19360
rect 11572 19320 11578 19332
rect 11701 19329 11713 19332
rect 11747 19329 11759 19363
rect 11701 19323 11759 19329
rect 11790 19320 11796 19372
rect 11848 19360 11854 19372
rect 11957 19363 12015 19369
rect 11957 19360 11969 19363
rect 11848 19332 11969 19360
rect 11848 19320 11854 19332
rect 11957 19329 11969 19332
rect 12003 19329 12015 19363
rect 13906 19360 13912 19372
rect 13867 19332 13912 19360
rect 11957 19323 12015 19329
rect 13906 19320 13912 19332
rect 13964 19320 13970 19372
rect 14918 19360 14924 19372
rect 14879 19332 14924 19360
rect 14918 19320 14924 19332
rect 14976 19320 14982 19372
rect 10042 19292 10048 19304
rect 10003 19264 10048 19292
rect 10042 19252 10048 19264
rect 10100 19252 10106 19304
rect 10226 19252 10232 19304
rect 10284 19292 10290 19304
rect 10321 19295 10379 19301
rect 10321 19292 10333 19295
rect 10284 19264 10333 19292
rect 10284 19252 10290 19264
rect 10321 19261 10333 19264
rect 10367 19261 10379 19295
rect 10321 19255 10379 19261
rect 14001 19295 14059 19301
rect 14001 19261 14013 19295
rect 14047 19261 14059 19295
rect 14001 19255 14059 19261
rect 14016 19224 14044 19255
rect 14090 19252 14096 19304
rect 14148 19292 14154 19304
rect 14829 19295 14887 19301
rect 14829 19292 14841 19295
rect 14148 19264 14841 19292
rect 14148 19252 14154 19264
rect 14829 19261 14841 19264
rect 14875 19261 14887 19295
rect 14829 19255 14887 19261
rect 15010 19252 15016 19304
rect 15068 19292 15074 19304
rect 15068 19264 16574 19292
rect 15068 19252 15074 19264
rect 15289 19227 15347 19233
rect 15289 19224 15301 19227
rect 14016 19196 15301 19224
rect 15289 19193 15301 19196
rect 15335 19193 15347 19227
rect 16546 19224 16574 19264
rect 17221 19227 17279 19233
rect 17221 19224 17233 19227
rect 16546 19196 17233 19224
rect 15289 19187 15347 19193
rect 17221 19193 17233 19196
rect 17267 19193 17279 19227
rect 17221 19187 17279 19193
rect 14185 19159 14243 19165
rect 14185 19125 14197 19159
rect 14231 19156 14243 19159
rect 15194 19156 15200 19168
rect 14231 19128 15200 19156
rect 14231 19125 14243 19128
rect 14185 19119 14243 19125
rect 15194 19116 15200 19128
rect 15252 19116 15258 19168
rect 17236 19156 17264 19187
rect 17604 19156 17632 19400
rect 17773 19397 17785 19400
rect 17819 19397 17831 19431
rect 17773 19391 17831 19397
rect 18693 19431 18751 19437
rect 18693 19397 18705 19431
rect 18739 19397 18751 19431
rect 18874 19428 18880 19440
rect 18835 19400 18880 19428
rect 18693 19391 18751 19397
rect 18874 19388 18880 19400
rect 18932 19388 18938 19440
rect 19705 19431 19763 19437
rect 19705 19397 19717 19431
rect 19751 19428 19763 19431
rect 20254 19428 20260 19440
rect 19751 19400 20260 19428
rect 19751 19397 19763 19400
rect 19705 19391 19763 19397
rect 20254 19388 20260 19400
rect 20312 19388 20318 19440
rect 22741 19431 22799 19437
rect 22741 19397 22753 19431
rect 22787 19428 22799 19431
rect 24762 19428 24768 19440
rect 22787 19400 24768 19428
rect 22787 19397 22799 19400
rect 22741 19391 22799 19397
rect 24762 19388 24768 19400
rect 24820 19388 24826 19440
rect 30282 19428 30288 19440
rect 25240 19400 30288 19428
rect 17862 19360 17868 19372
rect 17823 19332 17868 19360
rect 17862 19320 17868 19332
rect 17920 19320 17926 19372
rect 22922 19360 22928 19372
rect 22883 19332 22928 19360
rect 22922 19320 22928 19332
rect 22980 19320 22986 19372
rect 23106 19320 23112 19372
rect 23164 19360 23170 19372
rect 23201 19363 23259 19369
rect 23201 19360 23213 19363
rect 23164 19332 23213 19360
rect 23164 19320 23170 19332
rect 23201 19329 23213 19332
rect 23247 19329 23259 19363
rect 23201 19323 23259 19329
rect 23385 19363 23443 19369
rect 23385 19329 23397 19363
rect 23431 19329 23443 19363
rect 23385 19323 23443 19329
rect 24397 19363 24455 19369
rect 24397 19329 24409 19363
rect 24443 19360 24455 19363
rect 24854 19360 24860 19372
rect 24443 19332 24860 19360
rect 24443 19329 24455 19332
rect 24397 19323 24455 19329
rect 17681 19295 17739 19301
rect 17681 19261 17693 19295
rect 17727 19292 17739 19295
rect 19334 19292 19340 19304
rect 17727 19264 19340 19292
rect 17727 19261 17739 19264
rect 17681 19255 17739 19261
rect 19334 19252 19340 19264
rect 19392 19252 19398 19304
rect 22646 19252 22652 19304
rect 22704 19292 22710 19304
rect 23400 19292 23428 19323
rect 24854 19320 24860 19332
rect 24912 19320 24918 19372
rect 25240 19369 25268 19400
rect 30282 19388 30288 19400
rect 30340 19388 30346 19440
rect 32858 19388 32864 19440
rect 32916 19428 32922 19440
rect 35526 19428 35532 19440
rect 32916 19400 35204 19428
rect 32916 19388 32922 19400
rect 25225 19363 25283 19369
rect 25225 19329 25237 19363
rect 25271 19329 25283 19363
rect 25225 19323 25283 19329
rect 25492 19363 25550 19369
rect 25492 19329 25504 19363
rect 25538 19360 25550 19363
rect 26786 19360 26792 19372
rect 25538 19332 26792 19360
rect 25538 19329 25550 19332
rect 25492 19323 25550 19329
rect 26786 19320 26792 19332
rect 26844 19320 26850 19372
rect 27157 19363 27215 19369
rect 27157 19329 27169 19363
rect 27203 19329 27215 19363
rect 27338 19360 27344 19372
rect 27299 19332 27344 19360
rect 27157 19323 27215 19329
rect 22704 19264 23428 19292
rect 22704 19252 22710 19264
rect 20070 19224 20076 19236
rect 20031 19196 20076 19224
rect 20070 19184 20076 19196
rect 20128 19184 20134 19236
rect 20180 19196 25268 19224
rect 20180 19156 20208 19196
rect 17236 19128 20208 19156
rect 22462 19116 22468 19168
rect 22520 19156 22526 19168
rect 23750 19156 23756 19168
rect 22520 19128 23756 19156
rect 22520 19116 22526 19128
rect 23750 19116 23756 19128
rect 23808 19116 23814 19168
rect 24670 19156 24676 19168
rect 24631 19128 24676 19156
rect 24670 19116 24676 19128
rect 24728 19116 24734 19168
rect 25240 19156 25268 19196
rect 26326 19184 26332 19236
rect 26384 19224 26390 19236
rect 26605 19227 26663 19233
rect 26605 19224 26617 19227
rect 26384 19196 26617 19224
rect 26384 19184 26390 19196
rect 26605 19193 26617 19196
rect 26651 19224 26663 19227
rect 27172 19224 27200 19323
rect 27338 19320 27344 19332
rect 27396 19320 27402 19372
rect 27801 19363 27859 19369
rect 27801 19329 27813 19363
rect 27847 19360 27859 19363
rect 28258 19360 28264 19372
rect 27847 19332 28264 19360
rect 27847 19329 27859 19332
rect 27801 19323 27859 19329
rect 28258 19320 28264 19332
rect 28316 19320 28322 19372
rect 28537 19363 28595 19369
rect 28537 19329 28549 19363
rect 28583 19329 28595 19363
rect 28718 19360 28724 19372
rect 28679 19332 28724 19360
rect 28537 19323 28595 19329
rect 28074 19292 28080 19304
rect 28035 19264 28080 19292
rect 28074 19252 28080 19264
rect 28132 19252 28138 19304
rect 28552 19292 28580 19323
rect 28718 19320 28724 19332
rect 28776 19320 28782 19372
rect 29362 19360 29368 19372
rect 28828 19332 29368 19360
rect 28626 19292 28632 19304
rect 28539 19264 28632 19292
rect 28626 19252 28632 19264
rect 28684 19292 28690 19304
rect 28828 19292 28856 19332
rect 29362 19320 29368 19332
rect 29420 19320 29426 19372
rect 29549 19363 29607 19369
rect 29549 19329 29561 19363
rect 29595 19329 29607 19363
rect 29549 19323 29607 19329
rect 28684 19264 28856 19292
rect 29564 19292 29592 19323
rect 29914 19320 29920 19372
rect 29972 19360 29978 19372
rect 31018 19360 31024 19372
rect 29972 19332 31024 19360
rect 29972 19320 29978 19332
rect 31018 19320 31024 19332
rect 31076 19360 31082 19372
rect 31205 19363 31263 19369
rect 31205 19360 31217 19363
rect 31076 19332 31217 19360
rect 31076 19320 31082 19332
rect 31205 19329 31217 19332
rect 31251 19329 31263 19363
rect 31478 19360 31484 19372
rect 31439 19332 31484 19360
rect 31205 19323 31263 19329
rect 31478 19320 31484 19332
rect 31536 19320 31542 19372
rect 31665 19363 31723 19369
rect 31665 19329 31677 19363
rect 31711 19360 31723 19363
rect 32030 19360 32036 19372
rect 31711 19332 32036 19360
rect 31711 19329 31723 19332
rect 31665 19323 31723 19329
rect 32030 19320 32036 19332
rect 32088 19320 32094 19372
rect 33686 19320 33692 19372
rect 33744 19360 33750 19372
rect 33873 19363 33931 19369
rect 33873 19360 33885 19363
rect 33744 19332 33885 19360
rect 33744 19320 33750 19332
rect 33873 19329 33885 19332
rect 33919 19329 33931 19363
rect 33873 19323 33931 19329
rect 33962 19320 33968 19372
rect 34020 19360 34026 19372
rect 35176 19369 35204 19400
rect 35452 19400 35532 19428
rect 34241 19363 34299 19369
rect 34241 19360 34253 19363
rect 34020 19332 34253 19360
rect 34020 19320 34026 19332
rect 34241 19329 34253 19332
rect 34287 19329 34299 19363
rect 34241 19323 34299 19329
rect 35161 19363 35219 19369
rect 35161 19329 35173 19363
rect 35207 19329 35219 19363
rect 35342 19360 35348 19372
rect 35303 19332 35348 19360
rect 35161 19323 35219 19329
rect 35342 19320 35348 19332
rect 35400 19320 35406 19372
rect 31570 19292 31576 19304
rect 29564 19264 31576 19292
rect 28684 19252 28690 19264
rect 26651 19196 27200 19224
rect 26651 19193 26663 19196
rect 26605 19187 26663 19193
rect 27706 19184 27712 19236
rect 27764 19224 27770 19236
rect 28718 19224 28724 19236
rect 27764 19196 28724 19224
rect 27764 19184 27770 19196
rect 28718 19184 28724 19196
rect 28776 19224 28782 19236
rect 29564 19224 29592 19264
rect 31570 19252 31576 19264
rect 31628 19252 31634 19304
rect 33781 19295 33839 19301
rect 33781 19261 33793 19295
rect 33827 19292 33839 19295
rect 35250 19292 35256 19304
rect 33827 19264 35256 19292
rect 33827 19261 33839 19264
rect 33781 19255 33839 19261
rect 35250 19252 35256 19264
rect 35308 19252 35314 19304
rect 35452 19301 35480 19400
rect 35526 19388 35532 19400
rect 35584 19388 35590 19440
rect 35802 19388 35808 19440
rect 35860 19428 35866 19440
rect 36096 19428 36124 19468
rect 36541 19465 36553 19468
rect 36587 19465 36599 19499
rect 40126 19496 40132 19508
rect 40087 19468 40132 19496
rect 36541 19459 36599 19465
rect 40126 19456 40132 19468
rect 40184 19456 40190 19508
rect 43530 19496 43536 19508
rect 43491 19468 43536 19496
rect 43530 19456 43536 19468
rect 43588 19456 43594 19508
rect 43806 19496 43812 19508
rect 43719 19468 43812 19496
rect 37458 19428 37464 19440
rect 35860 19400 36124 19428
rect 36464 19400 37464 19428
rect 35860 19388 35866 19400
rect 36464 19369 36492 19400
rect 37458 19388 37464 19400
rect 37516 19388 37522 19440
rect 37645 19431 37703 19437
rect 37645 19397 37657 19431
rect 37691 19428 37703 19431
rect 38194 19428 38200 19440
rect 37691 19400 38200 19428
rect 37691 19397 37703 19400
rect 37645 19391 37703 19397
rect 35713 19363 35771 19369
rect 35713 19329 35725 19363
rect 35759 19360 35771 19363
rect 36449 19363 36507 19369
rect 36449 19360 36461 19363
rect 35759 19332 36461 19360
rect 35759 19329 35771 19332
rect 35713 19323 35771 19329
rect 36449 19329 36461 19332
rect 36495 19329 36507 19363
rect 36449 19323 36507 19329
rect 36633 19363 36691 19369
rect 36633 19329 36645 19363
rect 36679 19360 36691 19363
rect 37660 19360 37688 19391
rect 38194 19388 38200 19400
rect 38252 19388 38258 19440
rect 43438 19388 43444 19440
rect 43496 19428 43502 19440
rect 43732 19437 43760 19468
rect 43806 19456 43812 19468
rect 43864 19496 43870 19508
rect 44637 19499 44695 19505
rect 44637 19496 44649 19499
rect 43864 19468 44649 19496
rect 43864 19456 43870 19468
rect 44637 19465 44649 19468
rect 44683 19465 44695 19499
rect 44637 19459 44695 19465
rect 43717 19431 43775 19437
rect 43717 19428 43729 19431
rect 43496 19400 43729 19428
rect 43496 19388 43502 19400
rect 43717 19397 43729 19400
rect 43763 19397 43775 19431
rect 44266 19428 44272 19440
rect 43717 19391 43775 19397
rect 43824 19400 44272 19428
rect 39942 19360 39948 19372
rect 36679 19332 37688 19360
rect 39903 19332 39948 19360
rect 36679 19329 36691 19332
rect 36633 19323 36691 19329
rect 39942 19320 39948 19332
rect 40000 19320 40006 19372
rect 41874 19360 41880 19372
rect 41835 19332 41880 19360
rect 41874 19320 41880 19332
rect 41932 19320 41938 19372
rect 41969 19363 42027 19369
rect 41969 19329 41981 19363
rect 42015 19360 42027 19363
rect 42794 19360 42800 19372
rect 42015 19332 42800 19360
rect 42015 19329 42027 19332
rect 41969 19323 42027 19329
rect 42794 19320 42800 19332
rect 42852 19320 42858 19372
rect 43346 19360 43352 19372
rect 43307 19332 43352 19360
rect 43346 19320 43352 19332
rect 43404 19320 43410 19372
rect 43824 19369 43852 19400
rect 44266 19388 44272 19400
rect 44324 19428 44330 19440
rect 44324 19400 44772 19428
rect 44324 19388 44330 19400
rect 43809 19363 43867 19369
rect 43809 19329 43821 19363
rect 43855 19329 43867 19363
rect 44450 19360 44456 19372
rect 44363 19332 44456 19360
rect 43809 19323 43867 19329
rect 44450 19320 44456 19332
rect 44508 19320 44514 19372
rect 44744 19369 44772 19400
rect 44729 19363 44787 19369
rect 44729 19329 44741 19363
rect 44775 19329 44787 19363
rect 44729 19323 44787 19329
rect 47029 19363 47087 19369
rect 47029 19329 47041 19363
rect 47075 19360 47087 19363
rect 47302 19360 47308 19372
rect 47075 19332 47308 19360
rect 47075 19329 47087 19332
rect 47029 19323 47087 19329
rect 47302 19320 47308 19332
rect 47360 19320 47366 19372
rect 35437 19295 35495 19301
rect 35437 19261 35449 19295
rect 35483 19261 35495 19295
rect 35437 19255 35495 19261
rect 35529 19295 35587 19301
rect 35529 19261 35541 19295
rect 35575 19292 35587 19295
rect 35894 19292 35900 19304
rect 35575 19264 35900 19292
rect 35575 19261 35587 19264
rect 35529 19255 35587 19261
rect 35894 19252 35900 19264
rect 35952 19252 35958 19304
rect 39482 19252 39488 19304
rect 39540 19292 39546 19304
rect 39761 19295 39819 19301
rect 39761 19292 39773 19295
rect 39540 19264 39773 19292
rect 39540 19252 39546 19264
rect 39761 19261 39773 19264
rect 39807 19292 39819 19295
rect 40310 19292 40316 19304
rect 39807 19264 40316 19292
rect 39807 19261 39819 19264
rect 39761 19255 39819 19261
rect 40310 19252 40316 19264
rect 40368 19252 40374 19304
rect 43441 19295 43499 19301
rect 43441 19261 43453 19295
rect 43487 19292 43499 19295
rect 44468 19292 44496 19320
rect 43487 19264 44496 19292
rect 43487 19261 43499 19264
rect 43441 19255 43499 19261
rect 28776 19196 29592 19224
rect 28776 19184 28782 19196
rect 33594 19184 33600 19236
rect 33652 19224 33658 19236
rect 43456 19224 43484 19255
rect 33652 19196 43484 19224
rect 33652 19184 33658 19196
rect 27062 19156 27068 19168
rect 25240 19128 27068 19156
rect 27062 19116 27068 19128
rect 27120 19116 27126 19168
rect 27157 19159 27215 19165
rect 27157 19125 27169 19159
rect 27203 19156 27215 19159
rect 27522 19156 27528 19168
rect 27203 19128 27528 19156
rect 27203 19125 27215 19128
rect 27157 19119 27215 19125
rect 27522 19116 27528 19128
rect 27580 19116 27586 19168
rect 27893 19159 27951 19165
rect 27893 19125 27905 19159
rect 27939 19156 27951 19159
rect 28994 19156 29000 19168
rect 27939 19128 29000 19156
rect 27939 19125 27951 19128
rect 27893 19119 27951 19125
rect 28994 19116 29000 19128
rect 29052 19116 29058 19168
rect 34146 19156 34152 19168
rect 34107 19128 34152 19156
rect 34146 19116 34152 19128
rect 34204 19116 34210 19168
rect 34422 19156 34428 19168
rect 34383 19128 34428 19156
rect 34422 19116 34428 19128
rect 34480 19116 34486 19168
rect 36630 19116 36636 19168
rect 36688 19156 36694 19168
rect 37829 19159 37887 19165
rect 37829 19156 37841 19159
rect 36688 19128 37841 19156
rect 36688 19116 36694 19128
rect 37829 19125 37841 19128
rect 37875 19125 37887 19159
rect 37829 19119 37887 19125
rect 43070 19116 43076 19168
rect 43128 19156 43134 19168
rect 43165 19159 43223 19165
rect 43165 19156 43177 19159
rect 43128 19128 43177 19156
rect 43128 19116 43134 19128
rect 43165 19125 43177 19128
rect 43211 19125 43223 19159
rect 44266 19156 44272 19168
rect 44227 19128 44272 19156
rect 43165 19119 43223 19125
rect 44266 19116 44272 19128
rect 44324 19116 44330 19168
rect 47118 19156 47124 19168
rect 47079 19128 47124 19156
rect 47118 19116 47124 19128
rect 47176 19116 47182 19168
rect 47946 19156 47952 19168
rect 47907 19128 47952 19156
rect 47946 19116 47952 19128
rect 48004 19116 48010 19168
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 11701 18955 11759 18961
rect 11701 18921 11713 18955
rect 11747 18952 11759 18955
rect 11790 18952 11796 18964
rect 11747 18924 11796 18952
rect 11747 18921 11759 18924
rect 11701 18915 11759 18921
rect 11790 18912 11796 18924
rect 11848 18912 11854 18964
rect 22922 18912 22928 18964
rect 22980 18952 22986 18964
rect 23201 18955 23259 18961
rect 23201 18952 23213 18955
rect 22980 18924 23213 18952
rect 22980 18912 22986 18924
rect 23201 18921 23213 18924
rect 23247 18952 23259 18955
rect 26786 18952 26792 18964
rect 23247 18924 26648 18952
rect 26747 18924 26792 18952
rect 23247 18921 23259 18924
rect 23201 18915 23259 18921
rect 12989 18887 13047 18893
rect 12989 18853 13001 18887
rect 13035 18884 13047 18887
rect 13906 18884 13912 18896
rect 13035 18856 13912 18884
rect 13035 18853 13047 18856
rect 12989 18847 13047 18853
rect 13906 18844 13912 18856
rect 13964 18844 13970 18896
rect 24670 18844 24676 18896
rect 24728 18884 24734 18896
rect 24949 18887 25007 18893
rect 24949 18884 24961 18887
rect 24728 18856 24961 18884
rect 24728 18844 24734 18856
rect 24949 18853 24961 18856
rect 24995 18884 25007 18887
rect 25958 18884 25964 18896
rect 24995 18856 25964 18884
rect 24995 18853 25007 18856
rect 24949 18847 25007 18853
rect 25958 18844 25964 18856
rect 26016 18844 26022 18896
rect 26418 18884 26424 18896
rect 26068 18856 26424 18884
rect 12710 18816 12716 18828
rect 12671 18788 12716 18816
rect 12710 18776 12716 18788
rect 12768 18776 12774 18828
rect 2038 18708 2044 18760
rect 2096 18748 2102 18760
rect 2225 18751 2283 18757
rect 2225 18748 2237 18751
rect 2096 18720 2237 18748
rect 2096 18708 2102 18720
rect 2225 18717 2237 18720
rect 2271 18717 2283 18751
rect 2225 18711 2283 18717
rect 11885 18751 11943 18757
rect 11885 18717 11897 18751
rect 11931 18748 11943 18751
rect 12250 18748 12256 18760
rect 11931 18720 12256 18748
rect 11931 18717 11943 18720
rect 11885 18711 11943 18717
rect 12250 18708 12256 18720
rect 12308 18708 12314 18760
rect 12526 18708 12532 18760
rect 12584 18748 12590 18760
rect 12621 18751 12679 18757
rect 12621 18748 12633 18751
rect 12584 18720 12633 18748
rect 12584 18708 12590 18720
rect 12621 18717 12633 18720
rect 12667 18717 12679 18751
rect 12621 18711 12679 18717
rect 13906 18708 13912 18760
rect 13964 18748 13970 18760
rect 14921 18751 14979 18757
rect 14921 18748 14933 18751
rect 13964 18720 14933 18748
rect 13964 18708 13970 18720
rect 14921 18717 14933 18720
rect 14967 18717 14979 18751
rect 14921 18711 14979 18717
rect 15188 18751 15246 18757
rect 15188 18717 15200 18751
rect 15234 18748 15246 18751
rect 15470 18748 15476 18760
rect 15234 18720 15476 18748
rect 15234 18717 15246 18720
rect 15188 18711 15246 18717
rect 15470 18708 15476 18720
rect 15528 18708 15534 18760
rect 16758 18708 16764 18760
rect 16816 18748 16822 18760
rect 16945 18751 17003 18757
rect 16945 18748 16957 18751
rect 16816 18720 16957 18748
rect 16816 18708 16822 18720
rect 16945 18717 16957 18720
rect 16991 18748 17003 18751
rect 18138 18748 18144 18760
rect 16991 18720 18144 18748
rect 16991 18717 17003 18720
rect 16945 18711 17003 18717
rect 18138 18708 18144 18720
rect 18196 18708 18202 18760
rect 21821 18751 21879 18757
rect 21821 18717 21833 18751
rect 21867 18748 21879 18751
rect 24762 18748 24768 18760
rect 21867 18720 22784 18748
rect 24723 18720 24768 18748
rect 21867 18717 21879 18720
rect 21821 18711 21879 18717
rect 22756 18692 22784 18720
rect 24762 18708 24768 18720
rect 24820 18708 24826 18760
rect 26068 18757 26096 18856
rect 26418 18844 26424 18856
rect 26476 18844 26482 18896
rect 26326 18816 26332 18828
rect 26287 18788 26332 18816
rect 26326 18776 26332 18788
rect 26384 18776 26390 18828
rect 25041 18751 25099 18757
rect 25041 18717 25053 18751
rect 25087 18717 25099 18751
rect 25041 18711 25099 18717
rect 26053 18751 26111 18757
rect 26053 18717 26065 18751
rect 26099 18717 26111 18751
rect 26234 18748 26240 18760
rect 26195 18720 26240 18748
rect 26053 18711 26111 18717
rect 9950 18640 9956 18692
rect 10008 18680 10014 18692
rect 16390 18680 16396 18692
rect 10008 18652 16396 18680
rect 10008 18640 10014 18652
rect 16390 18640 16396 18652
rect 16448 18640 16454 18692
rect 17212 18683 17270 18689
rect 17212 18649 17224 18683
rect 17258 18680 17270 18683
rect 18230 18680 18236 18692
rect 17258 18652 18236 18680
rect 17258 18649 17270 18652
rect 17212 18643 17270 18649
rect 18230 18640 18236 18652
rect 18288 18640 18294 18692
rect 22088 18683 22146 18689
rect 22088 18649 22100 18683
rect 22134 18680 22146 18683
rect 22186 18680 22192 18692
rect 22134 18652 22192 18680
rect 22134 18649 22146 18652
rect 22088 18643 22146 18649
rect 22186 18640 22192 18652
rect 22244 18640 22250 18692
rect 22738 18640 22744 18692
rect 22796 18640 22802 18692
rect 16022 18572 16028 18624
rect 16080 18612 16086 18624
rect 16301 18615 16359 18621
rect 16301 18612 16313 18615
rect 16080 18584 16313 18612
rect 16080 18572 16086 18584
rect 16301 18581 16313 18584
rect 16347 18581 16359 18615
rect 16301 18575 16359 18581
rect 17862 18572 17868 18624
rect 17920 18612 17926 18624
rect 18325 18615 18383 18621
rect 18325 18612 18337 18615
rect 17920 18584 18337 18612
rect 17920 18572 17926 18584
rect 18325 18581 18337 18584
rect 18371 18581 18383 18615
rect 24578 18612 24584 18624
rect 24539 18584 24584 18612
rect 18325 18575 18383 18581
rect 24578 18572 24584 18584
rect 24636 18572 24642 18624
rect 25056 18612 25084 18711
rect 26234 18708 26240 18720
rect 26292 18708 26298 18760
rect 26620 18757 26648 18924
rect 26786 18912 26792 18924
rect 26844 18912 26850 18964
rect 27522 18912 27528 18964
rect 27580 18952 27586 18964
rect 28353 18955 28411 18961
rect 28353 18952 28365 18955
rect 27580 18924 28365 18952
rect 27580 18912 27586 18924
rect 28353 18921 28365 18924
rect 28399 18921 28411 18955
rect 28353 18915 28411 18921
rect 28721 18955 28779 18961
rect 28721 18921 28733 18955
rect 28767 18952 28779 18955
rect 28994 18952 29000 18964
rect 28767 18924 29000 18952
rect 28767 18921 28779 18924
rect 28721 18915 28779 18921
rect 28994 18912 29000 18924
rect 29052 18912 29058 18964
rect 31389 18955 31447 18961
rect 31389 18921 31401 18955
rect 31435 18952 31447 18955
rect 31478 18952 31484 18964
rect 31435 18924 31484 18952
rect 31435 18921 31447 18924
rect 31389 18915 31447 18921
rect 31478 18912 31484 18924
rect 31536 18912 31542 18964
rect 31570 18912 31576 18964
rect 31628 18952 31634 18964
rect 34146 18952 34152 18964
rect 31628 18924 34152 18952
rect 31628 18912 31634 18924
rect 34146 18912 34152 18924
rect 34204 18912 34210 18964
rect 35253 18955 35311 18961
rect 35253 18921 35265 18955
rect 35299 18952 35311 18955
rect 35434 18952 35440 18964
rect 35299 18924 35440 18952
rect 35299 18921 35311 18924
rect 35253 18915 35311 18921
rect 35434 18912 35440 18924
rect 35492 18912 35498 18964
rect 35526 18912 35532 18964
rect 35584 18952 35590 18964
rect 36262 18952 36268 18964
rect 35584 18924 36268 18952
rect 35584 18912 35590 18924
rect 36262 18912 36268 18924
rect 36320 18952 36326 18964
rect 38286 18952 38292 18964
rect 36320 18924 38292 18952
rect 36320 18912 36326 18924
rect 38286 18912 38292 18924
rect 38344 18912 38350 18964
rect 39022 18952 39028 18964
rect 38983 18924 39028 18952
rect 39022 18912 39028 18924
rect 39080 18912 39086 18964
rect 42150 18912 42156 18964
rect 42208 18952 42214 18964
rect 42613 18955 42671 18961
rect 42613 18952 42625 18955
rect 42208 18924 42625 18952
rect 42208 18912 42214 18924
rect 42613 18921 42625 18924
rect 42659 18921 42671 18955
rect 42613 18915 42671 18921
rect 27062 18844 27068 18896
rect 27120 18884 27126 18896
rect 31294 18884 31300 18896
rect 27120 18856 31300 18884
rect 27120 18844 27126 18856
rect 31294 18844 31300 18856
rect 31352 18844 31358 18896
rect 34514 18844 34520 18896
rect 34572 18884 34578 18896
rect 35894 18884 35900 18896
rect 34572 18856 35900 18884
rect 34572 18844 34578 18856
rect 35894 18844 35900 18856
rect 35952 18844 35958 18896
rect 37182 18844 37188 18896
rect 37240 18884 37246 18896
rect 40862 18884 40868 18896
rect 37240 18856 40868 18884
rect 37240 18844 37246 18856
rect 40862 18844 40868 18856
rect 40920 18884 40926 18896
rect 40920 18856 42932 18884
rect 40920 18844 40926 18856
rect 28534 18816 28540 18828
rect 26712 18788 28540 18816
rect 26421 18751 26479 18757
rect 26421 18717 26433 18751
rect 26467 18717 26479 18751
rect 26421 18711 26479 18717
rect 26605 18751 26663 18757
rect 26605 18717 26617 18751
rect 26651 18717 26663 18751
rect 26605 18711 26663 18717
rect 26436 18680 26464 18711
rect 26712 18680 26740 18788
rect 28534 18776 28540 18788
rect 28592 18776 28598 18828
rect 30834 18816 30840 18828
rect 30484 18788 30840 18816
rect 27522 18748 27528 18760
rect 27483 18720 27528 18748
rect 27522 18708 27528 18720
rect 27580 18708 27586 18760
rect 27801 18751 27859 18757
rect 27801 18717 27813 18751
rect 27847 18748 27859 18751
rect 28261 18751 28319 18757
rect 28261 18748 28273 18751
rect 27847 18720 28273 18748
rect 27847 18717 27859 18720
rect 27801 18711 27859 18717
rect 28261 18717 28273 18720
rect 28307 18717 28319 18751
rect 28261 18711 28319 18717
rect 30285 18751 30343 18757
rect 30285 18717 30297 18751
rect 30331 18748 30343 18751
rect 30374 18748 30380 18760
rect 30331 18720 30380 18748
rect 30331 18717 30343 18720
rect 30285 18711 30343 18717
rect 26436 18652 26740 18680
rect 27246 18640 27252 18692
rect 27304 18680 27310 18692
rect 27816 18680 27844 18711
rect 30374 18708 30380 18720
rect 30432 18708 30438 18760
rect 30484 18757 30512 18788
rect 30834 18776 30840 18788
rect 30892 18816 30898 18828
rect 31202 18816 31208 18828
rect 30892 18788 31208 18816
rect 30892 18776 30898 18788
rect 31202 18776 31208 18788
rect 31260 18776 31266 18828
rect 33134 18776 33140 18828
rect 33192 18816 33198 18828
rect 33778 18816 33784 18828
rect 33192 18788 33784 18816
rect 33192 18776 33198 18788
rect 33778 18776 33784 18788
rect 33836 18816 33842 18828
rect 34422 18816 34428 18828
rect 33836 18788 34428 18816
rect 33836 18776 33842 18788
rect 34422 18776 34428 18788
rect 34480 18776 34486 18828
rect 34790 18776 34796 18828
rect 34848 18816 34854 18828
rect 34848 18788 35112 18816
rect 34848 18776 34854 18788
rect 30469 18751 30527 18757
rect 30469 18717 30481 18751
rect 30515 18717 30527 18751
rect 30469 18711 30527 18717
rect 27304 18652 27844 18680
rect 27304 18640 27310 18652
rect 28534 18640 28540 18692
rect 28592 18680 28598 18692
rect 30484 18680 30512 18711
rect 30558 18708 30564 18760
rect 30616 18748 30622 18760
rect 33870 18748 33876 18760
rect 30616 18720 31754 18748
rect 33831 18720 33876 18748
rect 30616 18708 30622 18720
rect 31110 18680 31116 18692
rect 28592 18652 30512 18680
rect 31071 18652 31116 18680
rect 28592 18640 28598 18652
rect 31110 18640 31116 18652
rect 31168 18640 31174 18692
rect 26602 18612 26608 18624
rect 25056 18584 26608 18612
rect 26602 18572 26608 18584
rect 26660 18572 26666 18624
rect 27341 18615 27399 18621
rect 27341 18581 27353 18615
rect 27387 18612 27399 18615
rect 27430 18612 27436 18624
rect 27387 18584 27436 18612
rect 27387 18581 27399 18584
rect 27341 18575 27399 18581
rect 27430 18572 27436 18584
rect 27488 18572 27494 18624
rect 27709 18615 27767 18621
rect 27709 18581 27721 18615
rect 27755 18612 27767 18615
rect 29178 18612 29184 18624
rect 27755 18584 29184 18612
rect 27755 18581 27767 18584
rect 27709 18575 27767 18581
rect 29178 18572 29184 18584
rect 29236 18572 29242 18624
rect 30098 18612 30104 18624
rect 30059 18584 30104 18612
rect 30098 18572 30104 18584
rect 30156 18572 30162 18624
rect 31726 18612 31754 18720
rect 33870 18708 33876 18720
rect 33928 18708 33934 18760
rect 35084 18757 35112 18788
rect 35618 18776 35624 18828
rect 35676 18816 35682 18828
rect 35676 18788 35940 18816
rect 35676 18776 35682 18788
rect 33965 18751 34023 18757
rect 33965 18717 33977 18751
rect 34011 18748 34023 18751
rect 34977 18751 35035 18757
rect 34977 18748 34989 18751
rect 34011 18720 34989 18748
rect 34011 18717 34023 18720
rect 33965 18711 34023 18717
rect 34977 18717 34989 18720
rect 35023 18717 35035 18751
rect 34977 18711 35035 18717
rect 35069 18751 35127 18757
rect 35069 18717 35081 18751
rect 35115 18748 35127 18751
rect 35713 18751 35771 18757
rect 35713 18748 35725 18751
rect 35115 18720 35725 18748
rect 35115 18717 35127 18720
rect 35069 18711 35127 18717
rect 35713 18717 35725 18720
rect 35759 18748 35771 18751
rect 35802 18748 35808 18760
rect 35759 18720 35808 18748
rect 35759 18717 35771 18720
rect 35713 18711 35771 18717
rect 33686 18680 33692 18692
rect 33647 18652 33692 18680
rect 33686 18640 33692 18652
rect 33744 18640 33750 18692
rect 34882 18680 34888 18692
rect 33796 18652 34888 18680
rect 33796 18612 33824 18652
rect 34882 18640 34888 18652
rect 34940 18640 34946 18692
rect 34992 18680 35020 18711
rect 35802 18708 35808 18720
rect 35860 18708 35866 18760
rect 35912 18757 35940 18788
rect 42904 18760 42932 18856
rect 44450 18844 44456 18896
rect 44508 18844 44514 18896
rect 47946 18884 47952 18896
rect 46492 18856 47952 18884
rect 42981 18819 43039 18825
rect 42981 18785 42993 18819
rect 43027 18816 43039 18819
rect 44174 18816 44180 18828
rect 43027 18788 44180 18816
rect 43027 18785 43039 18788
rect 42981 18779 43039 18785
rect 35897 18751 35955 18757
rect 35897 18717 35909 18751
rect 35943 18717 35955 18751
rect 35897 18711 35955 18717
rect 38470 18708 38476 18760
rect 38528 18748 38534 18760
rect 38841 18751 38899 18757
rect 38841 18748 38853 18751
rect 38528 18720 38853 18748
rect 38528 18708 38534 18720
rect 38841 18717 38853 18720
rect 38887 18717 38899 18751
rect 38841 18711 38899 18717
rect 39114 18708 39120 18760
rect 39172 18748 39178 18760
rect 39172 18720 39217 18748
rect 39172 18708 39178 18720
rect 40126 18708 40132 18760
rect 40184 18748 40190 18760
rect 40770 18748 40776 18760
rect 40184 18720 40776 18748
rect 40184 18708 40190 18720
rect 40770 18708 40776 18720
rect 40828 18708 40834 18760
rect 42794 18748 42800 18760
rect 42755 18720 42800 18748
rect 42794 18708 42800 18720
rect 42852 18708 42858 18760
rect 42886 18708 42892 18760
rect 42944 18748 42950 18760
rect 42944 18720 42989 18748
rect 42944 18708 42950 18720
rect 43070 18708 43076 18760
rect 43128 18748 43134 18760
rect 44100 18757 44128 18788
rect 44174 18776 44180 18788
rect 44232 18776 44238 18828
rect 44468 18816 44496 18844
rect 46492 18825 46520 18856
rect 47946 18844 47952 18856
rect 48004 18844 48010 18896
rect 44376 18788 44496 18816
rect 46477 18819 46535 18825
rect 44085 18751 44143 18757
rect 43128 18720 43173 18748
rect 43128 18708 43134 18720
rect 44085 18717 44097 18751
rect 44131 18717 44143 18751
rect 44266 18748 44272 18760
rect 44227 18720 44272 18748
rect 44085 18711 44143 18717
rect 44266 18708 44272 18720
rect 44324 18708 44330 18760
rect 44376 18757 44404 18788
rect 46477 18785 46489 18819
rect 46523 18785 46535 18819
rect 46477 18779 46535 18785
rect 46661 18819 46719 18825
rect 46661 18785 46673 18819
rect 46707 18816 46719 18819
rect 47118 18816 47124 18828
rect 46707 18788 47124 18816
rect 46707 18785 46719 18788
rect 46661 18779 46719 18785
rect 47118 18776 47124 18788
rect 47176 18776 47182 18828
rect 48222 18816 48228 18828
rect 48183 18788 48228 18816
rect 48222 18776 48228 18788
rect 48280 18776 48286 18828
rect 44361 18751 44419 18757
rect 44361 18717 44373 18751
rect 44407 18717 44419 18751
rect 44361 18711 44419 18717
rect 44453 18751 44511 18757
rect 44453 18717 44465 18751
rect 44499 18717 44511 18751
rect 44453 18711 44511 18717
rect 36630 18680 36636 18692
rect 34992 18652 36636 18680
rect 36630 18640 36636 18652
rect 36688 18640 36694 18692
rect 41141 18683 41199 18689
rect 41141 18649 41153 18683
rect 41187 18680 41199 18683
rect 43346 18680 43352 18692
rect 41187 18652 43352 18680
rect 41187 18649 41199 18652
rect 41141 18643 41199 18649
rect 43346 18640 43352 18652
rect 43404 18680 43410 18692
rect 43530 18680 43536 18692
rect 43404 18652 43536 18680
rect 43404 18640 43410 18652
rect 43530 18640 43536 18652
rect 43588 18640 43594 18692
rect 44174 18640 44180 18692
rect 44232 18680 44238 18692
rect 44468 18680 44496 18711
rect 44232 18652 44496 18680
rect 44232 18640 44238 18652
rect 33962 18612 33968 18624
rect 31726 18584 33824 18612
rect 33923 18584 33968 18612
rect 33962 18572 33968 18584
rect 34020 18572 34026 18624
rect 35894 18612 35900 18624
rect 35855 18584 35900 18612
rect 35894 18572 35900 18584
rect 35952 18572 35958 18624
rect 38654 18612 38660 18624
rect 38615 18584 38660 18612
rect 38654 18572 38660 18584
rect 38712 18572 38718 18624
rect 44634 18612 44640 18624
rect 44595 18584 44640 18612
rect 44634 18572 44640 18584
rect 44692 18572 44698 18624
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 12250 18408 12256 18420
rect 12211 18380 12256 18408
rect 12250 18368 12256 18380
rect 12308 18368 12314 18420
rect 15933 18411 15991 18417
rect 15933 18377 15945 18411
rect 15979 18408 15991 18411
rect 15979 18380 16252 18408
rect 15979 18377 15991 18380
rect 15933 18371 15991 18377
rect 12621 18343 12679 18349
rect 12621 18309 12633 18343
rect 12667 18340 12679 18343
rect 16224 18340 16252 18380
rect 16390 18368 16396 18420
rect 16448 18408 16454 18420
rect 22281 18411 22339 18417
rect 16448 18380 21404 18408
rect 16448 18368 16454 18380
rect 17862 18340 17868 18352
rect 12667 18312 16068 18340
rect 16224 18312 17868 18340
rect 12667 18309 12679 18312
rect 12621 18303 12679 18309
rect 2038 18272 2044 18284
rect 1999 18244 2044 18272
rect 2038 18232 2044 18244
rect 2096 18232 2102 18284
rect 16040 18272 16068 18312
rect 17862 18300 17868 18312
rect 17920 18300 17926 18352
rect 21376 18340 21404 18380
rect 22281 18377 22293 18411
rect 22327 18408 22339 18411
rect 22370 18408 22376 18420
rect 22327 18380 22376 18408
rect 22327 18377 22339 18380
rect 22281 18371 22339 18377
rect 22370 18368 22376 18380
rect 22428 18368 22434 18420
rect 33594 18408 33600 18420
rect 23584 18380 33600 18408
rect 23584 18340 23612 18380
rect 33594 18368 33600 18380
rect 33652 18368 33658 18420
rect 36630 18408 36636 18420
rect 36591 18380 36636 18408
rect 36630 18368 36636 18380
rect 36688 18368 36694 18420
rect 38470 18408 38476 18420
rect 38431 18380 38476 18408
rect 38470 18368 38476 18380
rect 38528 18368 38534 18420
rect 41785 18411 41843 18417
rect 41785 18377 41797 18411
rect 41831 18377 41843 18411
rect 41785 18371 41843 18377
rect 21376 18312 23612 18340
rect 23652 18343 23710 18349
rect 23652 18309 23664 18343
rect 23698 18340 23710 18343
rect 24578 18340 24584 18352
rect 23698 18312 24584 18340
rect 23698 18309 23710 18312
rect 23652 18303 23710 18309
rect 24578 18300 24584 18312
rect 24636 18300 24642 18352
rect 26513 18343 26571 18349
rect 26513 18309 26525 18343
rect 26559 18340 26571 18343
rect 27246 18340 27252 18352
rect 26559 18312 27252 18340
rect 26559 18309 26571 18312
rect 26513 18303 26571 18309
rect 27246 18300 27252 18312
rect 27304 18300 27310 18352
rect 27522 18300 27528 18352
rect 27580 18340 27586 18352
rect 27580 18312 27936 18340
rect 27580 18300 27586 18312
rect 19058 18272 19064 18284
rect 16040 18244 19064 18272
rect 19058 18232 19064 18244
rect 19116 18232 19122 18284
rect 22278 18232 22284 18284
rect 22336 18272 22342 18284
rect 22465 18275 22523 18281
rect 22465 18272 22477 18275
rect 22336 18244 22477 18272
rect 22336 18232 22342 18244
rect 22465 18241 22477 18244
rect 22511 18241 22523 18275
rect 22741 18275 22799 18281
rect 22741 18272 22753 18275
rect 22465 18235 22523 18241
rect 22664 18244 22753 18272
rect 2222 18204 2228 18216
rect 2183 18176 2228 18204
rect 2222 18164 2228 18176
rect 2280 18164 2286 18216
rect 2774 18204 2780 18216
rect 2735 18176 2780 18204
rect 2774 18164 2780 18176
rect 2832 18164 2838 18216
rect 12710 18204 12716 18216
rect 12671 18176 12716 18204
rect 12710 18164 12716 18176
rect 12768 18164 12774 18216
rect 12897 18207 12955 18213
rect 12897 18173 12909 18207
rect 12943 18204 12955 18207
rect 13354 18204 13360 18216
rect 12943 18176 13360 18204
rect 12943 18173 12955 18176
rect 12897 18167 12955 18173
rect 13354 18164 13360 18176
rect 13412 18164 13418 18216
rect 16022 18204 16028 18216
rect 15983 18176 16028 18204
rect 16022 18164 16028 18176
rect 16080 18164 16086 18216
rect 16117 18207 16175 18213
rect 16117 18173 16129 18207
rect 16163 18173 16175 18207
rect 16117 18167 16175 18173
rect 19153 18207 19211 18213
rect 19153 18173 19165 18207
rect 19199 18173 19211 18207
rect 19153 18167 19211 18173
rect 19245 18207 19303 18213
rect 19245 18173 19257 18207
rect 19291 18204 19303 18207
rect 19334 18204 19340 18216
rect 19291 18176 19340 18204
rect 19291 18173 19303 18176
rect 19245 18167 19303 18173
rect 12618 18096 12624 18148
rect 12676 18136 12682 18148
rect 12676 18108 15700 18136
rect 12676 18096 12682 18108
rect 15194 18028 15200 18080
rect 15252 18068 15258 18080
rect 15565 18071 15623 18077
rect 15565 18068 15577 18071
rect 15252 18040 15577 18068
rect 15252 18028 15258 18040
rect 15565 18037 15577 18040
rect 15611 18037 15623 18071
rect 15672 18068 15700 18108
rect 15838 18096 15844 18148
rect 15896 18136 15902 18148
rect 16132 18136 16160 18167
rect 19168 18136 19196 18167
rect 19334 18164 19340 18176
rect 19392 18164 19398 18216
rect 22370 18164 22376 18216
rect 22428 18204 22434 18216
rect 22664 18204 22692 18244
rect 22741 18241 22753 18244
rect 22787 18241 22799 18275
rect 22922 18272 22928 18284
rect 22883 18244 22928 18272
rect 22741 18235 22799 18241
rect 22922 18232 22928 18244
rect 22980 18232 22986 18284
rect 26326 18232 26332 18284
rect 26384 18272 26390 18284
rect 26421 18275 26479 18281
rect 26421 18272 26433 18275
rect 26384 18244 26433 18272
rect 26384 18232 26390 18244
rect 26421 18241 26433 18244
rect 26467 18241 26479 18275
rect 26421 18235 26479 18241
rect 26602 18232 26608 18284
rect 26660 18272 26666 18284
rect 27338 18272 27344 18284
rect 26660 18244 27344 18272
rect 26660 18232 26666 18244
rect 27338 18232 27344 18244
rect 27396 18232 27402 18284
rect 27706 18272 27712 18284
rect 27667 18244 27712 18272
rect 27706 18232 27712 18244
rect 27764 18232 27770 18284
rect 27908 18281 27936 18312
rect 30098 18300 30104 18352
rect 30156 18340 30162 18352
rect 30622 18343 30680 18349
rect 30622 18340 30634 18343
rect 30156 18312 30634 18340
rect 30156 18300 30162 18312
rect 30622 18309 30634 18312
rect 30668 18309 30680 18343
rect 30622 18303 30680 18309
rect 33781 18343 33839 18349
rect 33781 18309 33793 18343
rect 33827 18340 33839 18343
rect 33870 18340 33876 18352
rect 33827 18312 33876 18340
rect 33827 18309 33839 18312
rect 33781 18303 33839 18309
rect 33870 18300 33876 18312
rect 33928 18300 33934 18352
rect 34011 18309 34069 18315
rect 34011 18306 34023 18309
rect 27893 18275 27951 18281
rect 27893 18241 27905 18275
rect 27939 18241 27951 18275
rect 27893 18235 27951 18241
rect 27985 18275 28043 18281
rect 27985 18241 27997 18275
rect 28031 18241 28043 18275
rect 27985 18235 28043 18241
rect 23385 18207 23443 18213
rect 23385 18204 23397 18207
rect 22428 18176 22692 18204
rect 22756 18176 23397 18204
rect 22428 18164 22434 18176
rect 22756 18148 22784 18176
rect 23385 18173 23397 18176
rect 23431 18173 23443 18207
rect 23385 18167 23443 18173
rect 22646 18136 22652 18148
rect 15896 18108 16160 18136
rect 16546 18108 22652 18136
rect 15896 18096 15902 18108
rect 16546 18068 16574 18108
rect 22646 18096 22652 18108
rect 22704 18096 22710 18148
rect 22738 18096 22744 18148
rect 22796 18096 22802 18148
rect 24765 18139 24823 18145
rect 24765 18105 24777 18139
rect 24811 18136 24823 18139
rect 26620 18136 26648 18232
rect 27522 18164 27528 18216
rect 27580 18204 27586 18216
rect 28000 18204 28028 18235
rect 28166 18232 28172 18284
rect 28224 18272 28230 18284
rect 28537 18275 28595 18281
rect 28537 18272 28549 18275
rect 28224 18244 28549 18272
rect 28224 18232 28230 18244
rect 28537 18241 28549 18244
rect 28583 18241 28595 18275
rect 28537 18235 28595 18241
rect 28626 18232 28632 18284
rect 28684 18272 28690 18284
rect 28684 18244 28729 18272
rect 28684 18232 28690 18244
rect 30282 18232 30288 18284
rect 30340 18272 30346 18284
rect 30377 18275 30435 18281
rect 30377 18272 30389 18275
rect 30340 18244 30389 18272
rect 30340 18232 30346 18244
rect 30377 18241 30389 18244
rect 30423 18241 30435 18275
rect 33229 18275 33287 18281
rect 33229 18272 33241 18275
rect 30377 18235 30435 18241
rect 30484 18244 33241 18272
rect 27580 18176 28028 18204
rect 27580 18164 27586 18176
rect 27801 18139 27859 18145
rect 24811 18108 26648 18136
rect 27172 18108 27752 18136
rect 24811 18105 24823 18108
rect 24765 18099 24823 18105
rect 18690 18068 18696 18080
rect 15672 18040 16574 18068
rect 18651 18040 18696 18068
rect 15565 18031 15623 18037
rect 18690 18028 18696 18040
rect 18748 18028 18754 18080
rect 23566 18028 23572 18080
rect 23624 18068 23630 18080
rect 27172 18068 27200 18108
rect 23624 18040 27200 18068
rect 23624 18028 23630 18040
rect 27246 18028 27252 18080
rect 27304 18068 27310 18080
rect 27525 18071 27583 18077
rect 27525 18068 27537 18071
rect 27304 18040 27537 18068
rect 27304 18028 27310 18040
rect 27525 18037 27537 18040
rect 27571 18037 27583 18071
rect 27724 18068 27752 18108
rect 27801 18105 27813 18139
rect 27847 18136 27859 18139
rect 27982 18136 27988 18148
rect 27847 18108 27988 18136
rect 27847 18105 27859 18108
rect 27801 18099 27859 18105
rect 27982 18096 27988 18108
rect 28040 18136 28046 18148
rect 28644 18136 28672 18232
rect 30484 18204 30512 18244
rect 33229 18241 33241 18244
rect 33275 18241 33287 18275
rect 33996 18275 34023 18306
rect 34057 18284 34069 18309
rect 35894 18300 35900 18352
rect 35952 18340 35958 18352
rect 35952 18312 36768 18340
rect 35952 18300 35958 18312
rect 34057 18275 34060 18284
rect 33996 18244 34060 18275
rect 33229 18235 33287 18241
rect 34054 18232 34060 18244
rect 34112 18232 34118 18284
rect 36446 18272 36452 18284
rect 36407 18244 36452 18272
rect 36446 18232 36452 18244
rect 36504 18232 36510 18284
rect 36740 18281 36768 18312
rect 37182 18300 37188 18352
rect 37240 18340 37246 18352
rect 37645 18343 37703 18349
rect 37645 18340 37657 18343
rect 37240 18312 37657 18340
rect 37240 18300 37246 18312
rect 37645 18309 37657 18312
rect 37691 18309 37703 18343
rect 40586 18340 40592 18352
rect 37645 18303 37703 18309
rect 38028 18312 40592 18340
rect 36725 18275 36783 18281
rect 36725 18241 36737 18275
rect 36771 18272 36783 18275
rect 36998 18272 37004 18284
rect 36771 18244 37004 18272
rect 36771 18241 36783 18244
rect 36725 18235 36783 18241
rect 36998 18232 37004 18244
rect 37056 18232 37062 18284
rect 37461 18275 37519 18281
rect 37461 18241 37473 18275
rect 37507 18272 37519 18275
rect 37550 18272 37556 18284
rect 37507 18244 37556 18272
rect 37507 18241 37519 18244
rect 37461 18235 37519 18241
rect 37550 18232 37556 18244
rect 37608 18232 37614 18284
rect 37918 18281 37924 18284
rect 37737 18278 37795 18281
rect 37721 18275 37795 18278
rect 37721 18272 37749 18275
rect 37660 18244 37749 18272
rect 32950 18204 32956 18216
rect 28920 18176 30512 18204
rect 32911 18176 32956 18204
rect 28920 18145 28948 18176
rect 32950 18164 32956 18176
rect 33008 18164 33014 18216
rect 33045 18207 33103 18213
rect 33045 18173 33057 18207
rect 33091 18173 33103 18207
rect 33045 18167 33103 18173
rect 28040 18108 28672 18136
rect 28905 18139 28963 18145
rect 28040 18096 28046 18108
rect 28905 18105 28917 18139
rect 28951 18105 28963 18139
rect 31754 18136 31760 18148
rect 31667 18108 31760 18136
rect 28905 18099 28963 18105
rect 31754 18096 31760 18108
rect 31812 18136 31818 18148
rect 33060 18136 33088 18167
rect 33134 18164 33140 18216
rect 33192 18204 33198 18216
rect 33192 18176 33237 18204
rect 33192 18164 33198 18176
rect 33318 18164 33324 18216
rect 33376 18204 33382 18216
rect 37660 18204 37688 18244
rect 37737 18241 37749 18244
rect 37783 18241 37795 18275
rect 37737 18235 37795 18241
rect 37865 18275 37924 18281
rect 37865 18241 37877 18275
rect 37911 18241 37924 18275
rect 37865 18235 37924 18241
rect 37918 18232 37924 18235
rect 37976 18272 37982 18284
rect 38028 18272 38056 18312
rect 40586 18300 40592 18312
rect 40644 18300 40650 18352
rect 41690 18300 41696 18352
rect 41748 18340 41754 18352
rect 41800 18340 41828 18371
rect 42610 18368 42616 18420
rect 42668 18408 42674 18420
rect 43641 18411 43699 18417
rect 43641 18408 43653 18411
rect 42668 18380 43653 18408
rect 42668 18368 42674 18380
rect 43641 18377 43653 18380
rect 43687 18377 43699 18411
rect 43806 18408 43812 18420
rect 43767 18380 43812 18408
rect 43641 18371 43699 18377
rect 43806 18368 43812 18380
rect 43864 18368 43870 18420
rect 44450 18368 44456 18420
rect 44508 18408 44514 18420
rect 46201 18411 46259 18417
rect 46201 18408 46213 18411
rect 44508 18380 46213 18408
rect 44508 18368 44514 18380
rect 46201 18377 46213 18380
rect 46247 18408 46259 18411
rect 46474 18408 46480 18420
rect 46247 18380 46480 18408
rect 46247 18377 46259 18380
rect 46201 18371 46259 18377
rect 46474 18368 46480 18380
rect 46532 18368 46538 18420
rect 42705 18343 42763 18349
rect 42705 18340 42717 18343
rect 41748 18312 42717 18340
rect 41748 18300 41754 18312
rect 42705 18309 42717 18312
rect 42751 18340 42763 18343
rect 43441 18343 43499 18349
rect 43441 18340 43453 18343
rect 42751 18312 43453 18340
rect 42751 18309 42763 18312
rect 42705 18303 42763 18309
rect 43441 18309 43453 18312
rect 43487 18340 43499 18343
rect 43990 18340 43996 18352
rect 43487 18312 43996 18340
rect 43487 18309 43499 18312
rect 43441 18303 43499 18309
rect 43990 18300 43996 18312
rect 44048 18300 44054 18352
rect 44634 18300 44640 18352
rect 44692 18340 44698 18352
rect 45066 18343 45124 18349
rect 45066 18340 45078 18343
rect 44692 18312 45078 18340
rect 44692 18300 44698 18312
rect 45066 18309 45078 18312
rect 45112 18309 45124 18343
rect 45066 18303 45124 18309
rect 38657 18275 38715 18281
rect 37976 18244 38069 18272
rect 37976 18232 37982 18244
rect 38657 18241 38669 18275
rect 38703 18272 38715 18275
rect 38746 18272 38752 18284
rect 38703 18244 38752 18272
rect 38703 18241 38715 18244
rect 38657 18235 38715 18241
rect 38746 18232 38752 18244
rect 38804 18232 38810 18284
rect 38930 18272 38936 18284
rect 38891 18244 38936 18272
rect 38930 18232 38936 18244
rect 38988 18232 38994 18284
rect 40678 18281 40684 18284
rect 39117 18275 39175 18281
rect 39117 18241 39129 18275
rect 39163 18241 39175 18275
rect 39117 18235 39175 18241
rect 40672 18235 40684 18281
rect 40736 18272 40742 18284
rect 40736 18244 40772 18272
rect 33376 18176 37688 18204
rect 33376 18164 33382 18176
rect 34146 18136 34152 18148
rect 31812 18108 32996 18136
rect 33060 18108 34008 18136
rect 34107 18108 34152 18136
rect 31812 18096 31818 18108
rect 28534 18068 28540 18080
rect 27724 18040 28540 18068
rect 27525 18031 27583 18037
rect 28534 18028 28540 18040
rect 28592 18028 28598 18080
rect 28721 18071 28779 18077
rect 28721 18037 28733 18071
rect 28767 18068 28779 18071
rect 28994 18068 29000 18080
rect 28767 18040 29000 18068
rect 28767 18037 28779 18040
rect 28721 18031 28779 18037
rect 28994 18028 29000 18040
rect 29052 18028 29058 18080
rect 31846 18028 31852 18080
rect 31904 18068 31910 18080
rect 32769 18071 32827 18077
rect 32769 18068 32781 18071
rect 31904 18040 32781 18068
rect 31904 18028 31910 18040
rect 32769 18037 32781 18040
rect 32815 18037 32827 18071
rect 32968 18068 32996 18108
rect 33980 18080 34008 18108
rect 34146 18096 34152 18108
rect 34204 18096 34210 18148
rect 34882 18096 34888 18148
rect 34940 18136 34946 18148
rect 39132 18136 39160 18235
rect 40678 18232 40684 18235
rect 40736 18232 40742 18244
rect 42058 18232 42064 18284
rect 42116 18272 42122 18284
rect 42610 18272 42616 18284
rect 42116 18244 42616 18272
rect 42116 18232 42122 18244
rect 42610 18232 42616 18244
rect 42668 18232 42674 18284
rect 42978 18272 42984 18284
rect 42939 18244 42984 18272
rect 42978 18232 42984 18244
rect 43036 18232 43042 18284
rect 44358 18232 44364 18284
rect 44416 18272 44422 18284
rect 44821 18275 44879 18281
rect 44821 18272 44833 18275
rect 44416 18244 44833 18272
rect 44416 18232 44422 18244
rect 44821 18241 44833 18244
rect 44867 18241 44879 18275
rect 44821 18235 44879 18241
rect 46566 18232 46572 18284
rect 46624 18272 46630 18284
rect 46753 18275 46811 18281
rect 46753 18272 46765 18275
rect 46624 18244 46765 18272
rect 46624 18232 46630 18244
rect 46753 18241 46765 18244
rect 46799 18241 46811 18275
rect 46753 18235 46811 18241
rect 47670 18232 47676 18284
rect 47728 18272 47734 18284
rect 47765 18275 47823 18281
rect 47765 18272 47777 18275
rect 47728 18244 47777 18272
rect 47728 18232 47734 18244
rect 47765 18241 47777 18244
rect 47811 18241 47823 18275
rect 47765 18235 47823 18241
rect 40402 18204 40408 18216
rect 40363 18176 40408 18204
rect 40402 18164 40408 18176
rect 40460 18164 40466 18216
rect 42702 18164 42708 18216
rect 42760 18204 42766 18216
rect 42797 18207 42855 18213
rect 42797 18204 42809 18207
rect 42760 18176 42809 18204
rect 42760 18164 42766 18176
rect 42797 18173 42809 18176
rect 42843 18173 42855 18207
rect 42797 18167 42855 18173
rect 39666 18136 39672 18148
rect 34940 18108 39672 18136
rect 34940 18096 34946 18108
rect 39666 18096 39672 18108
rect 39724 18096 39730 18148
rect 46750 18096 46756 18148
rect 46808 18136 46814 18148
rect 47857 18139 47915 18145
rect 47857 18136 47869 18139
rect 46808 18108 47869 18136
rect 46808 18096 46814 18108
rect 47857 18105 47869 18108
rect 47903 18105 47915 18139
rect 47857 18099 47915 18105
rect 33318 18068 33324 18080
rect 32968 18040 33324 18068
rect 32769 18031 32827 18037
rect 33318 18028 33324 18040
rect 33376 18028 33382 18080
rect 33962 18068 33968 18080
rect 33923 18040 33968 18068
rect 33962 18028 33968 18040
rect 34020 18028 34026 18080
rect 36449 18071 36507 18077
rect 36449 18037 36461 18071
rect 36495 18068 36507 18071
rect 36630 18068 36636 18080
rect 36495 18040 36636 18068
rect 36495 18037 36507 18040
rect 36449 18031 36507 18037
rect 36630 18028 36636 18040
rect 36688 18028 36694 18080
rect 37274 18028 37280 18080
rect 37332 18068 37338 18080
rect 37461 18071 37519 18077
rect 37461 18068 37473 18071
rect 37332 18040 37473 18068
rect 37332 18028 37338 18040
rect 37461 18037 37473 18040
rect 37507 18037 37519 18071
rect 37461 18031 37519 18037
rect 42981 18071 43039 18077
rect 42981 18037 42993 18071
rect 43027 18068 43039 18071
rect 43254 18068 43260 18080
rect 43027 18040 43260 18068
rect 43027 18037 43039 18040
rect 42981 18031 43039 18037
rect 43254 18028 43260 18040
rect 43312 18028 43318 18080
rect 43438 18028 43444 18080
rect 43496 18068 43502 18080
rect 43625 18071 43683 18077
rect 43625 18068 43637 18071
rect 43496 18040 43637 18068
rect 43496 18028 43502 18040
rect 43625 18037 43637 18040
rect 43671 18037 43683 18071
rect 43625 18031 43683 18037
rect 46658 18028 46664 18080
rect 46716 18068 46722 18080
rect 46845 18071 46903 18077
rect 46845 18068 46857 18071
rect 46716 18040 46857 18068
rect 46716 18028 46722 18040
rect 46845 18037 46857 18040
rect 46891 18037 46903 18071
rect 46845 18031 46903 18037
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 2222 17824 2228 17876
rect 2280 17864 2286 17876
rect 2317 17867 2375 17873
rect 2317 17864 2329 17867
rect 2280 17836 2329 17864
rect 2280 17824 2286 17836
rect 2317 17833 2329 17836
rect 2363 17833 2375 17867
rect 2317 17827 2375 17833
rect 12710 17824 12716 17876
rect 12768 17864 12774 17876
rect 12897 17867 12955 17873
rect 12897 17864 12909 17867
rect 12768 17836 12909 17864
rect 12768 17824 12774 17836
rect 12897 17833 12909 17836
rect 12943 17833 12955 17867
rect 23566 17864 23572 17876
rect 23527 17836 23572 17864
rect 12897 17827 12955 17833
rect 23566 17824 23572 17836
rect 23624 17824 23630 17876
rect 28074 17824 28080 17876
rect 28132 17864 28138 17876
rect 28813 17867 28871 17873
rect 28813 17864 28825 17867
rect 28132 17836 28825 17864
rect 28132 17824 28138 17836
rect 28813 17833 28825 17836
rect 28859 17833 28871 17867
rect 28813 17827 28871 17833
rect 30374 17824 30380 17876
rect 30432 17864 30438 17876
rect 30837 17867 30895 17873
rect 30837 17864 30849 17867
rect 30432 17836 30849 17864
rect 30432 17824 30438 17836
rect 30837 17833 30849 17836
rect 30883 17833 30895 17867
rect 30837 17827 30895 17833
rect 32950 17824 32956 17876
rect 33008 17864 33014 17876
rect 34054 17864 34060 17876
rect 33008 17836 34060 17864
rect 33008 17824 33014 17836
rect 34054 17824 34060 17836
rect 34112 17824 34118 17876
rect 35894 17864 35900 17876
rect 35636 17836 35900 17864
rect 18690 17796 18696 17808
rect 18651 17768 18696 17796
rect 18690 17756 18696 17768
rect 18748 17756 18754 17808
rect 28258 17796 28264 17808
rect 28219 17768 28264 17796
rect 28258 17756 28264 17768
rect 28316 17756 28322 17808
rect 11514 17728 11520 17740
rect 11475 17700 11520 17728
rect 11514 17688 11520 17700
rect 11572 17688 11578 17740
rect 18785 17731 18843 17737
rect 18785 17697 18797 17731
rect 18831 17728 18843 17731
rect 18831 17700 19656 17728
rect 18831 17697 18843 17700
rect 18785 17691 18843 17697
rect 2225 17663 2283 17669
rect 2225 17629 2237 17663
rect 2271 17660 2283 17663
rect 2314 17660 2320 17672
rect 2271 17632 2320 17660
rect 2271 17629 2283 17632
rect 2225 17623 2283 17629
rect 2314 17620 2320 17632
rect 2372 17620 2378 17672
rect 15194 17660 15200 17672
rect 15155 17632 15200 17660
rect 15194 17620 15200 17632
rect 15252 17620 15258 17672
rect 18325 17663 18383 17669
rect 18325 17629 18337 17663
rect 18371 17660 18383 17663
rect 18506 17660 18512 17672
rect 18371 17632 18512 17660
rect 18371 17629 18383 17632
rect 18325 17623 18383 17629
rect 18506 17620 18512 17632
rect 18564 17660 18570 17672
rect 18874 17660 18880 17672
rect 18564 17632 18880 17660
rect 18564 17620 18570 17632
rect 18874 17620 18880 17632
rect 18932 17620 18938 17672
rect 19628 17669 19656 17700
rect 27982 17688 27988 17740
rect 28040 17728 28046 17740
rect 28169 17731 28227 17737
rect 28169 17728 28181 17731
rect 28040 17700 28181 17728
rect 28040 17688 28046 17700
rect 28169 17697 28181 17700
rect 28215 17697 28227 17731
rect 28169 17691 28227 17697
rect 28353 17731 28411 17737
rect 28353 17697 28365 17731
rect 28399 17728 28411 17731
rect 29178 17728 29184 17740
rect 28399 17700 29184 17728
rect 28399 17697 28411 17700
rect 28353 17691 28411 17697
rect 29178 17688 29184 17700
rect 29236 17688 29242 17740
rect 19613 17663 19671 17669
rect 19613 17629 19625 17663
rect 19659 17629 19671 17663
rect 19613 17623 19671 17629
rect 22005 17663 22063 17669
rect 22005 17629 22017 17663
rect 22051 17660 22063 17663
rect 22094 17660 22100 17672
rect 22051 17632 22100 17660
rect 22051 17629 22063 17632
rect 22005 17623 22063 17629
rect 22094 17620 22100 17632
rect 22152 17620 22158 17672
rect 22646 17620 22652 17672
rect 22704 17660 22710 17672
rect 23477 17663 23535 17669
rect 23477 17660 23489 17663
rect 22704 17632 23489 17660
rect 22704 17620 22710 17632
rect 23477 17629 23489 17632
rect 23523 17660 23535 17663
rect 25130 17660 25136 17672
rect 23523 17632 25136 17660
rect 23523 17629 23535 17632
rect 23477 17623 23535 17629
rect 25130 17620 25136 17632
rect 25188 17620 25194 17672
rect 27706 17620 27712 17672
rect 27764 17660 27770 17672
rect 28077 17663 28135 17669
rect 28077 17660 28089 17663
rect 27764 17632 28089 17660
rect 27764 17620 27770 17632
rect 28077 17629 28089 17632
rect 28123 17629 28135 17663
rect 28077 17623 28135 17629
rect 28994 17620 29000 17672
rect 29052 17660 29058 17672
rect 29089 17663 29147 17669
rect 29089 17660 29101 17663
rect 29052 17632 29101 17660
rect 29052 17620 29058 17632
rect 29089 17629 29101 17632
rect 29135 17629 29147 17663
rect 31018 17660 31024 17672
rect 30979 17632 31024 17660
rect 29089 17623 29147 17629
rect 31018 17620 31024 17632
rect 31076 17620 31082 17672
rect 31297 17663 31355 17669
rect 31297 17629 31309 17663
rect 31343 17660 31355 17663
rect 31386 17660 31392 17672
rect 31343 17632 31392 17660
rect 31343 17629 31355 17632
rect 31297 17623 31355 17629
rect 31386 17620 31392 17632
rect 31444 17620 31450 17672
rect 31481 17663 31539 17669
rect 31481 17629 31493 17663
rect 31527 17660 31539 17663
rect 31754 17660 31760 17672
rect 31527 17632 31760 17660
rect 31527 17629 31539 17632
rect 31481 17623 31539 17629
rect 31754 17620 31760 17632
rect 31812 17620 31818 17672
rect 34606 17620 34612 17672
rect 34664 17660 34670 17672
rect 35636 17669 35664 17836
rect 35894 17824 35900 17836
rect 35952 17824 35958 17876
rect 39114 17824 39120 17876
rect 39172 17864 39178 17876
rect 39485 17867 39543 17873
rect 39485 17864 39497 17867
rect 39172 17836 39497 17864
rect 39172 17824 39178 17836
rect 39485 17833 39497 17836
rect 39531 17833 39543 17867
rect 39485 17827 39543 17833
rect 40678 17824 40684 17876
rect 40736 17864 40742 17876
rect 40865 17867 40923 17873
rect 40865 17864 40877 17867
rect 40736 17836 40877 17864
rect 40736 17824 40742 17836
rect 40865 17833 40877 17836
rect 40911 17833 40923 17867
rect 44177 17867 44235 17873
rect 44177 17864 44189 17867
rect 40865 17827 40923 17833
rect 41984 17836 44189 17864
rect 36722 17796 36728 17808
rect 35728 17768 36728 17796
rect 35529 17663 35587 17669
rect 35529 17660 35541 17663
rect 34664 17632 35541 17660
rect 34664 17620 34670 17632
rect 35529 17629 35541 17632
rect 35575 17629 35587 17663
rect 35529 17623 35587 17629
rect 35621 17663 35679 17669
rect 35621 17629 35633 17663
rect 35667 17629 35679 17663
rect 35621 17623 35679 17629
rect 11784 17595 11842 17601
rect 11784 17561 11796 17595
rect 11830 17592 11842 17595
rect 12066 17592 12072 17604
rect 11830 17564 12072 17592
rect 11830 17561 11842 17564
rect 11784 17555 11842 17561
rect 12066 17552 12072 17564
rect 12124 17552 12130 17604
rect 22738 17592 22744 17604
rect 22699 17564 22744 17592
rect 22738 17552 22744 17564
rect 22796 17552 22802 17604
rect 28442 17552 28448 17604
rect 28500 17592 28506 17604
rect 28626 17592 28632 17604
rect 28500 17564 28632 17592
rect 28500 17552 28506 17564
rect 28626 17552 28632 17564
rect 28684 17592 28690 17604
rect 28813 17595 28871 17601
rect 28813 17592 28825 17595
rect 28684 17564 28825 17592
rect 28684 17552 28690 17564
rect 28813 17561 28825 17564
rect 28859 17561 28871 17595
rect 28813 17555 28871 17561
rect 15010 17524 15016 17536
rect 14971 17496 15016 17524
rect 15010 17484 15016 17496
rect 15068 17484 15074 17536
rect 19426 17524 19432 17536
rect 19387 17496 19432 17524
rect 19426 17484 19432 17496
rect 19484 17484 19490 17536
rect 28258 17484 28264 17536
rect 28316 17524 28322 17536
rect 28997 17527 29055 17533
rect 28997 17524 29009 17527
rect 28316 17496 29009 17524
rect 28316 17484 28322 17496
rect 28997 17493 29009 17496
rect 29043 17493 29055 17527
rect 35342 17524 35348 17536
rect 35303 17496 35348 17524
rect 28997 17487 29055 17493
rect 35342 17484 35348 17496
rect 35400 17484 35406 17536
rect 35544 17524 35572 17623
rect 35728 17601 35756 17768
rect 36722 17756 36728 17768
rect 36780 17796 36786 17808
rect 36780 17768 37136 17796
rect 36780 17756 36786 17768
rect 36998 17728 37004 17740
rect 36959 17700 37004 17728
rect 36998 17688 37004 17700
rect 37056 17688 37062 17740
rect 37108 17737 37136 17768
rect 37093 17731 37151 17737
rect 37093 17697 37105 17731
rect 37139 17697 37151 17731
rect 41984 17728 42012 17836
rect 44177 17833 44189 17836
rect 44223 17833 44235 17867
rect 44177 17827 44235 17833
rect 44361 17799 44419 17805
rect 44361 17796 44373 17799
rect 37093 17691 37151 17697
rect 41892 17700 42012 17728
rect 43180 17768 44373 17796
rect 35986 17620 35992 17672
rect 36044 17660 36050 17672
rect 36446 17660 36452 17672
rect 36044 17632 36089 17660
rect 36188 17632 36452 17660
rect 36044 17620 36050 17632
rect 35713 17595 35771 17601
rect 35713 17561 35725 17595
rect 35759 17561 35771 17595
rect 35713 17555 35771 17561
rect 35802 17552 35808 17604
rect 35860 17601 35866 17604
rect 35860 17595 35889 17601
rect 35877 17561 35889 17595
rect 35860 17555 35889 17561
rect 35860 17552 35866 17555
rect 36188 17524 36216 17632
rect 36446 17620 36452 17632
rect 36504 17660 36510 17672
rect 36906 17660 36912 17672
rect 36504 17632 36912 17660
rect 36504 17620 36510 17632
rect 36906 17620 36912 17632
rect 36964 17620 36970 17672
rect 37185 17663 37243 17669
rect 37185 17629 37197 17663
rect 37231 17660 37243 17663
rect 37366 17660 37372 17672
rect 37231 17632 37372 17660
rect 37231 17629 37243 17632
rect 37185 17623 37243 17629
rect 37366 17620 37372 17632
rect 37424 17620 37430 17672
rect 37458 17620 37464 17672
rect 37516 17660 37522 17672
rect 38105 17663 38163 17669
rect 38105 17660 38117 17663
rect 37516 17632 38117 17660
rect 37516 17620 37522 17632
rect 38105 17629 38117 17632
rect 38151 17629 38163 17663
rect 38105 17623 38163 17629
rect 38372 17663 38430 17669
rect 38372 17629 38384 17663
rect 38418 17660 38430 17663
rect 38654 17660 38660 17672
rect 38418 17632 38660 17660
rect 38418 17629 38430 17632
rect 38372 17623 38430 17629
rect 38654 17620 38660 17632
rect 38712 17620 38718 17672
rect 41046 17660 41052 17672
rect 41007 17632 41052 17660
rect 41046 17620 41052 17632
rect 41104 17620 41110 17672
rect 41690 17660 41696 17672
rect 41651 17632 41696 17660
rect 41690 17620 41696 17632
rect 41748 17620 41754 17672
rect 41892 17669 41920 17700
rect 41877 17663 41935 17669
rect 41877 17629 41889 17663
rect 41923 17629 41935 17663
rect 41877 17623 41935 17629
rect 41969 17663 42027 17669
rect 41969 17629 41981 17663
rect 42015 17660 42027 17663
rect 42058 17660 42064 17672
rect 42015 17632 42064 17660
rect 42015 17629 42027 17632
rect 41969 17623 42027 17629
rect 40770 17552 40776 17604
rect 40828 17592 40834 17604
rect 41892 17592 41920 17623
rect 42058 17620 42064 17632
rect 42116 17620 42122 17672
rect 43180 17669 43208 17768
rect 44361 17765 44373 17768
rect 44407 17765 44419 17799
rect 44361 17759 44419 17765
rect 43438 17728 43444 17740
rect 43399 17700 43444 17728
rect 43438 17688 43444 17700
rect 43496 17688 43502 17740
rect 46474 17728 46480 17740
rect 46435 17700 46480 17728
rect 46474 17688 46480 17700
rect 46532 17688 46538 17740
rect 46658 17728 46664 17740
rect 46619 17700 46664 17728
rect 46658 17688 46664 17700
rect 46716 17688 46722 17740
rect 48038 17728 48044 17740
rect 47999 17700 48044 17728
rect 48038 17688 48044 17700
rect 48096 17688 48102 17740
rect 43165 17663 43223 17669
rect 43165 17629 43177 17663
rect 43211 17629 43223 17663
rect 43165 17623 43223 17629
rect 40828 17564 41920 17592
rect 42076 17592 42104 17620
rect 43990 17592 43996 17604
rect 42076 17564 43392 17592
rect 43951 17564 43996 17592
rect 40828 17552 40834 17564
rect 36722 17524 36728 17536
rect 35544 17496 36216 17524
rect 36683 17496 36728 17524
rect 36722 17484 36728 17496
rect 36780 17484 36786 17536
rect 41509 17527 41567 17533
rect 41509 17493 41521 17527
rect 41555 17524 41567 17527
rect 41598 17524 41604 17536
rect 41555 17496 41604 17524
rect 41555 17493 41567 17496
rect 41509 17487 41567 17493
rect 41598 17484 41604 17496
rect 41656 17484 41662 17536
rect 42794 17524 42800 17536
rect 42755 17496 42800 17524
rect 42794 17484 42800 17496
rect 42852 17484 42858 17536
rect 43254 17524 43260 17536
rect 43215 17496 43260 17524
rect 43254 17484 43260 17496
rect 43312 17484 43318 17536
rect 43364 17524 43392 17564
rect 43990 17552 43996 17564
rect 44048 17552 44054 17604
rect 44193 17527 44251 17533
rect 44193 17524 44205 17527
rect 43364 17496 44205 17524
rect 44193 17493 44205 17496
rect 44239 17493 44251 17527
rect 44193 17487 44251 17493
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 12066 17320 12072 17332
rect 12027 17292 12072 17320
rect 12066 17280 12072 17292
rect 12124 17280 12130 17332
rect 19058 17280 19064 17332
rect 19116 17320 19122 17332
rect 19797 17323 19855 17329
rect 19797 17320 19809 17323
rect 19116 17292 19809 17320
rect 19116 17280 19122 17292
rect 19797 17289 19809 17292
rect 19843 17289 19855 17323
rect 26234 17320 26240 17332
rect 26195 17292 26240 17320
rect 19797 17283 19855 17289
rect 26234 17280 26240 17292
rect 26292 17280 26298 17332
rect 35805 17323 35863 17329
rect 35805 17320 35817 17323
rect 33888 17292 35817 17320
rect 11514 17212 11520 17264
rect 11572 17252 11578 17264
rect 13906 17252 13912 17264
rect 11572 17224 13912 17252
rect 11572 17212 11578 17224
rect 13906 17212 13912 17224
rect 13964 17252 13970 17264
rect 14544 17255 14602 17261
rect 13964 17224 14320 17252
rect 13964 17212 13970 17224
rect 12253 17187 12311 17193
rect 12253 17153 12265 17187
rect 12299 17184 12311 17187
rect 12710 17184 12716 17196
rect 12299 17156 12716 17184
rect 12299 17153 12311 17156
rect 12253 17147 12311 17153
rect 12710 17144 12716 17156
rect 12768 17144 12774 17196
rect 13170 17144 13176 17196
rect 13228 17184 13234 17196
rect 14292 17193 14320 17224
rect 14544 17221 14556 17255
rect 14590 17252 14602 17255
rect 15010 17252 15016 17264
rect 14590 17224 15016 17252
rect 14590 17221 14602 17224
rect 14544 17215 14602 17221
rect 15010 17212 15016 17224
rect 15068 17212 15074 17264
rect 18684 17255 18742 17261
rect 18684 17221 18696 17255
rect 18730 17252 18742 17255
rect 19426 17252 19432 17264
rect 18730 17224 19432 17252
rect 18730 17221 18742 17224
rect 18684 17215 18742 17221
rect 19426 17212 19432 17224
rect 19484 17212 19490 17264
rect 23284 17255 23342 17261
rect 23284 17221 23296 17255
rect 23330 17252 23342 17255
rect 23474 17252 23480 17264
rect 23330 17224 23480 17252
rect 23330 17221 23342 17224
rect 23284 17215 23342 17221
rect 23474 17212 23480 17224
rect 23532 17212 23538 17264
rect 30190 17212 30196 17264
rect 30248 17252 30254 17264
rect 33888 17261 33916 17292
rect 35805 17289 35817 17292
rect 35851 17289 35863 17323
rect 39114 17320 39120 17332
rect 35805 17283 35863 17289
rect 36556 17292 39120 17320
rect 33873 17255 33931 17261
rect 30248 17224 31340 17252
rect 30248 17212 30254 17224
rect 13449 17187 13507 17193
rect 13449 17184 13461 17187
rect 13228 17156 13461 17184
rect 13228 17144 13234 17156
rect 13449 17153 13461 17156
rect 13495 17153 13507 17187
rect 13449 17147 13507 17153
rect 14277 17187 14335 17193
rect 14277 17153 14289 17187
rect 14323 17153 14335 17187
rect 14277 17147 14335 17153
rect 17037 17187 17095 17193
rect 17037 17153 17049 17187
rect 17083 17184 17095 17187
rect 18322 17184 18328 17196
rect 17083 17156 18328 17184
rect 17083 17153 17095 17156
rect 17037 17147 17095 17153
rect 18322 17144 18328 17156
rect 18380 17144 18386 17196
rect 22186 17184 22192 17196
rect 22147 17156 22192 17184
rect 22186 17144 22192 17156
rect 22244 17144 22250 17196
rect 22465 17187 22523 17193
rect 22465 17153 22477 17187
rect 22511 17184 22523 17187
rect 22554 17184 22560 17196
rect 22511 17156 22560 17184
rect 22511 17153 22523 17156
rect 22465 17147 22523 17153
rect 22554 17144 22560 17156
rect 22612 17184 22618 17196
rect 23842 17184 23848 17196
rect 22612 17156 23848 17184
rect 22612 17144 22618 17156
rect 23842 17144 23848 17156
rect 23900 17144 23906 17196
rect 24394 17144 24400 17196
rect 24452 17184 24458 17196
rect 25225 17187 25283 17193
rect 25225 17184 25237 17187
rect 24452 17156 25237 17184
rect 24452 17144 24458 17156
rect 25225 17153 25237 17156
rect 25271 17153 25283 17187
rect 26142 17184 26148 17196
rect 25225 17147 25283 17153
rect 25516 17156 26148 17184
rect 13541 17119 13599 17125
rect 13541 17085 13553 17119
rect 13587 17085 13599 17119
rect 13541 17079 13599 17085
rect 13817 17119 13875 17125
rect 13817 17085 13829 17119
rect 13863 17116 13875 17119
rect 14090 17116 14096 17128
rect 13863 17088 14096 17116
rect 13863 17085 13875 17088
rect 13817 17079 13875 17085
rect 13556 17048 13584 17079
rect 14090 17076 14096 17088
rect 14148 17076 14154 17128
rect 18414 17116 18420 17128
rect 18375 17088 18420 17116
rect 18414 17076 18420 17088
rect 18472 17076 18478 17128
rect 23017 17119 23075 17125
rect 23017 17085 23029 17119
rect 23063 17085 23075 17119
rect 25314 17116 25320 17128
rect 25275 17088 25320 17116
rect 23017 17079 23075 17085
rect 13556 17020 14320 17048
rect 1578 16940 1584 16992
rect 1636 16980 1642 16992
rect 2317 16983 2375 16989
rect 2317 16980 2329 16983
rect 1636 16952 2329 16980
rect 1636 16940 1642 16952
rect 2317 16949 2329 16952
rect 2363 16949 2375 16983
rect 14292 16980 14320 17020
rect 22094 17008 22100 17060
rect 22152 17048 22158 17060
rect 22738 17048 22744 17060
rect 22152 17020 22744 17048
rect 22152 17008 22158 17020
rect 22738 17008 22744 17020
rect 22796 17048 22802 17060
rect 23032 17048 23060 17079
rect 25314 17076 25320 17088
rect 25372 17076 25378 17128
rect 25516 17125 25544 17156
rect 26142 17144 26148 17156
rect 26200 17144 26206 17196
rect 30742 17144 30748 17196
rect 30800 17184 30806 17196
rect 31312 17193 31340 17224
rect 33873 17221 33885 17255
rect 33919 17221 33931 17255
rect 34606 17252 34612 17264
rect 34567 17224 34612 17252
rect 33873 17215 33931 17221
rect 34606 17212 34612 17224
rect 34664 17212 34670 17264
rect 34790 17212 34796 17264
rect 34848 17261 34854 17264
rect 34848 17255 34867 17261
rect 34855 17221 34867 17255
rect 34848 17215 34867 17221
rect 35437 17255 35495 17261
rect 35437 17221 35449 17255
rect 35483 17221 35495 17255
rect 35437 17215 35495 17221
rect 34848 17212 34854 17215
rect 31021 17187 31079 17193
rect 31021 17184 31033 17187
rect 30800 17156 31033 17184
rect 30800 17144 30806 17156
rect 31021 17153 31033 17156
rect 31067 17153 31079 17187
rect 31021 17147 31079 17153
rect 31297 17187 31355 17193
rect 31297 17153 31309 17187
rect 31343 17153 31355 17187
rect 31297 17147 31355 17153
rect 31481 17187 31539 17193
rect 31481 17153 31493 17187
rect 31527 17153 31539 17187
rect 31481 17147 31539 17153
rect 25501 17119 25559 17125
rect 25501 17085 25513 17119
rect 25547 17085 25559 17119
rect 25501 17079 25559 17085
rect 30926 17076 30932 17128
rect 30984 17116 30990 17128
rect 31496 17116 31524 17147
rect 33318 17144 33324 17196
rect 33376 17184 33382 17196
rect 34057 17187 34115 17193
rect 34057 17184 34069 17187
rect 33376 17156 34069 17184
rect 33376 17144 33382 17156
rect 34057 17153 34069 17156
rect 34103 17153 34115 17187
rect 34057 17147 34115 17153
rect 34149 17187 34207 17193
rect 34149 17153 34161 17187
rect 34195 17184 34207 17187
rect 34514 17184 34520 17196
rect 34195 17156 34520 17184
rect 34195 17153 34207 17156
rect 34149 17147 34207 17153
rect 34514 17144 34520 17156
rect 34572 17144 34578 17196
rect 35452 17184 35480 17215
rect 35526 17212 35532 17264
rect 35584 17252 35590 17264
rect 35637 17255 35695 17261
rect 35637 17252 35649 17255
rect 35584 17224 35649 17252
rect 35584 17212 35590 17224
rect 35637 17221 35649 17224
rect 35683 17221 35695 17255
rect 35637 17215 35695 17221
rect 35986 17184 35992 17196
rect 35452 17156 35992 17184
rect 35986 17144 35992 17156
rect 36044 17184 36050 17196
rect 36556 17193 36584 17292
rect 39114 17280 39120 17292
rect 39172 17280 39178 17332
rect 41046 17280 41052 17332
rect 41104 17320 41110 17332
rect 41785 17323 41843 17329
rect 41785 17320 41797 17323
rect 41104 17292 41797 17320
rect 41104 17280 41110 17292
rect 41785 17289 41797 17292
rect 41831 17289 41843 17323
rect 41785 17283 41843 17289
rect 43438 17280 43444 17332
rect 43496 17320 43502 17332
rect 44913 17323 44971 17329
rect 44913 17320 44925 17323
rect 43496 17292 44925 17320
rect 43496 17280 43502 17292
rect 44913 17289 44925 17292
rect 44959 17289 44971 17323
rect 44913 17283 44971 17289
rect 37366 17212 37372 17264
rect 37424 17252 37430 17264
rect 39393 17255 39451 17261
rect 39393 17252 39405 17255
rect 37424 17224 39405 17252
rect 37424 17212 37430 17224
rect 39393 17221 39405 17224
rect 39439 17221 39451 17255
rect 44358 17252 44364 17264
rect 39393 17215 39451 17221
rect 43548 17224 44364 17252
rect 36541 17187 36599 17193
rect 36541 17184 36553 17187
rect 36044 17156 36553 17184
rect 36044 17144 36050 17156
rect 36541 17153 36553 17156
rect 36587 17153 36599 17187
rect 36541 17147 36599 17153
rect 36814 17144 36820 17196
rect 36872 17184 36878 17196
rect 37717 17187 37775 17193
rect 37717 17184 37729 17187
rect 36872 17156 37729 17184
rect 36872 17144 36878 17156
rect 37717 17153 37729 17156
rect 37763 17153 37775 17187
rect 37717 17147 37775 17153
rect 39301 17187 39359 17193
rect 39301 17153 39313 17187
rect 39347 17153 39359 17187
rect 39482 17184 39488 17196
rect 39443 17156 39488 17184
rect 39301 17147 39359 17153
rect 30984 17088 31524 17116
rect 30984 17076 30990 17088
rect 33686 17076 33692 17128
rect 33744 17116 33750 17128
rect 36633 17119 36691 17125
rect 33744 17088 35020 17116
rect 33744 17076 33750 17088
rect 22796 17020 23060 17048
rect 22796 17008 22802 17020
rect 26234 17008 26240 17060
rect 26292 17048 26298 17060
rect 27430 17048 27436 17060
rect 26292 17020 27436 17048
rect 26292 17008 26298 17020
rect 27430 17008 27436 17020
rect 27488 17048 27494 17060
rect 33410 17048 33416 17060
rect 27488 17020 33416 17048
rect 27488 17008 27494 17020
rect 33410 17008 33416 17020
rect 33468 17048 33474 17060
rect 33873 17051 33931 17057
rect 33468 17020 33732 17048
rect 33468 17008 33474 17020
rect 15010 16980 15016 16992
rect 14292 16952 15016 16980
rect 2317 16943 2375 16949
rect 15010 16940 15016 16952
rect 15068 16980 15074 16992
rect 15657 16983 15715 16989
rect 15657 16980 15669 16983
rect 15068 16952 15669 16980
rect 15068 16940 15074 16952
rect 15657 16949 15669 16952
rect 15703 16949 15715 16983
rect 16850 16980 16856 16992
rect 16811 16952 16856 16980
rect 15657 16943 15715 16949
rect 16850 16940 16856 16952
rect 16908 16940 16914 16992
rect 22002 16980 22008 16992
rect 21963 16952 22008 16980
rect 22002 16940 22008 16952
rect 22060 16940 22066 16992
rect 22373 16983 22431 16989
rect 22373 16949 22385 16983
rect 22419 16980 22431 16983
rect 22554 16980 22560 16992
rect 22419 16952 22560 16980
rect 22419 16949 22431 16952
rect 22373 16943 22431 16949
rect 22554 16940 22560 16952
rect 22612 16940 22618 16992
rect 24394 16980 24400 16992
rect 24355 16952 24400 16980
rect 24394 16940 24400 16952
rect 24452 16940 24458 16992
rect 24854 16980 24860 16992
rect 24815 16952 24860 16980
rect 24854 16940 24860 16952
rect 24912 16940 24918 16992
rect 30837 16983 30895 16989
rect 30837 16949 30849 16983
rect 30883 16980 30895 16983
rect 32490 16980 32496 16992
rect 30883 16952 32496 16980
rect 30883 16949 30895 16952
rect 30837 16943 30895 16949
rect 32490 16940 32496 16952
rect 32548 16940 32554 16992
rect 33704 16980 33732 17020
rect 33873 17017 33885 17051
rect 33919 17048 33931 17051
rect 34054 17048 34060 17060
rect 33919 17020 34060 17048
rect 33919 17017 33931 17020
rect 33873 17011 33931 17017
rect 34054 17008 34060 17020
rect 34112 17008 34118 17060
rect 34422 16980 34428 16992
rect 33704 16952 34428 16980
rect 34422 16940 34428 16952
rect 34480 16940 34486 16992
rect 34698 16940 34704 16992
rect 34756 16980 34762 16992
rect 34992 16989 35020 17088
rect 36633 17085 36645 17119
rect 36679 17085 36691 17119
rect 36906 17116 36912 17128
rect 36867 17088 36912 17116
rect 36633 17079 36691 17085
rect 34793 16983 34851 16989
rect 34793 16980 34805 16983
rect 34756 16952 34805 16980
rect 34756 16940 34762 16952
rect 34793 16949 34805 16952
rect 34839 16949 34851 16983
rect 34793 16943 34851 16949
rect 34977 16983 35035 16989
rect 34977 16949 34989 16983
rect 35023 16949 35035 16983
rect 34977 16943 35035 16949
rect 35621 16983 35679 16989
rect 35621 16949 35633 16983
rect 35667 16980 35679 16983
rect 35802 16980 35808 16992
rect 35667 16952 35808 16980
rect 35667 16949 35679 16952
rect 35621 16943 35679 16949
rect 35802 16940 35808 16952
rect 35860 16980 35866 16992
rect 36648 16980 36676 17079
rect 36906 17076 36912 17088
rect 36964 17076 36970 17128
rect 37458 17116 37464 17128
rect 37419 17088 37464 17116
rect 37458 17076 37464 17088
rect 37516 17076 37522 17128
rect 39316 17116 39344 17147
rect 39482 17144 39488 17156
rect 39540 17144 39546 17196
rect 41598 17184 41604 17196
rect 41559 17156 41604 17184
rect 41598 17144 41604 17156
rect 41656 17144 41662 17196
rect 42705 17187 42763 17193
rect 42705 17153 42717 17187
rect 42751 17184 42763 17187
rect 42886 17184 42892 17196
rect 42751 17156 42892 17184
rect 42751 17153 42763 17156
rect 42705 17147 42763 17153
rect 42886 17144 42892 17156
rect 42944 17144 42950 17196
rect 43548 17193 43576 17224
rect 44358 17212 44364 17224
rect 44416 17212 44422 17264
rect 45557 17255 45615 17261
rect 45557 17221 45569 17255
rect 45603 17252 45615 17255
rect 47118 17252 47124 17264
rect 45603 17224 47124 17252
rect 45603 17221 45615 17224
rect 45557 17215 45615 17221
rect 47118 17212 47124 17224
rect 47176 17212 47182 17264
rect 43533 17187 43591 17193
rect 43533 17153 43545 17187
rect 43579 17153 43591 17187
rect 43533 17147 43591 17153
rect 39942 17116 39948 17128
rect 39316 17088 39948 17116
rect 39942 17076 39948 17088
rect 40000 17076 40006 17128
rect 41417 17119 41475 17125
rect 41417 17085 41429 17119
rect 41463 17116 41475 17119
rect 43254 17116 43260 17128
rect 41463 17088 43260 17116
rect 41463 17085 41475 17088
rect 41417 17079 41475 17085
rect 43254 17076 43260 17088
rect 43312 17076 43318 17128
rect 42702 17008 42708 17060
rect 42760 17048 42766 17060
rect 43548 17048 43576 17147
rect 43622 17144 43628 17196
rect 43680 17184 43686 17196
rect 43789 17187 43847 17193
rect 43789 17184 43801 17187
rect 43680 17156 43801 17184
rect 43680 17144 43686 17156
rect 43789 17153 43801 17156
rect 43835 17153 43847 17187
rect 43789 17147 43847 17153
rect 45373 17119 45431 17125
rect 45373 17085 45385 17119
rect 45419 17116 45431 17119
rect 46382 17116 46388 17128
rect 45419 17088 46388 17116
rect 45419 17085 45431 17088
rect 45373 17079 45431 17085
rect 46382 17076 46388 17088
rect 46440 17076 46446 17128
rect 46842 17116 46848 17128
rect 46803 17088 46848 17116
rect 46842 17076 46848 17088
rect 46900 17076 46906 17128
rect 42760 17020 43576 17048
rect 42760 17008 42766 17020
rect 37642 16980 37648 16992
rect 35860 16952 37648 16980
rect 35860 16940 35866 16952
rect 37642 16940 37648 16952
rect 37700 16980 37706 16992
rect 38841 16983 38899 16989
rect 38841 16980 38853 16983
rect 37700 16952 38853 16980
rect 37700 16940 37706 16952
rect 38841 16949 38853 16952
rect 38887 16949 38899 16983
rect 38841 16943 38899 16949
rect 42981 16983 43039 16989
rect 42981 16949 42993 16983
rect 43027 16980 43039 16983
rect 43806 16980 43812 16992
rect 43027 16952 43812 16980
rect 43027 16949 43039 16952
rect 42981 16943 43039 16949
rect 43806 16940 43812 16952
rect 43864 16980 43870 16992
rect 44174 16980 44180 16992
rect 43864 16952 44180 16980
rect 43864 16940 43870 16952
rect 44174 16940 44180 16952
rect 44232 16940 44238 16992
rect 46474 16940 46480 16992
rect 46532 16980 46538 16992
rect 47949 16983 48007 16989
rect 47949 16980 47961 16983
rect 46532 16952 47961 16980
rect 46532 16940 46538 16952
rect 47949 16949 47961 16952
rect 47995 16949 48007 16983
rect 47949 16943 48007 16949
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 12710 16776 12716 16788
rect 12671 16748 12716 16776
rect 12710 16736 12716 16748
rect 12768 16736 12774 16788
rect 16758 16776 16764 16788
rect 16408 16748 16764 16776
rect 1578 16640 1584 16652
rect 1539 16612 1584 16640
rect 1578 16600 1584 16612
rect 1636 16600 1642 16652
rect 2774 16640 2780 16652
rect 2735 16612 2780 16640
rect 2774 16600 2780 16612
rect 2832 16600 2838 16652
rect 13170 16640 13176 16652
rect 13131 16612 13176 16640
rect 13170 16600 13176 16612
rect 13228 16600 13234 16652
rect 13354 16640 13360 16652
rect 13315 16612 13360 16640
rect 13354 16600 13360 16612
rect 13412 16600 13418 16652
rect 16408 16649 16436 16748
rect 16758 16736 16764 16748
rect 16816 16736 16822 16788
rect 22094 16776 22100 16788
rect 20824 16748 22100 16776
rect 18414 16668 18420 16720
rect 18472 16668 18478 16720
rect 16393 16643 16451 16649
rect 16393 16609 16405 16643
rect 16439 16609 16451 16643
rect 18432 16640 18460 16668
rect 20824 16649 20852 16748
rect 22094 16736 22100 16748
rect 22152 16736 22158 16788
rect 23474 16776 23480 16788
rect 23435 16748 23480 16776
rect 23474 16736 23480 16748
rect 23532 16736 23538 16788
rect 26142 16736 26148 16788
rect 26200 16776 26206 16788
rect 26237 16779 26295 16785
rect 26237 16776 26249 16779
rect 26200 16748 26249 16776
rect 26200 16736 26206 16748
rect 26237 16745 26249 16748
rect 26283 16745 26295 16779
rect 26237 16739 26295 16745
rect 27614 16736 27620 16788
rect 27672 16776 27678 16788
rect 27801 16779 27859 16785
rect 27801 16776 27813 16779
rect 27672 16748 27813 16776
rect 27672 16736 27678 16748
rect 27801 16745 27813 16748
rect 27847 16745 27859 16779
rect 27801 16739 27859 16745
rect 30282 16736 30288 16788
rect 30340 16776 30346 16788
rect 30340 16748 31754 16776
rect 30340 16736 30346 16748
rect 26326 16708 26332 16720
rect 25056 16680 26332 16708
rect 20809 16643 20867 16649
rect 20809 16640 20821 16643
rect 18432 16612 20821 16640
rect 16393 16603 16451 16609
rect 20809 16609 20821 16612
rect 20855 16609 20867 16643
rect 20809 16603 20867 16609
rect 24486 16600 24492 16652
rect 24544 16640 24550 16652
rect 25056 16649 25084 16680
rect 26326 16668 26332 16680
rect 26384 16668 26390 16720
rect 25041 16643 25099 16649
rect 24544 16612 24992 16640
rect 24544 16600 24550 16612
rect 21076 16575 21134 16581
rect 21076 16541 21088 16575
rect 21122 16572 21134 16575
rect 22002 16572 22008 16584
rect 21122 16544 22008 16572
rect 21122 16541 21134 16544
rect 21076 16535 21134 16541
rect 22002 16532 22008 16544
rect 22060 16532 22066 16584
rect 23661 16575 23719 16581
rect 23661 16541 23673 16575
rect 23707 16572 23719 16575
rect 24854 16572 24860 16584
rect 23707 16544 24860 16572
rect 23707 16541 23719 16544
rect 23661 16535 23719 16541
rect 24854 16532 24860 16544
rect 24912 16532 24918 16584
rect 24964 16572 24992 16612
rect 25041 16609 25053 16643
rect 25087 16609 25099 16643
rect 25222 16640 25228 16652
rect 25183 16612 25228 16640
rect 25041 16603 25099 16609
rect 25222 16600 25228 16612
rect 25280 16640 25286 16652
rect 25774 16640 25780 16652
rect 25280 16612 25780 16640
rect 25280 16600 25286 16612
rect 25774 16600 25780 16612
rect 25832 16600 25838 16652
rect 25958 16600 25964 16652
rect 26016 16640 26022 16652
rect 26881 16643 26939 16649
rect 26881 16640 26893 16643
rect 26016 16612 26893 16640
rect 26016 16600 26022 16612
rect 26881 16609 26893 16612
rect 26927 16609 26939 16643
rect 27893 16643 27951 16649
rect 27893 16640 27905 16643
rect 26881 16603 26939 16609
rect 27356 16612 27905 16640
rect 27356 16584 27384 16612
rect 27893 16609 27905 16612
rect 27939 16609 27951 16643
rect 30282 16640 30288 16652
rect 30243 16612 30288 16640
rect 27893 16603 27951 16609
rect 30282 16600 30288 16612
rect 30340 16600 30346 16652
rect 31726 16640 31754 16748
rect 34698 16736 34704 16788
rect 34756 16776 34762 16788
rect 35253 16779 35311 16785
rect 35253 16776 35265 16779
rect 34756 16748 35265 16776
rect 34756 16736 34762 16748
rect 35253 16745 35265 16748
rect 35299 16776 35311 16779
rect 35526 16776 35532 16788
rect 35299 16748 35532 16776
rect 35299 16745 35311 16748
rect 35253 16739 35311 16745
rect 35526 16736 35532 16748
rect 35584 16736 35590 16788
rect 36722 16776 36728 16788
rect 36683 16748 36728 16776
rect 36722 16736 36728 16748
rect 36780 16736 36786 16788
rect 36814 16736 36820 16788
rect 36872 16776 36878 16788
rect 43441 16779 43499 16785
rect 36872 16748 36917 16776
rect 36872 16736 36878 16748
rect 43441 16745 43453 16779
rect 43487 16776 43499 16779
rect 43622 16776 43628 16788
rect 43487 16748 43628 16776
rect 43487 16745 43499 16748
rect 43441 16739 43499 16745
rect 43622 16736 43628 16748
rect 43680 16736 43686 16788
rect 33318 16668 33324 16720
rect 33376 16708 33382 16720
rect 35066 16708 35072 16720
rect 33376 16680 35072 16708
rect 33376 16668 33382 16680
rect 35066 16668 35072 16680
rect 35124 16708 35130 16720
rect 38286 16708 38292 16720
rect 35124 16680 35940 16708
rect 38199 16680 38292 16708
rect 35124 16668 35130 16680
rect 32125 16643 32183 16649
rect 32125 16640 32137 16643
rect 31726 16612 32137 16640
rect 32125 16609 32137 16612
rect 32171 16609 32183 16643
rect 35342 16640 35348 16652
rect 32125 16603 32183 16609
rect 34256 16612 35348 16640
rect 25869 16575 25927 16581
rect 24964 16544 25452 16572
rect 1765 16507 1823 16513
rect 1765 16473 1777 16507
rect 1811 16504 1823 16507
rect 2590 16504 2596 16516
rect 1811 16476 2596 16504
rect 1811 16473 1823 16476
rect 1765 16467 1823 16473
rect 2590 16464 2596 16476
rect 2648 16464 2654 16516
rect 16660 16507 16718 16513
rect 16660 16473 16672 16507
rect 16706 16504 16718 16507
rect 16850 16504 16856 16516
rect 16706 16476 16856 16504
rect 16706 16473 16718 16476
rect 16660 16467 16718 16473
rect 16850 16464 16856 16476
rect 16908 16464 16914 16516
rect 25314 16504 25320 16516
rect 24596 16476 25320 16504
rect 13081 16439 13139 16445
rect 13081 16405 13093 16439
rect 13127 16436 13139 16439
rect 17494 16436 17500 16448
rect 13127 16408 17500 16436
rect 13127 16405 13139 16408
rect 13081 16399 13139 16405
rect 17494 16396 17500 16408
rect 17552 16436 17558 16448
rect 17773 16439 17831 16445
rect 17773 16436 17785 16439
rect 17552 16408 17785 16436
rect 17552 16396 17558 16408
rect 17773 16405 17785 16408
rect 17819 16405 17831 16439
rect 17773 16399 17831 16405
rect 22189 16439 22247 16445
rect 22189 16405 22201 16439
rect 22235 16436 22247 16439
rect 22646 16436 22652 16448
rect 22235 16408 22652 16436
rect 22235 16405 22247 16408
rect 22189 16399 22247 16405
rect 22646 16396 22652 16408
rect 22704 16396 22710 16448
rect 24596 16445 24624 16476
rect 25314 16464 25320 16476
rect 25372 16464 25378 16516
rect 24581 16439 24639 16445
rect 24581 16405 24593 16439
rect 24627 16405 24639 16439
rect 24946 16436 24952 16448
rect 24907 16408 24952 16436
rect 24581 16399 24639 16405
rect 24946 16396 24952 16408
rect 25004 16396 25010 16448
rect 25424 16436 25452 16544
rect 25869 16541 25881 16575
rect 25915 16572 25927 16575
rect 26694 16572 26700 16584
rect 25915 16544 26700 16572
rect 25915 16541 25927 16544
rect 25869 16535 25927 16541
rect 26694 16532 26700 16544
rect 26752 16532 26758 16584
rect 27062 16572 27068 16584
rect 27023 16544 27068 16572
rect 27062 16532 27068 16544
rect 27120 16532 27126 16584
rect 27246 16572 27252 16584
rect 27207 16544 27252 16572
rect 27246 16532 27252 16544
rect 27304 16532 27310 16584
rect 27338 16532 27344 16584
rect 27396 16572 27402 16584
rect 27801 16575 27859 16581
rect 27396 16544 27441 16572
rect 27396 16532 27402 16544
rect 27801 16541 27813 16575
rect 27847 16541 27859 16575
rect 27801 16535 27859 16541
rect 34057 16575 34115 16581
rect 34057 16541 34069 16575
rect 34103 16572 34115 16575
rect 34256 16572 34284 16612
rect 35342 16600 35348 16612
rect 35400 16600 35406 16652
rect 34103 16544 34284 16572
rect 34333 16575 34391 16581
rect 34103 16541 34115 16544
rect 34057 16535 34115 16541
rect 34333 16541 34345 16575
rect 34379 16572 34391 16575
rect 34790 16572 34796 16584
rect 34379 16544 34796 16572
rect 34379 16541 34391 16544
rect 34333 16535 34391 16541
rect 26050 16464 26056 16516
rect 26108 16504 26114 16516
rect 26418 16504 26424 16516
rect 26108 16476 26424 16504
rect 26108 16464 26114 16476
rect 26418 16464 26424 16476
rect 26476 16464 26482 16516
rect 26510 16464 26516 16516
rect 26568 16504 26574 16516
rect 27816 16504 27844 16535
rect 34790 16532 34796 16544
rect 34848 16572 34854 16584
rect 35710 16572 35716 16584
rect 34848 16544 35204 16572
rect 35671 16544 35716 16572
rect 34848 16532 34854 16544
rect 28258 16504 28264 16516
rect 26568 16476 27844 16504
rect 27908 16476 28264 16504
rect 26568 16464 26574 16476
rect 27908 16436 27936 16476
rect 28258 16464 28264 16476
rect 28316 16464 28322 16516
rect 30558 16513 30564 16516
rect 30552 16467 30564 16513
rect 30616 16504 30622 16516
rect 32398 16513 32404 16516
rect 30616 16476 30652 16504
rect 30558 16464 30564 16467
rect 30616 16464 30622 16476
rect 32392 16467 32404 16513
rect 32456 16504 32462 16516
rect 34241 16507 34299 16513
rect 32456 16476 32492 16504
rect 32398 16464 32404 16467
rect 32456 16464 32462 16476
rect 34241 16473 34253 16507
rect 34287 16504 34299 16507
rect 34698 16504 34704 16516
rect 34287 16476 34704 16504
rect 34287 16473 34299 16476
rect 34241 16467 34299 16473
rect 34698 16464 34704 16476
rect 34756 16464 34762 16516
rect 34885 16507 34943 16513
rect 34885 16473 34897 16507
rect 34931 16473 34943 16507
rect 35066 16504 35072 16516
rect 35027 16476 35072 16504
rect 34885 16467 34943 16473
rect 28166 16436 28172 16448
rect 25424 16408 27936 16436
rect 28127 16408 28172 16436
rect 28166 16396 28172 16408
rect 28224 16396 28230 16448
rect 31478 16396 31484 16448
rect 31536 16436 31542 16448
rect 31665 16439 31723 16445
rect 31665 16436 31677 16439
rect 31536 16408 31677 16436
rect 31536 16396 31542 16408
rect 31665 16405 31677 16408
rect 31711 16405 31723 16439
rect 31665 16399 31723 16405
rect 33318 16396 33324 16448
rect 33376 16436 33382 16448
rect 33505 16439 33563 16445
rect 33505 16436 33517 16439
rect 33376 16408 33517 16436
rect 33376 16396 33382 16408
rect 33505 16405 33517 16408
rect 33551 16405 33563 16439
rect 34146 16436 34152 16448
rect 34204 16445 34210 16448
rect 34113 16408 34152 16436
rect 33505 16399 33563 16405
rect 34146 16396 34152 16408
rect 34204 16399 34213 16445
rect 34204 16396 34210 16399
rect 34514 16396 34520 16448
rect 34572 16436 34578 16448
rect 34900 16436 34928 16467
rect 35066 16464 35072 16476
rect 35124 16464 35130 16516
rect 35176 16504 35204 16544
rect 35710 16532 35716 16544
rect 35768 16532 35774 16584
rect 35912 16581 35940 16680
rect 38286 16668 38292 16680
rect 38344 16708 38350 16720
rect 44542 16708 44548 16720
rect 38344 16680 44548 16708
rect 38344 16668 38350 16680
rect 44542 16668 44548 16680
rect 44600 16668 44606 16720
rect 36909 16643 36967 16649
rect 36909 16609 36921 16643
rect 36955 16640 36967 16643
rect 37274 16640 37280 16652
rect 36955 16612 37280 16640
rect 36955 16609 36967 16612
rect 36909 16603 36967 16609
rect 37274 16600 37280 16612
rect 37332 16600 37338 16652
rect 37458 16600 37464 16652
rect 37516 16640 37522 16652
rect 40402 16640 40408 16652
rect 37516 16612 40408 16640
rect 37516 16600 37522 16612
rect 40402 16600 40408 16612
rect 40460 16640 40466 16652
rect 40770 16640 40776 16652
rect 40460 16612 40776 16640
rect 40460 16600 40466 16612
rect 40770 16600 40776 16612
rect 40828 16600 40834 16652
rect 41782 16640 41788 16652
rect 40880 16612 41788 16640
rect 35897 16575 35955 16581
rect 35897 16541 35909 16575
rect 35943 16541 35955 16575
rect 36630 16572 36636 16584
rect 36591 16544 36636 16572
rect 35897 16535 35955 16541
rect 36630 16532 36636 16544
rect 36688 16532 36694 16584
rect 37366 16532 37372 16584
rect 37424 16572 37430 16584
rect 38013 16575 38071 16581
rect 38013 16572 38025 16575
rect 37424 16544 38025 16572
rect 37424 16532 37430 16544
rect 38013 16541 38025 16544
rect 38059 16541 38071 16575
rect 38013 16535 38071 16541
rect 39482 16532 39488 16584
rect 39540 16572 39546 16584
rect 40880 16572 40908 16612
rect 41782 16600 41788 16612
rect 41840 16600 41846 16652
rect 46474 16640 46480 16652
rect 46435 16612 46480 16640
rect 46474 16600 46480 16612
rect 46532 16600 46538 16652
rect 48222 16640 48228 16652
rect 48183 16612 48228 16640
rect 48222 16600 48228 16612
rect 48280 16600 48286 16652
rect 39540 16544 40908 16572
rect 39540 16532 39546 16544
rect 42794 16532 42800 16584
rect 42852 16572 42858 16584
rect 43625 16575 43683 16581
rect 43625 16572 43637 16575
rect 42852 16544 43637 16572
rect 42852 16532 42858 16544
rect 43625 16541 43637 16544
rect 43671 16541 43683 16575
rect 43625 16535 43683 16541
rect 35805 16507 35863 16513
rect 35805 16504 35817 16507
rect 35176 16476 35817 16504
rect 35805 16473 35817 16476
rect 35851 16473 35863 16507
rect 35805 16467 35863 16473
rect 46661 16507 46719 16513
rect 46661 16473 46673 16507
rect 46707 16504 46719 16507
rect 46750 16504 46756 16516
rect 46707 16476 46756 16504
rect 46707 16473 46719 16476
rect 46661 16467 46719 16473
rect 46750 16464 46756 16476
rect 46808 16464 46814 16516
rect 35710 16436 35716 16448
rect 34572 16408 35716 16436
rect 34572 16396 34578 16408
rect 35710 16396 35716 16408
rect 35768 16396 35774 16448
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 2590 16232 2596 16244
rect 2551 16204 2596 16232
rect 2590 16192 2596 16204
rect 2648 16192 2654 16244
rect 13170 16192 13176 16244
rect 13228 16232 13234 16244
rect 13449 16235 13507 16241
rect 13449 16232 13461 16235
rect 13228 16204 13461 16232
rect 13228 16192 13234 16204
rect 13449 16201 13461 16204
rect 13495 16201 13507 16235
rect 13449 16195 13507 16201
rect 17129 16235 17187 16241
rect 17129 16201 17141 16235
rect 17175 16201 17187 16235
rect 17494 16232 17500 16244
rect 17455 16204 17500 16232
rect 17129 16195 17187 16201
rect 14737 16167 14795 16173
rect 14737 16133 14749 16167
rect 14783 16164 14795 16167
rect 17034 16164 17040 16176
rect 14783 16136 17040 16164
rect 14783 16133 14795 16136
rect 14737 16127 14795 16133
rect 17034 16124 17040 16136
rect 17092 16124 17098 16176
rect 17144 16164 17172 16195
rect 17494 16192 17500 16204
rect 17552 16192 17558 16244
rect 18414 16192 18420 16244
rect 18472 16232 18478 16244
rect 18693 16235 18751 16241
rect 18693 16232 18705 16235
rect 18472 16204 18705 16232
rect 18472 16192 18478 16204
rect 18693 16201 18705 16204
rect 18739 16201 18751 16235
rect 18693 16195 18751 16201
rect 22005 16235 22063 16241
rect 22005 16201 22017 16235
rect 22051 16232 22063 16235
rect 22186 16232 22192 16244
rect 22051 16204 22192 16232
rect 22051 16201 22063 16204
rect 22005 16195 22063 16201
rect 22186 16192 22192 16204
rect 22244 16192 22250 16244
rect 26237 16235 26295 16241
rect 26237 16201 26249 16235
rect 26283 16232 26295 16235
rect 26326 16232 26332 16244
rect 26283 16204 26332 16232
rect 26283 16201 26295 16204
rect 26237 16195 26295 16201
rect 26326 16192 26332 16204
rect 26384 16192 26390 16244
rect 26418 16192 26424 16244
rect 26476 16232 26482 16244
rect 32309 16235 32367 16241
rect 26476 16204 31754 16232
rect 26476 16192 26482 16204
rect 18325 16167 18383 16173
rect 18325 16164 18337 16167
rect 17144 16136 18337 16164
rect 18325 16133 18337 16136
rect 18371 16133 18383 16167
rect 24946 16164 24952 16176
rect 18325 16127 18383 16133
rect 23299 16136 24952 16164
rect 2406 16056 2412 16108
rect 2464 16096 2470 16108
rect 2501 16099 2559 16105
rect 2501 16096 2513 16099
rect 2464 16068 2513 16096
rect 2464 16056 2470 16068
rect 2501 16065 2513 16068
rect 2547 16065 2559 16099
rect 2501 16059 2559 16065
rect 12069 16099 12127 16105
rect 12069 16065 12081 16099
rect 12115 16096 12127 16099
rect 12158 16096 12164 16108
rect 12115 16068 12164 16096
rect 12115 16065 12127 16068
rect 12069 16059 12127 16065
rect 12158 16056 12164 16068
rect 12216 16056 12222 16108
rect 12336 16099 12394 16105
rect 12336 16065 12348 16099
rect 12382 16096 12394 16099
rect 12894 16096 12900 16108
rect 12382 16068 12900 16096
rect 12382 16065 12394 16068
rect 12336 16059 12394 16065
rect 12894 16056 12900 16068
rect 12952 16056 12958 16108
rect 14829 16099 14887 16105
rect 14829 16065 14841 16099
rect 14875 16096 14887 16099
rect 15194 16096 15200 16108
rect 14875 16068 15200 16096
rect 14875 16065 14887 16068
rect 14829 16059 14887 16065
rect 15194 16056 15200 16068
rect 15252 16056 15258 16108
rect 18509 16099 18567 16105
rect 18509 16065 18521 16099
rect 18555 16096 18567 16099
rect 18598 16096 18604 16108
rect 18555 16068 18604 16096
rect 18555 16065 18567 16068
rect 18509 16059 18567 16065
rect 18598 16056 18604 16068
rect 18656 16056 18662 16108
rect 18874 16056 18880 16108
rect 18932 16096 18938 16108
rect 19337 16099 19395 16105
rect 19337 16096 19349 16099
rect 18932 16068 19349 16096
rect 18932 16056 18938 16068
rect 19337 16065 19349 16068
rect 19383 16065 19395 16099
rect 22186 16096 22192 16108
rect 22147 16068 22192 16096
rect 19337 16059 19395 16065
rect 22186 16056 22192 16068
rect 22244 16056 22250 16108
rect 22462 16096 22468 16108
rect 22423 16068 22468 16096
rect 22462 16056 22468 16068
rect 22520 16056 22526 16108
rect 22646 16056 22652 16108
rect 22704 16096 22710 16108
rect 23299 16096 23327 16136
rect 24946 16124 24952 16136
rect 25004 16124 25010 16176
rect 25133 16167 25191 16173
rect 25133 16133 25145 16167
rect 25179 16164 25191 16167
rect 28166 16164 28172 16176
rect 25179 16136 27292 16164
rect 25179 16133 25191 16136
rect 25133 16127 25191 16133
rect 24394 16096 24400 16108
rect 22704 16068 23327 16096
rect 24307 16068 24400 16096
rect 22704 16056 22710 16068
rect 24394 16056 24400 16068
rect 24452 16056 24458 16108
rect 24578 16096 24584 16108
rect 24539 16068 24584 16096
rect 24578 16056 24584 16068
rect 24636 16056 24642 16108
rect 24762 16056 24768 16108
rect 24820 16096 24826 16108
rect 25041 16099 25099 16105
rect 25041 16096 25053 16099
rect 24820 16068 25053 16096
rect 24820 16056 24826 16068
rect 25041 16065 25053 16068
rect 25087 16065 25099 16099
rect 25041 16059 25099 16065
rect 25225 16099 25283 16105
rect 25225 16065 25237 16099
rect 25271 16065 25283 16099
rect 25225 16059 25283 16065
rect 25869 16099 25927 16105
rect 25869 16065 25881 16099
rect 25915 16096 25927 16099
rect 26234 16096 26240 16108
rect 25915 16068 26240 16096
rect 25915 16065 25927 16068
rect 25869 16059 25927 16065
rect 13354 15988 13360 16040
rect 13412 16028 13418 16040
rect 14921 16031 14979 16037
rect 14921 16028 14933 16031
rect 13412 16000 14933 16028
rect 13412 15988 13418 16000
rect 14921 15997 14933 16000
rect 14967 16028 14979 16031
rect 15102 16028 15108 16040
rect 14967 16000 15108 16028
rect 14967 15997 14979 16000
rect 14921 15991 14979 15997
rect 15102 15988 15108 16000
rect 15160 15988 15166 16040
rect 17586 16028 17592 16040
rect 17547 16000 17592 16028
rect 17586 15988 17592 16000
rect 17644 15988 17650 16040
rect 17678 15988 17684 16040
rect 17736 16028 17742 16040
rect 17736 16000 17781 16028
rect 17736 15988 17742 16000
rect 24412 15960 24440 16056
rect 24596 16028 24624 16056
rect 25240 16028 25268 16059
rect 26234 16056 26240 16068
rect 26292 16056 26298 16108
rect 27264 16105 27292 16136
rect 27448 16136 28172 16164
rect 27448 16105 27476 16136
rect 28166 16124 28172 16136
rect 28224 16124 28230 16176
rect 31386 16164 31392 16176
rect 31312 16136 31392 16164
rect 27249 16099 27307 16105
rect 27249 16065 27261 16099
rect 27295 16065 27307 16099
rect 27249 16059 27307 16065
rect 27433 16099 27491 16105
rect 27433 16065 27445 16099
rect 27479 16065 27491 16099
rect 27433 16059 27491 16065
rect 27522 16056 27528 16108
rect 27580 16096 27586 16108
rect 27801 16099 27859 16105
rect 27580 16068 27625 16096
rect 27580 16056 27586 16068
rect 27801 16065 27813 16099
rect 27847 16065 27859 16099
rect 31018 16096 31024 16108
rect 30979 16068 31024 16096
rect 27801 16059 27859 16065
rect 25958 16028 25964 16040
rect 24596 16000 25268 16028
rect 25919 16000 25964 16028
rect 25958 15988 25964 16000
rect 26016 15988 26022 16040
rect 27614 16028 27620 16040
rect 26436 16000 27620 16028
rect 24762 15960 24768 15972
rect 24412 15932 24768 15960
rect 24762 15920 24768 15932
rect 24820 15920 24826 15972
rect 26436 15904 26464 16000
rect 27614 15988 27620 16000
rect 27672 15988 27678 16040
rect 27062 15920 27068 15972
rect 27120 15960 27126 15972
rect 27816 15960 27844 16059
rect 31018 16056 31024 16068
rect 31076 16056 31082 16108
rect 31312 16105 31340 16136
rect 31386 16124 31392 16136
rect 31444 16124 31450 16176
rect 31726 16164 31754 16204
rect 32309 16201 32321 16235
rect 32355 16232 32367 16235
rect 32398 16232 32404 16244
rect 32355 16204 32404 16232
rect 32355 16201 32367 16204
rect 32309 16195 32367 16201
rect 32398 16192 32404 16204
rect 32456 16192 32462 16244
rect 34911 16235 34969 16241
rect 34532 16204 34836 16232
rect 34532 16164 34560 16204
rect 34698 16164 34704 16176
rect 31726 16136 34560 16164
rect 34659 16136 34704 16164
rect 34698 16124 34704 16136
rect 34756 16124 34762 16176
rect 34808 16164 34836 16204
rect 34911 16201 34923 16235
rect 34957 16232 34969 16235
rect 35342 16232 35348 16244
rect 34957 16204 35348 16232
rect 34957 16201 34969 16204
rect 34911 16195 34969 16201
rect 35342 16192 35348 16204
rect 35400 16192 35406 16244
rect 41598 16192 41604 16244
rect 41656 16232 41662 16244
rect 42813 16235 42871 16241
rect 42813 16232 42825 16235
rect 41656 16204 42825 16232
rect 41656 16192 41662 16204
rect 42813 16201 42825 16204
rect 42859 16201 42871 16235
rect 47118 16232 47124 16244
rect 47079 16204 47124 16232
rect 42813 16195 42871 16201
rect 47118 16192 47124 16204
rect 47176 16192 47182 16244
rect 39482 16164 39488 16176
rect 34808 16136 39488 16164
rect 39482 16124 39488 16136
rect 39540 16124 39546 16176
rect 41874 16164 41880 16176
rect 41386 16136 41880 16164
rect 31297 16099 31355 16105
rect 31297 16065 31309 16099
rect 31343 16065 31355 16099
rect 31478 16096 31484 16108
rect 31439 16068 31484 16096
rect 31297 16059 31355 16065
rect 31478 16056 31484 16068
rect 31536 16096 31542 16108
rect 32490 16096 32496 16108
rect 31536 16068 31754 16096
rect 32451 16068 32496 16096
rect 31536 16056 31542 16068
rect 27982 16028 27988 16040
rect 27943 16000 27988 16028
rect 27982 15988 27988 16000
rect 28040 15988 28046 16040
rect 30466 15960 30472 15972
rect 27120 15932 27844 15960
rect 27908 15932 30472 15960
rect 27120 15920 27126 15932
rect 13078 15852 13084 15904
rect 13136 15892 13142 15904
rect 14369 15895 14427 15901
rect 14369 15892 14381 15895
rect 13136 15864 14381 15892
rect 13136 15852 13142 15864
rect 14369 15861 14381 15864
rect 14415 15861 14427 15895
rect 19150 15892 19156 15904
rect 19111 15864 19156 15892
rect 14369 15855 14427 15861
rect 19150 15852 19156 15864
rect 19208 15852 19214 15904
rect 24397 15895 24455 15901
rect 24397 15861 24409 15895
rect 24443 15892 24455 15895
rect 26418 15892 26424 15904
rect 24443 15864 26424 15892
rect 24443 15861 24455 15864
rect 24397 15855 24455 15861
rect 26418 15852 26424 15864
rect 26476 15852 26482 15904
rect 26786 15852 26792 15904
rect 26844 15892 26850 15904
rect 27908 15892 27936 15932
rect 30466 15920 30472 15932
rect 30524 15920 30530 15972
rect 31726 15960 31754 16068
rect 32490 16056 32496 16068
rect 32548 16056 32554 16108
rect 32674 16096 32680 16108
rect 32635 16068 32680 16096
rect 32674 16056 32680 16068
rect 32732 16056 32738 16108
rect 32769 16099 32827 16105
rect 32769 16065 32781 16099
rect 32815 16096 32827 16099
rect 33318 16096 33324 16108
rect 32815 16068 33324 16096
rect 32815 16065 32827 16068
rect 32769 16059 32827 16065
rect 33318 16056 33324 16068
rect 33376 16056 33382 16108
rect 33410 16056 33416 16108
rect 33468 16096 33474 16108
rect 33468 16068 33513 16096
rect 33468 16056 33474 16068
rect 33594 16056 33600 16108
rect 33652 16096 33658 16108
rect 33652 16068 34100 16096
rect 33652 16056 33658 16068
rect 33689 16031 33747 16037
rect 33689 15997 33701 16031
rect 33735 15997 33747 16031
rect 34072 16028 34100 16068
rect 34146 16056 34152 16108
rect 34204 16096 34210 16108
rect 35529 16099 35587 16105
rect 35529 16096 35541 16099
rect 34204 16068 35541 16096
rect 34204 16056 34210 16068
rect 35529 16065 35541 16068
rect 35575 16065 35587 16099
rect 35529 16059 35587 16065
rect 39298 16056 39304 16108
rect 39356 16096 39362 16108
rect 40017 16099 40075 16105
rect 40017 16096 40029 16099
rect 39356 16068 40029 16096
rect 39356 16056 39362 16068
rect 40017 16065 40029 16068
rect 40063 16065 40075 16099
rect 40017 16059 40075 16065
rect 35805 16031 35863 16037
rect 35805 16028 35817 16031
rect 34072 16000 35817 16028
rect 33689 15991 33747 15997
rect 35805 15997 35817 16000
rect 35851 16028 35863 16031
rect 39758 16028 39764 16040
rect 35851 16000 36860 16028
rect 39719 16000 39764 16028
rect 35851 15997 35863 16000
rect 35805 15991 35863 15997
rect 33704 15960 33732 15991
rect 31726 15932 33732 15960
rect 26844 15864 27936 15892
rect 26844 15852 26850 15864
rect 30650 15852 30656 15904
rect 30708 15892 30714 15904
rect 30837 15895 30895 15901
rect 30837 15892 30849 15895
rect 30708 15864 30849 15892
rect 30708 15852 30714 15864
rect 30837 15861 30849 15864
rect 30883 15861 30895 15895
rect 33226 15892 33232 15904
rect 33187 15864 33232 15892
rect 30837 15855 30895 15861
rect 33226 15852 33232 15864
rect 33284 15852 33290 15904
rect 34790 15852 34796 15904
rect 34848 15892 34854 15904
rect 34885 15895 34943 15901
rect 34885 15892 34897 15895
rect 34848 15864 34897 15892
rect 34848 15852 34854 15864
rect 34885 15861 34897 15864
rect 34931 15861 34943 15895
rect 34885 15855 34943 15861
rect 35069 15895 35127 15901
rect 35069 15861 35081 15895
rect 35115 15892 35127 15895
rect 35621 15895 35679 15901
rect 35621 15892 35633 15895
rect 35115 15864 35633 15892
rect 35115 15861 35127 15864
rect 35069 15855 35127 15861
rect 35621 15861 35633 15864
rect 35667 15861 35679 15895
rect 35621 15855 35679 15861
rect 35710 15852 35716 15904
rect 35768 15892 35774 15904
rect 36832 15892 36860 16000
rect 39758 15988 39764 16000
rect 39816 15988 39822 16040
rect 41141 15963 41199 15969
rect 41141 15929 41153 15963
rect 41187 15960 41199 15963
rect 41386 15960 41414 16136
rect 41874 16124 41880 16136
rect 41932 16164 41938 16176
rect 42613 16167 42671 16173
rect 42613 16164 42625 16167
rect 41932 16136 42625 16164
rect 41932 16124 41938 16136
rect 42613 16133 42625 16136
rect 42659 16133 42671 16167
rect 42613 16127 42671 16133
rect 41601 16099 41659 16105
rect 41601 16065 41613 16099
rect 41647 16065 41659 16099
rect 41782 16096 41788 16108
rect 41743 16068 41788 16096
rect 41601 16059 41659 16065
rect 41187 15932 41414 15960
rect 41616 15960 41644 16059
rect 41782 16056 41788 16068
rect 41840 16056 41846 16108
rect 46934 16056 46940 16108
rect 46992 16096 46998 16108
rect 47029 16099 47087 16105
rect 47029 16096 47041 16099
rect 46992 16068 47041 16096
rect 46992 16056 46998 16068
rect 47029 16065 47041 16068
rect 47075 16065 47087 16099
rect 47029 16059 47087 16065
rect 46382 15988 46388 16040
rect 46440 16028 46446 16040
rect 47949 16031 48007 16037
rect 47949 16028 47961 16031
rect 46440 16000 47961 16028
rect 46440 15988 46446 16000
rect 47949 15997 47961 16000
rect 47995 15997 48007 16031
rect 47949 15991 48007 15997
rect 42058 15960 42064 15972
rect 41616 15932 42064 15960
rect 41187 15929 41199 15932
rect 41141 15923 41199 15929
rect 42058 15920 42064 15932
rect 42116 15960 42122 15972
rect 42981 15963 43039 15969
rect 42981 15960 42993 15963
rect 42116 15932 42993 15960
rect 42116 15920 42122 15932
rect 42981 15929 42993 15932
rect 43027 15929 43039 15963
rect 42981 15923 43039 15929
rect 40126 15892 40132 15904
rect 35768 15864 35813 15892
rect 36832 15864 40132 15892
rect 35768 15852 35774 15864
rect 40126 15852 40132 15864
rect 40184 15852 40190 15904
rect 41690 15892 41696 15904
rect 41651 15864 41696 15892
rect 41690 15852 41696 15864
rect 41748 15852 41754 15904
rect 41966 15852 41972 15904
rect 42024 15892 42030 15904
rect 42797 15895 42855 15901
rect 42797 15892 42809 15895
rect 42024 15864 42809 15892
rect 42024 15852 42030 15864
rect 42797 15861 42809 15864
rect 42843 15861 42855 15895
rect 42797 15855 42855 15861
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 12894 15688 12900 15700
rect 12855 15660 12900 15688
rect 12894 15648 12900 15660
rect 12952 15648 12958 15700
rect 18874 15688 18880 15700
rect 18835 15660 18880 15688
rect 18874 15648 18880 15660
rect 18932 15648 18938 15700
rect 26234 15688 26240 15700
rect 19628 15660 26096 15688
rect 26195 15660 26240 15688
rect 17494 15580 17500 15632
rect 17552 15620 17558 15632
rect 19628 15620 19656 15660
rect 17552 15592 19656 15620
rect 26068 15620 26096 15660
rect 26234 15648 26240 15660
rect 26292 15648 26298 15700
rect 30469 15691 30527 15697
rect 26988 15660 28212 15688
rect 26988 15620 27016 15660
rect 26068 15592 27016 15620
rect 17552 15580 17558 15592
rect 27062 15580 27068 15632
rect 27120 15580 27126 15632
rect 28077 15623 28135 15629
rect 28077 15589 28089 15623
rect 28123 15589 28135 15623
rect 28077 15583 28135 15589
rect 2774 15552 2780 15564
rect 2735 15524 2780 15552
rect 2774 15512 2780 15524
rect 2832 15512 2838 15564
rect 15010 15552 15016 15564
rect 14971 15524 15016 15552
rect 15010 15512 15016 15524
rect 15068 15512 15074 15564
rect 15102 15512 15108 15564
rect 15160 15552 15166 15564
rect 17678 15552 17684 15564
rect 15160 15524 15205 15552
rect 17591 15524 17684 15552
rect 15160 15512 15166 15524
rect 17678 15512 17684 15524
rect 17736 15552 17742 15564
rect 19334 15552 19340 15564
rect 17736 15524 19340 15552
rect 17736 15512 17742 15524
rect 19334 15512 19340 15524
rect 19392 15552 19398 15564
rect 19981 15555 20039 15561
rect 19981 15552 19993 15555
rect 19392 15524 19993 15552
rect 19392 15512 19398 15524
rect 19981 15521 19993 15524
rect 20027 15521 20039 15555
rect 19981 15515 20039 15521
rect 22094 15512 22100 15564
rect 22152 15552 22158 15564
rect 22649 15555 22707 15561
rect 22649 15552 22661 15555
rect 22152 15524 22661 15552
rect 22152 15512 22158 15524
rect 22649 15521 22661 15524
rect 22695 15521 22707 15555
rect 22649 15515 22707 15521
rect 24762 15512 24768 15564
rect 24820 15552 24826 15564
rect 25777 15555 25835 15561
rect 24820 15524 25636 15552
rect 24820 15512 24826 15524
rect 1578 15484 1584 15496
rect 1539 15456 1584 15484
rect 1578 15444 1584 15456
rect 1636 15444 1642 15496
rect 13078 15484 13084 15496
rect 13039 15456 13084 15484
rect 13078 15444 13084 15456
rect 13136 15444 13142 15496
rect 13725 15487 13783 15493
rect 13725 15453 13737 15487
rect 13771 15484 13783 15487
rect 13771 15456 14596 15484
rect 13771 15453 13783 15456
rect 13725 15447 13783 15453
rect 1765 15419 1823 15425
rect 1765 15385 1777 15419
rect 1811 15385 1823 15419
rect 1765 15379 1823 15385
rect 1780 15348 1808 15379
rect 1946 15376 1952 15428
rect 2004 15416 2010 15428
rect 2406 15416 2412 15428
rect 2004 15388 2412 15416
rect 2004 15376 2010 15388
rect 2406 15376 2412 15388
rect 2464 15376 2470 15428
rect 2866 15348 2872 15360
rect 1780 15320 2872 15348
rect 2866 15308 2872 15320
rect 2924 15308 2930 15360
rect 13541 15351 13599 15357
rect 13541 15317 13553 15351
rect 13587 15348 13599 15351
rect 14090 15348 14096 15360
rect 13587 15320 14096 15348
rect 13587 15317 13599 15320
rect 13541 15311 13599 15317
rect 14090 15308 14096 15320
rect 14148 15308 14154 15360
rect 14568 15357 14596 15456
rect 17034 15444 17040 15496
rect 17092 15484 17098 15496
rect 17402 15484 17408 15496
rect 17092 15456 17408 15484
rect 17092 15444 17098 15456
rect 17402 15444 17408 15456
rect 17460 15444 17466 15496
rect 19797 15487 19855 15493
rect 19797 15484 19809 15487
rect 18432 15456 19809 15484
rect 14921 15419 14979 15425
rect 14921 15385 14933 15419
rect 14967 15416 14979 15419
rect 18432 15416 18460 15456
rect 19797 15453 19809 15456
rect 19843 15453 19855 15487
rect 19797 15447 19855 15453
rect 19889 15487 19947 15493
rect 19889 15453 19901 15487
rect 19935 15484 19947 15487
rect 19935 15456 24532 15484
rect 19935 15453 19947 15456
rect 19889 15447 19947 15453
rect 14967 15388 18460 15416
rect 18509 15419 18567 15425
rect 14967 15385 14979 15388
rect 14921 15379 14979 15385
rect 18509 15385 18521 15419
rect 18555 15385 18567 15419
rect 18509 15379 18567 15385
rect 14553 15351 14611 15357
rect 14553 15317 14565 15351
rect 14599 15317 14611 15351
rect 14553 15311 14611 15317
rect 17037 15351 17095 15357
rect 17037 15317 17049 15351
rect 17083 15348 17095 15351
rect 17126 15348 17132 15360
rect 17083 15320 17132 15348
rect 17083 15317 17095 15320
rect 17037 15311 17095 15317
rect 17126 15308 17132 15320
rect 17184 15308 17190 15360
rect 17494 15348 17500 15360
rect 17455 15320 17500 15348
rect 17494 15308 17500 15320
rect 17552 15308 17558 15360
rect 18524 15348 18552 15379
rect 18598 15376 18604 15428
rect 18656 15416 18662 15428
rect 18693 15419 18751 15425
rect 18693 15416 18705 15419
rect 18656 15388 18705 15416
rect 18656 15376 18662 15388
rect 18693 15385 18705 15388
rect 18739 15385 18751 15419
rect 19812 15416 19840 15447
rect 19978 15416 19984 15428
rect 19812 15388 19984 15416
rect 18693 15379 18751 15385
rect 19978 15376 19984 15388
rect 20036 15376 20042 15428
rect 22916 15419 22974 15425
rect 22916 15385 22928 15419
rect 22962 15416 22974 15419
rect 23198 15416 23204 15428
rect 22962 15388 23204 15416
rect 22962 15385 22974 15388
rect 22916 15379 22974 15385
rect 23198 15376 23204 15388
rect 23256 15376 23262 15428
rect 24504 15416 24532 15456
rect 24578 15444 24584 15496
rect 24636 15484 24642 15496
rect 25608 15493 25636 15524
rect 25777 15521 25789 15555
rect 25823 15552 25835 15555
rect 26510 15552 26516 15564
rect 25823 15524 26516 15552
rect 25823 15521 25835 15524
rect 25777 15515 25835 15521
rect 26252 15493 26280 15524
rect 26510 15512 26516 15524
rect 26568 15512 26574 15564
rect 27080 15552 27108 15580
rect 26896 15524 27108 15552
rect 25409 15487 25467 15493
rect 25409 15484 25421 15487
rect 24636 15456 25421 15484
rect 24636 15444 24642 15456
rect 25409 15453 25421 15456
rect 25455 15453 25467 15487
rect 25409 15447 25467 15453
rect 25593 15487 25651 15493
rect 25593 15453 25605 15487
rect 25639 15453 25651 15487
rect 25593 15447 25651 15453
rect 26237 15487 26295 15493
rect 26237 15453 26249 15487
rect 26283 15453 26295 15487
rect 26418 15484 26424 15496
rect 26379 15456 26424 15484
rect 26237 15447 26295 15453
rect 26418 15444 26424 15456
rect 26476 15444 26482 15496
rect 26896 15493 26924 15524
rect 27246 15512 27252 15564
rect 27304 15552 27310 15564
rect 27617 15555 27675 15561
rect 27617 15552 27629 15555
rect 27304 15524 27629 15552
rect 27304 15512 27310 15524
rect 27617 15521 27629 15524
rect 27663 15521 27675 15555
rect 27617 15515 27675 15521
rect 26881 15487 26939 15493
rect 26881 15453 26893 15487
rect 26927 15453 26939 15487
rect 27062 15484 27068 15496
rect 27023 15456 27068 15484
rect 26881 15447 26939 15453
rect 27062 15444 27068 15456
rect 27120 15444 27126 15496
rect 27709 15487 27767 15493
rect 27709 15453 27721 15487
rect 27755 15453 27767 15487
rect 28092 15484 28120 15583
rect 28184 15552 28212 15660
rect 30469 15657 30481 15691
rect 30515 15688 30527 15691
rect 30558 15688 30564 15700
rect 30515 15660 30564 15688
rect 30515 15657 30527 15660
rect 30469 15651 30527 15657
rect 30558 15648 30564 15660
rect 30616 15648 30622 15700
rect 30834 15688 30840 15700
rect 30795 15660 30840 15688
rect 30834 15648 30840 15660
rect 30892 15648 30898 15700
rect 39298 15688 39304 15700
rect 39259 15660 39304 15688
rect 39298 15648 39304 15660
rect 39356 15648 39362 15700
rect 40770 15648 40776 15700
rect 40828 15688 40834 15700
rect 42702 15688 42708 15700
rect 40828 15660 42708 15688
rect 40828 15648 40834 15660
rect 42702 15648 42708 15660
rect 42760 15648 42766 15700
rect 28258 15580 28264 15632
rect 28316 15620 28322 15632
rect 28316 15592 37412 15620
rect 28316 15580 28322 15592
rect 30926 15552 30932 15564
rect 28184 15524 30932 15552
rect 30926 15512 30932 15524
rect 30984 15512 30990 15564
rect 35710 15552 35716 15564
rect 35084 15524 35716 15552
rect 28537 15487 28595 15493
rect 28537 15484 28549 15487
rect 28092 15456 28549 15484
rect 27709 15447 27767 15453
rect 28537 15453 28549 15456
rect 28583 15453 28595 15487
rect 28537 15447 28595 15453
rect 26786 15416 26792 15428
rect 24504 15388 26792 15416
rect 26786 15376 26792 15388
rect 26844 15376 26850 15428
rect 26973 15419 27031 15425
rect 26973 15385 26985 15419
rect 27019 15416 27031 15419
rect 27338 15416 27344 15428
rect 27019 15388 27344 15416
rect 27019 15385 27031 15388
rect 26973 15379 27031 15385
rect 27338 15376 27344 15388
rect 27396 15416 27402 15428
rect 27724 15416 27752 15447
rect 28626 15444 28632 15496
rect 28684 15484 28690 15496
rect 28721 15487 28779 15493
rect 28721 15484 28733 15487
rect 28684 15456 28733 15484
rect 28684 15444 28690 15456
rect 28721 15453 28733 15456
rect 28767 15453 28779 15487
rect 30650 15484 30656 15496
rect 30611 15456 30656 15484
rect 28721 15447 28779 15453
rect 30650 15444 30656 15456
rect 30708 15444 30714 15496
rect 33226 15444 33232 15496
rect 33284 15484 33290 15496
rect 35084 15493 35112 15524
rect 35710 15512 35716 15524
rect 35768 15512 35774 15564
rect 34885 15487 34943 15493
rect 34885 15484 34897 15487
rect 33284 15456 34897 15484
rect 33284 15444 33290 15456
rect 34885 15453 34897 15456
rect 34931 15453 34943 15487
rect 34885 15447 34943 15453
rect 35069 15487 35127 15493
rect 35069 15453 35081 15487
rect 35115 15453 35127 15487
rect 35069 15447 35127 15453
rect 35253 15487 35311 15493
rect 35253 15453 35265 15487
rect 35299 15484 35311 15487
rect 37090 15484 37096 15496
rect 35299 15456 37096 15484
rect 35299 15453 35311 15456
rect 35253 15447 35311 15453
rect 37090 15444 37096 15456
rect 37148 15444 37154 15496
rect 37384 15493 37412 15592
rect 40770 15552 40776 15564
rect 40731 15524 40776 15552
rect 40770 15512 40776 15524
rect 40828 15512 40834 15564
rect 41782 15552 41788 15564
rect 41743 15524 41788 15552
rect 41782 15512 41788 15524
rect 41840 15512 41846 15564
rect 41874 15512 41880 15564
rect 41932 15552 41938 15564
rect 42702 15552 42708 15564
rect 41932 15524 41977 15552
rect 42663 15524 42708 15552
rect 41932 15512 41938 15524
rect 42702 15512 42708 15524
rect 42760 15512 42766 15564
rect 46477 15555 46535 15561
rect 46477 15521 46489 15555
rect 46523 15552 46535 15555
rect 47946 15552 47952 15564
rect 46523 15524 47952 15552
rect 46523 15521 46535 15524
rect 46477 15515 46535 15521
rect 47946 15512 47952 15524
rect 48004 15512 48010 15564
rect 48222 15552 48228 15564
rect 48183 15524 48228 15552
rect 48222 15512 48228 15524
rect 48280 15512 48286 15564
rect 37369 15487 37427 15493
rect 37369 15453 37381 15487
rect 37415 15453 37427 15487
rect 37369 15447 37427 15453
rect 37645 15487 37703 15493
rect 37645 15453 37657 15487
rect 37691 15484 37703 15487
rect 38930 15484 38936 15496
rect 37691 15456 38936 15484
rect 37691 15453 37703 15456
rect 37645 15447 37703 15453
rect 38930 15444 38936 15456
rect 38988 15444 38994 15496
rect 39485 15487 39543 15493
rect 39485 15453 39497 15487
rect 39531 15484 39543 15487
rect 40494 15484 40500 15496
rect 39531 15456 40500 15484
rect 39531 15453 39543 15456
rect 39485 15447 39543 15453
rect 40494 15444 40500 15456
rect 40552 15444 40558 15496
rect 41598 15484 41604 15496
rect 41559 15456 41604 15484
rect 41598 15444 41604 15456
rect 41656 15444 41662 15496
rect 41693 15487 41751 15493
rect 41693 15453 41705 15487
rect 41739 15484 41751 15487
rect 41966 15484 41972 15496
rect 41739 15456 41972 15484
rect 41739 15453 41751 15456
rect 41693 15447 41751 15453
rect 41966 15444 41972 15456
rect 42024 15444 42030 15496
rect 29270 15416 29276 15428
rect 27396 15388 27752 15416
rect 28460 15388 29276 15416
rect 27396 15376 27402 15388
rect 19429 15351 19487 15357
rect 19429 15348 19441 15351
rect 18524 15320 19441 15348
rect 19429 15317 19441 15320
rect 19475 15317 19487 15351
rect 19429 15311 19487 15317
rect 23658 15308 23664 15360
rect 23716 15348 23722 15360
rect 24029 15351 24087 15357
rect 24029 15348 24041 15351
rect 23716 15320 24041 15348
rect 23716 15308 23722 15320
rect 24029 15317 24041 15320
rect 24075 15348 24087 15351
rect 24578 15348 24584 15360
rect 24075 15320 24584 15348
rect 24075 15317 24087 15320
rect 24029 15311 24087 15317
rect 24578 15308 24584 15320
rect 24636 15308 24642 15360
rect 26694 15308 26700 15360
rect 26752 15348 26758 15360
rect 28460 15348 28488 15388
rect 29270 15376 29276 15388
rect 29328 15376 29334 15428
rect 34514 15376 34520 15428
rect 34572 15416 34578 15428
rect 35161 15419 35219 15425
rect 35161 15416 35173 15419
rect 34572 15388 35173 15416
rect 34572 15376 34578 15388
rect 35161 15385 35173 15388
rect 35207 15416 35219 15419
rect 35710 15416 35716 15428
rect 35207 15388 35716 15416
rect 35207 15385 35219 15388
rect 35161 15379 35219 15385
rect 35710 15376 35716 15388
rect 35768 15376 35774 15428
rect 40034 15416 40040 15428
rect 39995 15388 40040 15416
rect 40034 15376 40040 15388
rect 40092 15376 40098 15428
rect 42972 15419 43030 15425
rect 42972 15385 42984 15419
rect 43018 15416 43030 15419
rect 43070 15416 43076 15428
rect 43018 15388 43076 15416
rect 43018 15385 43030 15388
rect 42972 15379 43030 15385
rect 43070 15376 43076 15388
rect 43128 15376 43134 15428
rect 46661 15419 46719 15425
rect 46661 15385 46673 15419
rect 46707 15416 46719 15419
rect 47118 15416 47124 15428
rect 46707 15388 47124 15416
rect 46707 15385 46719 15388
rect 46661 15379 46719 15385
rect 47118 15376 47124 15388
rect 47176 15376 47182 15428
rect 26752 15320 28488 15348
rect 26752 15308 26758 15320
rect 28534 15308 28540 15360
rect 28592 15348 28598 15360
rect 28629 15351 28687 15357
rect 28629 15348 28641 15351
rect 28592 15320 28641 15348
rect 28592 15308 28598 15320
rect 28629 15317 28641 15320
rect 28675 15317 28687 15351
rect 35434 15348 35440 15360
rect 35395 15320 35440 15348
rect 28629 15311 28687 15317
rect 35434 15308 35440 15320
rect 35492 15308 35498 15360
rect 37185 15351 37243 15357
rect 37185 15317 37197 15351
rect 37231 15348 37243 15351
rect 37366 15348 37372 15360
rect 37231 15320 37372 15348
rect 37231 15317 37243 15320
rect 37185 15311 37243 15317
rect 37366 15308 37372 15320
rect 37424 15308 37430 15360
rect 37553 15351 37611 15357
rect 37553 15317 37565 15351
rect 37599 15348 37611 15351
rect 38930 15348 38936 15360
rect 37599 15320 38936 15348
rect 37599 15317 37611 15320
rect 37553 15311 37611 15317
rect 38930 15308 38936 15320
rect 38988 15308 38994 15360
rect 41414 15308 41420 15360
rect 41472 15348 41478 15360
rect 44082 15348 44088 15360
rect 41472 15320 41517 15348
rect 44043 15320 44088 15348
rect 41472 15308 41478 15320
rect 44082 15308 44088 15320
rect 44140 15308 44146 15360
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 2866 15144 2872 15156
rect 2827 15116 2872 15144
rect 2866 15104 2872 15116
rect 2924 15104 2930 15156
rect 15194 15144 15200 15156
rect 15155 15116 15200 15144
rect 15194 15104 15200 15116
rect 15252 15104 15258 15156
rect 17313 15147 17371 15153
rect 17313 15144 17325 15147
rect 16546 15116 17325 15144
rect 4614 15076 4620 15088
rect 3804 15048 4620 15076
rect 1578 14968 1584 15020
rect 1636 15008 1642 15020
rect 2317 15011 2375 15017
rect 2317 15008 2329 15011
rect 1636 14980 2329 15008
rect 1636 14968 1642 14980
rect 2317 14977 2329 14980
rect 2363 14977 2375 15011
rect 2317 14971 2375 14977
rect 2498 14968 2504 15020
rect 2556 15008 2562 15020
rect 2777 15011 2835 15017
rect 2777 15008 2789 15011
rect 2556 14980 2789 15008
rect 2556 14968 2562 14980
rect 2777 14977 2789 14980
rect 2823 15008 2835 15011
rect 3234 15008 3240 15020
rect 2823 14980 3240 15008
rect 2823 14977 2835 14980
rect 2777 14971 2835 14977
rect 3234 14968 3240 14980
rect 3292 14968 3298 15020
rect 3804 15017 3832 15048
rect 4614 15036 4620 15048
rect 4672 15036 4678 15088
rect 14090 15085 14096 15088
rect 14084 15076 14096 15085
rect 14051 15048 14096 15076
rect 14084 15039 14096 15048
rect 14090 15036 14096 15039
rect 14148 15036 14154 15088
rect 3789 15011 3847 15017
rect 3789 14977 3801 15011
rect 3835 14977 3847 15011
rect 3789 14971 3847 14977
rect 13817 15011 13875 15017
rect 13817 14977 13829 15011
rect 13863 15008 13875 15011
rect 13906 15008 13912 15020
rect 13863 14980 13912 15008
rect 13863 14977 13875 14980
rect 13817 14971 13875 14977
rect 13906 14968 13912 14980
rect 13964 14968 13970 15020
rect 16301 15011 16359 15017
rect 16301 14977 16313 15011
rect 16347 15008 16359 15011
rect 16546 15008 16574 15116
rect 17313 15113 17325 15116
rect 17359 15113 17371 15147
rect 17313 15107 17371 15113
rect 19889 15147 19947 15153
rect 19889 15113 19901 15147
rect 19935 15144 19947 15147
rect 19978 15144 19984 15156
rect 19935 15116 19984 15144
rect 19935 15113 19947 15116
rect 19889 15107 19947 15113
rect 19978 15104 19984 15116
rect 20036 15104 20042 15156
rect 27154 15104 27160 15156
rect 27212 15144 27218 15156
rect 27249 15147 27307 15153
rect 27249 15144 27261 15147
rect 27212 15116 27261 15144
rect 27212 15104 27218 15116
rect 27249 15113 27261 15116
rect 27295 15113 27307 15147
rect 35710 15144 35716 15156
rect 35671 15116 35716 15144
rect 27249 15107 27307 15113
rect 35710 15104 35716 15116
rect 35768 15104 35774 15156
rect 40339 15147 40397 15153
rect 40339 15113 40351 15147
rect 40385 15144 40397 15147
rect 41414 15144 41420 15156
rect 40385 15116 41420 15144
rect 40385 15113 40397 15116
rect 40339 15107 40397 15113
rect 41414 15104 41420 15116
rect 41472 15104 41478 15156
rect 43070 15144 43076 15156
rect 43031 15116 43076 15144
rect 43070 15104 43076 15116
rect 43128 15104 43134 15156
rect 47118 15144 47124 15156
rect 43180 15116 43576 15144
rect 47079 15116 47124 15144
rect 16853 15079 16911 15085
rect 16853 15045 16865 15079
rect 16899 15076 16911 15079
rect 18598 15076 18604 15088
rect 16899 15048 18604 15076
rect 16899 15045 16911 15048
rect 16853 15039 16911 15045
rect 18598 15036 18604 15048
rect 18656 15036 18662 15088
rect 18776 15079 18834 15085
rect 18776 15045 18788 15079
rect 18822 15076 18834 15079
rect 19150 15076 19156 15088
rect 18822 15048 19156 15076
rect 18822 15045 18834 15048
rect 18776 15039 18834 15045
rect 19150 15036 19156 15048
rect 19208 15036 19214 15088
rect 29086 15076 29092 15088
rect 28736 15048 29092 15076
rect 16347 14980 16574 15008
rect 16347 14977 16359 14980
rect 16301 14971 16359 14977
rect 16758 14968 16764 15020
rect 16816 15008 16822 15020
rect 18509 15011 18567 15017
rect 18509 15008 18521 15011
rect 16816 14980 18521 15008
rect 16816 14968 16822 14980
rect 18509 14977 18521 14980
rect 18555 14977 18567 15011
rect 18509 14971 18567 14977
rect 23014 14968 23020 15020
rect 23072 15008 23078 15020
rect 23385 15011 23443 15017
rect 23385 15008 23397 15011
rect 23072 14980 23397 15008
rect 23072 14968 23078 14980
rect 23385 14977 23397 14980
rect 23431 14977 23443 15011
rect 23385 14971 23443 14977
rect 23661 15011 23719 15017
rect 23661 14977 23673 15011
rect 23707 14977 23719 15011
rect 23842 15008 23848 15020
rect 23803 14980 23848 15008
rect 23661 14971 23719 14977
rect 3973 14943 4031 14949
rect 3973 14909 3985 14943
rect 4019 14940 4031 14943
rect 4062 14940 4068 14952
rect 4019 14912 4068 14940
rect 4019 14909 4031 14912
rect 3973 14903 4031 14909
rect 4062 14900 4068 14912
rect 4120 14900 4126 14952
rect 5350 14940 5356 14952
rect 5311 14912 5356 14940
rect 5350 14900 5356 14912
rect 5408 14900 5414 14952
rect 23106 14900 23112 14952
rect 23164 14940 23170 14952
rect 23676 14940 23704 14971
rect 23842 14968 23848 14980
rect 23900 14968 23906 15020
rect 27157 15011 27215 15017
rect 27157 14977 27169 15011
rect 27203 14977 27215 15011
rect 27157 14971 27215 14977
rect 23164 14912 23704 14940
rect 23164 14900 23170 14912
rect 26326 14900 26332 14952
rect 26384 14940 26390 14952
rect 27172 14940 27200 14971
rect 27246 14968 27252 15020
rect 27304 15008 27310 15020
rect 28736 15017 28764 15048
rect 29086 15036 29092 15048
rect 29144 15076 29150 15088
rect 30282 15076 30288 15088
rect 29144 15048 30288 15076
rect 29144 15036 29150 15048
rect 30282 15036 30288 15048
rect 30340 15036 30346 15088
rect 30374 15036 30380 15088
rect 30432 15076 30438 15088
rect 34600 15079 34658 15085
rect 30432 15048 32904 15076
rect 30432 15036 30438 15048
rect 28994 15017 29000 15020
rect 27341 15011 27399 15017
rect 27341 15008 27353 15011
rect 27304 14980 27353 15008
rect 27304 14968 27310 14980
rect 27341 14977 27353 14980
rect 27387 14977 27399 15011
rect 27341 14971 27399 14977
rect 28721 15011 28779 15017
rect 28721 14977 28733 15011
rect 28767 14977 28779 15011
rect 28721 14971 28779 14977
rect 28988 14971 29000 15017
rect 29052 15008 29058 15020
rect 32674 15008 32680 15020
rect 29052 14980 29088 15008
rect 32635 14980 32680 15008
rect 28994 14968 29000 14971
rect 29052 14968 29058 14980
rect 32674 14968 32680 14980
rect 32732 14968 32738 15020
rect 32876 15017 32904 15048
rect 34600 15045 34612 15079
rect 34646 15076 34658 15079
rect 35434 15076 35440 15088
rect 34646 15048 35440 15076
rect 34646 15045 34658 15048
rect 34600 15039 34658 15045
rect 35434 15036 35440 15048
rect 35492 15036 35498 15088
rect 37366 15036 37372 15088
rect 37424 15076 37430 15088
rect 37706 15079 37764 15085
rect 37706 15076 37718 15079
rect 37424 15048 37718 15076
rect 37424 15036 37430 15048
rect 37706 15045 37718 15048
rect 37752 15045 37764 15079
rect 37706 15039 37764 15045
rect 40129 15079 40187 15085
rect 40129 15045 40141 15079
rect 40175 15076 40187 15079
rect 40218 15076 40224 15088
rect 40175 15048 40224 15076
rect 40175 15045 40187 15048
rect 40129 15039 40187 15045
rect 40218 15036 40224 15048
rect 40276 15036 40282 15088
rect 42794 15036 42800 15088
rect 42852 15076 42858 15088
rect 43180 15076 43208 15116
rect 42852 15048 43208 15076
rect 43548 15085 43576 15116
rect 47118 15104 47124 15116
rect 47176 15104 47182 15156
rect 43548 15079 43617 15085
rect 43548 15048 43571 15079
rect 42852 15036 42858 15048
rect 43559 15045 43571 15048
rect 43605 15045 43617 15079
rect 43559 15039 43617 15045
rect 32861 15011 32919 15017
rect 32861 14977 32873 15011
rect 32907 14977 32919 15011
rect 37458 15008 37464 15020
rect 37419 14980 37464 15008
rect 32861 14971 32919 14977
rect 37458 14968 37464 14980
rect 37516 14968 37522 15020
rect 43257 15011 43315 15017
rect 43257 14977 43269 15011
rect 43303 14977 43315 15011
rect 43257 14971 43315 14977
rect 43349 15011 43407 15017
rect 43349 14977 43361 15011
rect 43395 14977 43407 15011
rect 43349 14971 43407 14977
rect 26384 14912 28764 14940
rect 26384 14900 26390 14912
rect 17126 14872 17132 14884
rect 17087 14844 17132 14872
rect 17126 14832 17132 14844
rect 17184 14832 17190 14884
rect 28736 14816 28764 14912
rect 32766 14900 32772 14952
rect 32824 14940 32830 14952
rect 32953 14943 33011 14949
rect 32953 14940 32965 14943
rect 32824 14912 32965 14940
rect 32824 14900 32830 14912
rect 32953 14909 32965 14912
rect 32999 14909 33011 14943
rect 32953 14903 33011 14909
rect 34333 14943 34391 14949
rect 34333 14909 34345 14943
rect 34379 14909 34391 14943
rect 34333 14903 34391 14909
rect 30282 14832 30288 14884
rect 30340 14872 30346 14884
rect 33686 14872 33692 14884
rect 30340 14844 33692 14872
rect 30340 14832 30346 14844
rect 33686 14832 33692 14844
rect 33744 14872 33750 14884
rect 34348 14872 34376 14903
rect 41690 14872 41696 14884
rect 33744 14844 34376 14872
rect 40328 14844 41696 14872
rect 33744 14832 33750 14844
rect 16114 14804 16120 14816
rect 16075 14776 16120 14804
rect 16114 14764 16120 14776
rect 16172 14764 16178 14816
rect 23201 14807 23259 14813
rect 23201 14773 23213 14807
rect 23247 14804 23259 14807
rect 23382 14804 23388 14816
rect 23247 14776 23388 14804
rect 23247 14773 23259 14776
rect 23201 14767 23259 14773
rect 23382 14764 23388 14776
rect 23440 14764 23446 14816
rect 28718 14764 28724 14816
rect 28776 14804 28782 14816
rect 30101 14807 30159 14813
rect 30101 14804 30113 14807
rect 28776 14776 30113 14804
rect 28776 14764 28782 14776
rect 30101 14773 30113 14776
rect 30147 14773 30159 14807
rect 30101 14767 30159 14773
rect 32493 14807 32551 14813
rect 32493 14773 32505 14807
rect 32539 14804 32551 14807
rect 32582 14804 32588 14816
rect 32539 14776 32588 14804
rect 32539 14773 32551 14776
rect 32493 14767 32551 14773
rect 32582 14764 32588 14776
rect 32640 14764 32646 14816
rect 38194 14764 38200 14816
rect 38252 14804 38258 14816
rect 40328 14813 40356 14844
rect 41690 14832 41696 14844
rect 41748 14832 41754 14884
rect 43272 14872 43300 14971
rect 43364 14940 43392 14971
rect 43438 14968 43444 15020
rect 43496 15008 43502 15020
rect 43496 14980 43541 15008
rect 43496 14968 43502 14980
rect 43714 14968 43720 15020
rect 43772 15008 43778 15020
rect 44082 15008 44088 15020
rect 43772 14980 44088 15008
rect 43772 14968 43778 14980
rect 44082 14968 44088 14980
rect 44140 14968 44146 15020
rect 44174 14968 44180 15020
rect 44232 15008 44238 15020
rect 47026 15008 47032 15020
rect 44232 14980 44277 15008
rect 46987 14980 47032 15008
rect 44232 14968 44238 14980
rect 47026 14968 47032 14980
rect 47084 14968 47090 15020
rect 47946 15008 47952 15020
rect 47907 14980 47952 15008
rect 47946 14968 47952 14980
rect 48004 14968 48010 15020
rect 44358 14940 44364 14952
rect 43364 14912 44364 14940
rect 44358 14900 44364 14912
rect 44416 14900 44422 14952
rect 44450 14900 44456 14952
rect 44508 14940 44514 14952
rect 44508 14912 44553 14940
rect 44508 14900 44514 14912
rect 43272 14844 44404 14872
rect 38841 14807 38899 14813
rect 38841 14804 38853 14807
rect 38252 14776 38853 14804
rect 38252 14764 38258 14776
rect 38841 14773 38853 14776
rect 38887 14773 38899 14807
rect 38841 14767 38899 14773
rect 40313 14807 40371 14813
rect 40313 14773 40325 14807
rect 40359 14773 40371 14807
rect 40494 14804 40500 14816
rect 40455 14776 40500 14804
rect 40313 14767 40371 14773
rect 40494 14764 40500 14776
rect 40552 14764 40558 14816
rect 44266 14804 44272 14816
rect 44227 14776 44272 14804
rect 44266 14764 44272 14776
rect 44324 14764 44330 14816
rect 44376 14813 44404 14844
rect 44361 14807 44419 14813
rect 44361 14773 44373 14807
rect 44407 14773 44419 14807
rect 44361 14767 44419 14773
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 4062 14600 4068 14612
rect 4023 14572 4068 14600
rect 4062 14560 4068 14572
rect 4120 14560 4126 14612
rect 17402 14600 17408 14612
rect 17363 14572 17408 14600
rect 17402 14560 17408 14572
rect 17460 14560 17466 14612
rect 23198 14600 23204 14612
rect 23159 14572 23204 14600
rect 23198 14560 23204 14572
rect 23256 14560 23262 14612
rect 23569 14603 23627 14609
rect 23569 14569 23581 14603
rect 23615 14600 23627 14603
rect 25038 14600 25044 14612
rect 23615 14572 25044 14600
rect 23615 14569 23627 14572
rect 23569 14563 23627 14569
rect 25038 14560 25044 14572
rect 25096 14560 25102 14612
rect 26697 14603 26755 14609
rect 26697 14569 26709 14603
rect 26743 14600 26755 14603
rect 27062 14600 27068 14612
rect 26743 14572 27068 14600
rect 26743 14569 26755 14572
rect 26697 14563 26755 14569
rect 27062 14560 27068 14572
rect 27120 14560 27126 14612
rect 28994 14560 29000 14612
rect 29052 14600 29058 14612
rect 29181 14603 29239 14609
rect 29181 14600 29193 14603
rect 29052 14572 29193 14600
rect 29052 14560 29058 14572
rect 29181 14569 29193 14572
rect 29227 14569 29239 14603
rect 29181 14563 29239 14569
rect 29270 14560 29276 14612
rect 29328 14600 29334 14612
rect 38930 14600 38936 14612
rect 29328 14572 30512 14600
rect 38891 14572 38936 14600
rect 29328 14560 29334 14572
rect 22554 14492 22560 14544
rect 22612 14532 22618 14544
rect 23014 14532 23020 14544
rect 22612 14504 23020 14532
rect 22612 14492 22618 14504
rect 23014 14492 23020 14504
rect 23072 14532 23078 14544
rect 23072 14504 27568 14532
rect 23072 14492 23078 14504
rect 2774 14464 2780 14476
rect 2735 14436 2780 14464
rect 2774 14424 2780 14436
rect 2832 14424 2838 14476
rect 23658 14464 23664 14476
rect 23619 14436 23664 14464
rect 23658 14424 23664 14436
rect 23716 14424 23722 14476
rect 27540 14473 27568 14504
rect 27798 14492 27804 14544
rect 27856 14532 27862 14544
rect 27856 14504 30052 14532
rect 27856 14492 27862 14504
rect 27525 14467 27583 14473
rect 27525 14433 27537 14467
rect 27571 14464 27583 14467
rect 29822 14464 29828 14476
rect 27571 14436 29828 14464
rect 27571 14433 27583 14436
rect 27525 14427 27583 14433
rect 29822 14424 29828 14436
rect 29880 14424 29886 14476
rect 30024 14464 30052 14504
rect 30098 14492 30104 14544
rect 30156 14532 30162 14544
rect 30374 14532 30380 14544
rect 30156 14504 30380 14532
rect 30156 14492 30162 14504
rect 30374 14492 30380 14504
rect 30432 14492 30438 14544
rect 30484 14464 30512 14572
rect 38930 14560 38936 14572
rect 38988 14560 38994 14612
rect 41141 14603 41199 14609
rect 41141 14569 41153 14603
rect 41187 14600 41199 14603
rect 41966 14600 41972 14612
rect 41187 14572 41972 14600
rect 41187 14569 41199 14572
rect 41141 14563 41199 14569
rect 41966 14560 41972 14572
rect 42024 14560 42030 14612
rect 44266 14600 44272 14612
rect 44227 14572 44272 14600
rect 44266 14560 44272 14572
rect 44324 14560 44330 14612
rect 44358 14560 44364 14612
rect 44416 14600 44422 14612
rect 44637 14603 44695 14609
rect 44637 14600 44649 14603
rect 44416 14572 44649 14600
rect 44416 14560 44422 14572
rect 44637 14569 44649 14572
rect 44683 14569 44695 14603
rect 44637 14563 44695 14569
rect 37918 14532 37924 14544
rect 31864 14504 37924 14532
rect 31864 14464 31892 14504
rect 37918 14492 37924 14504
rect 37976 14492 37982 14544
rect 33686 14464 33692 14476
rect 30024 14436 30144 14464
rect 30484 14436 31892 14464
rect 33647 14436 33692 14464
rect 1578 14396 1584 14408
rect 1539 14368 1584 14396
rect 1578 14356 1584 14368
rect 1636 14356 1642 14408
rect 3786 14356 3792 14408
rect 3844 14396 3850 14408
rect 3973 14399 4031 14405
rect 3973 14396 3985 14399
rect 3844 14368 3985 14396
rect 3844 14356 3850 14368
rect 3973 14365 3985 14368
rect 4019 14365 4031 14399
rect 3973 14359 4031 14365
rect 16025 14399 16083 14405
rect 16025 14365 16037 14399
rect 16071 14396 16083 14399
rect 16758 14396 16764 14408
rect 16071 14368 16764 14396
rect 16071 14365 16083 14368
rect 16025 14359 16083 14365
rect 16758 14356 16764 14368
rect 16816 14356 16822 14408
rect 23382 14396 23388 14408
rect 23343 14368 23388 14396
rect 23382 14356 23388 14368
rect 23440 14356 23446 14408
rect 24854 14396 24860 14408
rect 24815 14368 24860 14396
rect 24854 14356 24860 14368
rect 24912 14356 24918 14408
rect 25133 14399 25191 14405
rect 25133 14365 25145 14399
rect 25179 14396 25191 14399
rect 25682 14396 25688 14408
rect 25179 14368 25688 14396
rect 25179 14365 25191 14368
rect 25133 14359 25191 14365
rect 25682 14356 25688 14368
rect 25740 14396 25746 14408
rect 26513 14399 26571 14405
rect 26513 14396 26525 14399
rect 25740 14368 26525 14396
rect 25740 14356 25746 14368
rect 26513 14365 26525 14368
rect 26559 14396 26571 14399
rect 27246 14396 27252 14408
rect 26559 14368 27252 14396
rect 26559 14365 26571 14368
rect 26513 14359 26571 14365
rect 27246 14356 27252 14368
rect 27304 14356 27310 14408
rect 27341 14399 27399 14405
rect 27341 14365 27353 14399
rect 27387 14365 27399 14399
rect 27341 14359 27399 14365
rect 27617 14399 27675 14405
rect 27617 14365 27629 14399
rect 27663 14396 27675 14399
rect 27706 14396 27712 14408
rect 27663 14368 27712 14396
rect 27663 14365 27675 14368
rect 27617 14359 27675 14365
rect 1762 14328 1768 14340
rect 1723 14300 1768 14328
rect 1762 14288 1768 14300
rect 1820 14288 1826 14340
rect 16114 14288 16120 14340
rect 16172 14328 16178 14340
rect 16270 14331 16328 14337
rect 16270 14328 16282 14331
rect 16172 14300 16282 14328
rect 16172 14288 16178 14300
rect 16270 14297 16282 14300
rect 16316 14297 16328 14331
rect 26326 14328 26332 14340
rect 26287 14300 26332 14328
rect 16270 14291 16328 14297
rect 26326 14288 26332 14300
rect 26384 14288 26390 14340
rect 24578 14220 24584 14272
rect 24636 14260 24642 14272
rect 24673 14263 24731 14269
rect 24673 14260 24685 14263
rect 24636 14232 24685 14260
rect 24636 14220 24642 14232
rect 24673 14229 24685 14232
rect 24719 14229 24731 14263
rect 24673 14223 24731 14229
rect 27157 14263 27215 14269
rect 27157 14229 27169 14263
rect 27203 14260 27215 14263
rect 27246 14260 27252 14272
rect 27203 14232 27252 14260
rect 27203 14229 27215 14232
rect 27157 14223 27215 14229
rect 27246 14220 27252 14232
rect 27304 14220 27310 14272
rect 27356 14260 27384 14359
rect 27706 14356 27712 14368
rect 27764 14356 27770 14408
rect 28534 14396 28540 14408
rect 28495 14368 28540 14396
rect 28534 14356 28540 14368
rect 28592 14356 28598 14408
rect 28718 14405 28724 14408
rect 28685 14399 28724 14405
rect 28685 14365 28697 14399
rect 28685 14359 28724 14365
rect 28718 14356 28724 14359
rect 28776 14356 28782 14408
rect 29043 14399 29101 14405
rect 29043 14365 29055 14399
rect 29089 14396 29101 14399
rect 29270 14396 29276 14408
rect 29089 14368 29276 14396
rect 29089 14365 29101 14368
rect 29043 14359 29101 14365
rect 29270 14356 29276 14368
rect 29328 14356 29334 14408
rect 29917 14399 29975 14405
rect 29917 14365 29929 14399
rect 29963 14365 29975 14399
rect 30116 14396 30144 14436
rect 30173 14399 30231 14405
rect 30173 14396 30185 14399
rect 30116 14368 30185 14396
rect 29917 14359 29975 14365
rect 30173 14365 30185 14368
rect 30219 14365 30231 14399
rect 31478 14396 31484 14408
rect 31439 14368 31484 14396
rect 30173 14359 30231 14365
rect 28813 14331 28871 14337
rect 28813 14297 28825 14331
rect 28859 14297 28871 14331
rect 28813 14291 28871 14297
rect 27614 14260 27620 14272
rect 27356 14232 27620 14260
rect 27614 14220 27620 14232
rect 27672 14220 27678 14272
rect 28828 14260 28856 14291
rect 28902 14288 28908 14340
rect 28960 14328 28966 14340
rect 29822 14328 29828 14340
rect 28960 14300 29005 14328
rect 29656 14300 29828 14328
rect 28960 14288 28966 14300
rect 29656 14260 29684 14300
rect 29822 14288 29828 14300
rect 29880 14288 29886 14340
rect 29932 14328 29960 14359
rect 31478 14356 31484 14368
rect 31536 14356 31542 14408
rect 31570 14356 31576 14408
rect 31628 14396 31634 14408
rect 31864 14405 31892 14436
rect 33686 14424 33692 14436
rect 33744 14424 33750 14476
rect 43533 14467 43591 14473
rect 43533 14433 43545 14467
rect 43579 14464 43591 14467
rect 43714 14464 43720 14476
rect 43579 14436 43720 14464
rect 43579 14433 43591 14436
rect 43533 14427 43591 14433
rect 43714 14424 43720 14436
rect 43772 14424 43778 14476
rect 43809 14467 43867 14473
rect 43809 14433 43821 14467
rect 43855 14433 43867 14467
rect 43809 14427 43867 14433
rect 31757 14399 31815 14405
rect 31757 14396 31769 14399
rect 31628 14368 31769 14396
rect 31628 14356 31634 14368
rect 31757 14365 31769 14368
rect 31803 14365 31815 14399
rect 31757 14359 31815 14365
rect 31849 14399 31907 14405
rect 31849 14365 31861 14399
rect 31895 14365 31907 14399
rect 31849 14359 31907 14365
rect 31938 14356 31944 14408
rect 31996 14396 32002 14408
rect 32490 14396 32496 14408
rect 31996 14368 32496 14396
rect 31996 14356 32002 14368
rect 32490 14356 32496 14368
rect 32548 14396 32554 14408
rect 32953 14399 33011 14405
rect 32953 14396 32965 14399
rect 32548 14368 32965 14396
rect 32548 14356 32554 14368
rect 32953 14365 32965 14368
rect 32999 14365 33011 14399
rect 32953 14359 33011 14365
rect 37921 14399 37979 14405
rect 37921 14365 37933 14399
rect 37967 14396 37979 14399
rect 38194 14396 38200 14408
rect 37967 14368 38200 14396
rect 37967 14365 37979 14368
rect 37921 14359 37979 14365
rect 38194 14356 38200 14368
rect 38252 14356 38258 14408
rect 38289 14399 38347 14405
rect 38289 14365 38301 14399
rect 38335 14396 38347 14399
rect 38746 14396 38752 14408
rect 38335 14368 38752 14396
rect 38335 14365 38347 14368
rect 38289 14359 38347 14365
rect 38746 14356 38752 14368
rect 38804 14356 38810 14408
rect 38930 14356 38936 14408
rect 38988 14396 38994 14408
rect 40957 14399 41015 14405
rect 40957 14396 40969 14399
rect 38988 14368 40969 14396
rect 38988 14356 38994 14368
rect 40957 14365 40969 14368
rect 41003 14396 41015 14399
rect 42886 14396 42892 14408
rect 41003 14368 42892 14396
rect 41003 14365 41015 14368
rect 40957 14359 41015 14365
rect 42886 14356 42892 14368
rect 42944 14396 42950 14408
rect 43441 14399 43499 14405
rect 43441 14396 43453 14399
rect 42944 14368 43453 14396
rect 42944 14356 42950 14368
rect 43441 14365 43453 14368
rect 43487 14365 43499 14399
rect 43824 14396 43852 14427
rect 44174 14424 44180 14476
rect 44232 14464 44238 14476
rect 44361 14467 44419 14473
rect 44361 14464 44373 14467
rect 44232 14436 44373 14464
rect 44232 14424 44238 14436
rect 44361 14433 44373 14436
rect 44407 14433 44419 14467
rect 44361 14427 44419 14433
rect 44266 14396 44272 14408
rect 43824 14368 44272 14396
rect 43441 14359 43499 14365
rect 44266 14356 44272 14368
rect 44324 14396 44330 14408
rect 44450 14396 44456 14408
rect 44324 14368 44456 14396
rect 44324 14356 44330 14368
rect 44450 14356 44456 14368
rect 44508 14356 44514 14408
rect 29932 14300 30144 14328
rect 28828 14232 29684 14260
rect 29733 14263 29791 14269
rect 29733 14229 29745 14263
rect 29779 14260 29791 14263
rect 30006 14260 30012 14272
rect 29779 14232 30012 14260
rect 29779 14229 29791 14232
rect 29733 14223 29791 14229
rect 30006 14220 30012 14232
rect 30064 14220 30070 14272
rect 30116 14260 30144 14300
rect 30282 14288 30288 14340
rect 30340 14328 30346 14340
rect 31665 14331 31723 14337
rect 31665 14328 31677 14331
rect 30340 14300 31677 14328
rect 30340 14288 30346 14300
rect 31665 14297 31677 14300
rect 31711 14328 31723 14331
rect 37182 14328 37188 14340
rect 31711 14300 37188 14328
rect 31711 14297 31723 14300
rect 31665 14291 31723 14297
rect 37182 14288 37188 14300
rect 37240 14288 37246 14340
rect 40770 14328 40776 14340
rect 40731 14300 40776 14328
rect 40770 14288 40776 14300
rect 40828 14288 40834 14340
rect 30374 14260 30380 14272
rect 30116 14232 30380 14260
rect 30374 14220 30380 14232
rect 30432 14220 30438 14272
rect 32030 14260 32036 14272
rect 31991 14232 32036 14260
rect 32030 14220 32036 14232
rect 32088 14220 32094 14272
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 1762 14016 1768 14068
rect 1820 14056 1826 14068
rect 2869 14059 2927 14065
rect 2869 14056 2881 14059
rect 1820 14028 2881 14056
rect 1820 14016 1826 14028
rect 2869 14025 2881 14028
rect 2915 14025 2927 14059
rect 25682 14056 25688 14068
rect 25643 14028 25688 14056
rect 2869 14019 2927 14025
rect 25682 14016 25688 14028
rect 25740 14016 25746 14068
rect 28258 14016 28264 14068
rect 28316 14056 28322 14068
rect 28537 14059 28595 14065
rect 28537 14056 28549 14059
rect 28316 14028 28549 14056
rect 28316 14016 28322 14028
rect 28537 14025 28549 14028
rect 28583 14056 28595 14059
rect 28902 14056 28908 14068
rect 28583 14028 28908 14056
rect 28583 14025 28595 14028
rect 28537 14019 28595 14025
rect 28902 14016 28908 14028
rect 28960 14016 28966 14068
rect 31018 14016 31024 14068
rect 31076 14056 31082 14068
rect 31113 14059 31171 14065
rect 31113 14056 31125 14059
rect 31076 14028 31125 14056
rect 31076 14016 31082 14028
rect 31113 14025 31125 14028
rect 31159 14056 31171 14059
rect 31570 14056 31576 14068
rect 31159 14028 31576 14056
rect 31159 14025 31171 14028
rect 31113 14019 31171 14025
rect 31570 14016 31576 14028
rect 31628 14016 31634 14068
rect 38010 14016 38016 14068
rect 38068 14056 38074 14068
rect 38841 14059 38899 14065
rect 38841 14056 38853 14059
rect 38068 14028 38853 14056
rect 38068 14016 38074 14028
rect 38841 14025 38853 14028
rect 38887 14025 38899 14059
rect 40770 14056 40776 14068
rect 40731 14028 40776 14056
rect 38841 14019 38899 14025
rect 40770 14016 40776 14028
rect 40828 14016 40834 14068
rect 44174 14016 44180 14068
rect 44232 14056 44238 14068
rect 44637 14059 44695 14065
rect 44637 14056 44649 14059
rect 44232 14028 44649 14056
rect 44232 14016 44238 14028
rect 44637 14025 44649 14028
rect 44683 14025 44695 14059
rect 44637 14019 44695 14025
rect 45462 14016 45468 14068
rect 45520 14056 45526 14068
rect 46569 14059 46627 14065
rect 46569 14056 46581 14059
rect 45520 14028 46581 14056
rect 45520 14016 45526 14028
rect 46569 14025 46581 14028
rect 46615 14025 46627 14059
rect 46569 14019 46627 14025
rect 22554 13988 22560 14000
rect 21100 13960 22560 13988
rect 1578 13880 1584 13932
rect 1636 13920 1642 13932
rect 2317 13923 2375 13929
rect 2317 13920 2329 13923
rect 1636 13892 2329 13920
rect 1636 13880 1642 13892
rect 2317 13889 2329 13892
rect 2363 13889 2375 13923
rect 2317 13883 2375 13889
rect 2777 13923 2835 13929
rect 2777 13889 2789 13923
rect 2823 13920 2835 13923
rect 2958 13920 2964 13932
rect 2823 13892 2964 13920
rect 2823 13889 2835 13892
rect 2777 13883 2835 13889
rect 2958 13880 2964 13892
rect 3016 13880 3022 13932
rect 21100 13852 21128 13960
rect 22554 13948 22560 13960
rect 22612 13948 22618 14000
rect 29086 13988 29092 14000
rect 24320 13960 24716 13988
rect 21177 13923 21235 13929
rect 21177 13889 21189 13923
rect 21223 13920 21235 13923
rect 22005 13923 22063 13929
rect 22005 13920 22017 13923
rect 21223 13892 22017 13920
rect 21223 13889 21235 13892
rect 21177 13883 21235 13889
rect 22005 13889 22017 13892
rect 22051 13889 22063 13923
rect 22186 13920 22192 13932
rect 22147 13892 22192 13920
rect 22005 13883 22063 13889
rect 22186 13880 22192 13892
rect 22244 13880 22250 13932
rect 22462 13920 22468 13932
rect 22423 13892 22468 13920
rect 22462 13880 22468 13892
rect 22520 13880 22526 13932
rect 22646 13880 22652 13932
rect 22704 13920 22710 13932
rect 24320 13929 24348 13960
rect 24578 13929 24584 13932
rect 24305 13923 24363 13929
rect 22704 13892 23796 13920
rect 22704 13880 22710 13892
rect 21361 13855 21419 13861
rect 21361 13852 21373 13855
rect 21100 13824 21373 13852
rect 21361 13821 21373 13824
rect 21407 13821 21419 13855
rect 21361 13815 21419 13821
rect 21453 13855 21511 13861
rect 21453 13821 21465 13855
rect 21499 13852 21511 13855
rect 23290 13852 23296 13864
rect 21499 13824 23296 13852
rect 21499 13821 21511 13824
rect 21453 13815 21511 13821
rect 23290 13812 23296 13824
rect 23348 13812 23354 13864
rect 20990 13716 20996 13728
rect 20951 13688 20996 13716
rect 20990 13676 20996 13688
rect 21048 13676 21054 13728
rect 23768 13716 23796 13892
rect 24305 13889 24317 13923
rect 24351 13889 24363 13923
rect 24572 13920 24584 13929
rect 24539 13892 24584 13920
rect 24305 13883 24363 13889
rect 24572 13883 24584 13892
rect 24578 13880 24584 13883
rect 24636 13880 24642 13932
rect 24688 13920 24716 13960
rect 25700 13960 29092 13988
rect 25700 13920 25728 13960
rect 24688 13892 25728 13920
rect 25774 13880 25780 13932
rect 25832 13920 25838 13932
rect 27172 13929 27200 13960
rect 29086 13948 29092 13960
rect 29144 13948 29150 14000
rect 30006 13997 30012 14000
rect 30000 13988 30012 13997
rect 29967 13960 30012 13988
rect 30000 13951 30012 13960
rect 30006 13948 30012 13951
rect 30064 13948 30070 14000
rect 32582 13997 32588 14000
rect 32576 13988 32588 13997
rect 32543 13960 32588 13988
rect 32576 13951 32588 13960
rect 32582 13948 32588 13951
rect 32640 13948 32646 14000
rect 39758 13988 39764 14000
rect 37476 13960 39764 13988
rect 26145 13923 26203 13929
rect 26145 13920 26157 13923
rect 25832 13892 26157 13920
rect 25832 13880 25838 13892
rect 26145 13889 26157 13892
rect 26191 13889 26203 13923
rect 26145 13883 26203 13889
rect 26329 13923 26387 13929
rect 26329 13889 26341 13923
rect 26375 13889 26387 13923
rect 26329 13883 26387 13889
rect 27157 13923 27215 13929
rect 27157 13889 27169 13923
rect 27203 13889 27215 13923
rect 27157 13883 27215 13889
rect 26344 13716 26372 13883
rect 27246 13880 27252 13932
rect 27304 13920 27310 13932
rect 27413 13923 27471 13929
rect 27413 13920 27425 13923
rect 27304 13892 27425 13920
rect 27304 13880 27310 13892
rect 27413 13889 27425 13892
rect 27459 13889 27471 13923
rect 29104 13920 29132 13948
rect 37476 13929 37504 13960
rect 29733 13923 29791 13929
rect 29733 13920 29745 13923
rect 29104 13892 29745 13920
rect 27413 13883 27471 13889
rect 29733 13889 29745 13892
rect 29779 13889 29791 13923
rect 29733 13883 29791 13889
rect 37461 13923 37519 13929
rect 37461 13889 37473 13923
rect 37507 13889 37519 13923
rect 37461 13883 37519 13889
rect 37550 13880 37556 13932
rect 37608 13920 37614 13932
rect 39408 13929 39436 13960
rect 39758 13948 39764 13960
rect 39816 13988 39822 14000
rect 40862 13988 40868 14000
rect 39816 13960 40868 13988
rect 39816 13948 39822 13960
rect 40862 13948 40868 13960
rect 40920 13948 40926 14000
rect 41506 13948 41512 14000
rect 41564 13988 41570 14000
rect 45480 13988 45508 14016
rect 41564 13960 41736 13988
rect 41564 13948 41570 13960
rect 37717 13923 37775 13929
rect 37717 13920 37729 13923
rect 37608 13892 37729 13920
rect 37608 13880 37614 13892
rect 37717 13889 37729 13892
rect 37763 13889 37775 13923
rect 37717 13883 37775 13889
rect 39393 13923 39451 13929
rect 39393 13889 39405 13923
rect 39439 13889 39451 13923
rect 39393 13883 39451 13889
rect 39660 13923 39718 13929
rect 39660 13889 39672 13923
rect 39706 13920 39718 13923
rect 40126 13920 40132 13932
rect 39706 13892 40132 13920
rect 39706 13889 39718 13892
rect 39660 13883 39718 13889
rect 40126 13880 40132 13892
rect 40184 13880 40190 13932
rect 40218 13880 40224 13932
rect 40276 13920 40282 13932
rect 41233 13923 41291 13929
rect 41233 13920 41245 13923
rect 40276 13892 41245 13920
rect 40276 13880 40282 13892
rect 41233 13889 41245 13892
rect 41279 13889 41291 13923
rect 41233 13883 41291 13889
rect 41417 13923 41475 13929
rect 41417 13889 41429 13923
rect 41463 13889 41475 13923
rect 41598 13920 41604 13932
rect 41559 13892 41604 13920
rect 41417 13883 41475 13889
rect 26510 13852 26516 13864
rect 26471 13824 26516 13852
rect 26510 13812 26516 13824
rect 26568 13812 26574 13864
rect 32306 13852 32312 13864
rect 32267 13824 32312 13852
rect 32306 13812 32312 13824
rect 32364 13812 32370 13864
rect 41432 13852 41460 13883
rect 41598 13880 41604 13892
rect 41656 13880 41662 13932
rect 41708 13929 41736 13960
rect 44468 13960 45508 13988
rect 41693 13923 41751 13929
rect 41693 13889 41705 13923
rect 41739 13920 41751 13923
rect 41966 13920 41972 13932
rect 41739 13892 41972 13920
rect 41739 13889 41751 13892
rect 41693 13883 41751 13889
rect 41966 13880 41972 13892
rect 42024 13880 42030 13932
rect 42886 13880 42892 13932
rect 42944 13920 42950 13932
rect 43533 13923 43591 13929
rect 43533 13920 43545 13923
rect 42944 13892 43545 13920
rect 42944 13880 42950 13892
rect 43533 13889 43545 13892
rect 43579 13889 43591 13923
rect 43714 13920 43720 13932
rect 43675 13892 43720 13920
rect 43533 13883 43591 13889
rect 41782 13852 41788 13864
rect 41432 13824 41788 13852
rect 41782 13812 41788 13824
rect 41840 13812 41846 13864
rect 43548 13852 43576 13883
rect 43714 13880 43720 13892
rect 43772 13880 43778 13932
rect 44468 13929 44496 13960
rect 43809 13923 43867 13929
rect 43809 13889 43821 13923
rect 43855 13920 43867 13923
rect 44453 13923 44511 13929
rect 44453 13920 44465 13923
rect 43855 13892 44465 13920
rect 43855 13889 43867 13892
rect 43809 13883 43867 13889
rect 44453 13889 44465 13892
rect 44499 13889 44511 13923
rect 44453 13883 44511 13889
rect 45456 13923 45514 13929
rect 45456 13889 45468 13923
rect 45502 13920 45514 13923
rect 45738 13920 45744 13932
rect 45502 13892 45744 13920
rect 45502 13889 45514 13892
rect 45456 13883 45514 13889
rect 43622 13852 43628 13864
rect 43548 13824 43628 13852
rect 43622 13812 43628 13824
rect 43680 13812 43686 13864
rect 43530 13744 43536 13796
rect 43588 13784 43594 13796
rect 43824 13784 43852 13883
rect 45738 13880 45744 13892
rect 45796 13880 45802 13932
rect 47026 13920 47032 13932
rect 46987 13892 47032 13920
rect 47026 13880 47032 13892
rect 47084 13880 47090 13932
rect 44269 13855 44327 13861
rect 44269 13821 44281 13855
rect 44315 13852 44327 13855
rect 44634 13852 44640 13864
rect 44315 13824 44640 13852
rect 44315 13821 44327 13824
rect 44269 13815 44327 13821
rect 44634 13812 44640 13824
rect 44692 13812 44698 13864
rect 45094 13812 45100 13864
rect 45152 13852 45158 13864
rect 45189 13855 45247 13861
rect 45189 13852 45201 13855
rect 45152 13824 45201 13852
rect 45152 13812 45158 13824
rect 45189 13821 45201 13824
rect 45235 13821 45247 13855
rect 45189 13815 45247 13821
rect 43588 13756 43852 13784
rect 43588 13744 43594 13756
rect 23768 13688 26372 13716
rect 33689 13719 33747 13725
rect 33689 13685 33701 13719
rect 33735 13716 33747 13719
rect 33778 13716 33784 13728
rect 33735 13688 33784 13716
rect 33735 13685 33747 13688
rect 33689 13679 33747 13685
rect 33778 13676 33784 13688
rect 33836 13676 33842 13728
rect 43349 13719 43407 13725
rect 43349 13685 43361 13719
rect 43395 13716 43407 13719
rect 43622 13716 43628 13728
rect 43395 13688 43628 13716
rect 43395 13685 43407 13688
rect 43349 13679 43407 13685
rect 43622 13676 43628 13688
rect 43680 13676 43686 13728
rect 47118 13716 47124 13728
rect 47079 13688 47124 13716
rect 47118 13676 47124 13688
rect 47176 13676 47182 13728
rect 47946 13716 47952 13728
rect 47907 13688 47952 13716
rect 47946 13676 47952 13688
rect 48004 13676 48010 13728
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 21542 13472 21548 13524
rect 21600 13512 21606 13524
rect 22189 13515 22247 13521
rect 21600 13484 22094 13512
rect 21600 13472 21606 13484
rect 22066 13376 22094 13484
rect 22189 13481 22201 13515
rect 22235 13512 22247 13515
rect 22646 13512 22652 13524
rect 22235 13484 22652 13512
rect 22235 13481 22247 13484
rect 22189 13475 22247 13481
rect 22646 13472 22652 13484
rect 22704 13472 22710 13524
rect 23014 13512 23020 13524
rect 22975 13484 23020 13512
rect 23014 13472 23020 13484
rect 23072 13472 23078 13524
rect 24765 13515 24823 13521
rect 24765 13481 24777 13515
rect 24811 13512 24823 13515
rect 24854 13512 24860 13524
rect 24811 13484 24860 13512
rect 24811 13481 24823 13484
rect 24765 13475 24823 13481
rect 24854 13472 24860 13484
rect 24912 13472 24918 13524
rect 27614 13512 27620 13524
rect 27575 13484 27620 13512
rect 27614 13472 27620 13484
rect 27672 13472 27678 13524
rect 30374 13512 30380 13524
rect 30335 13484 30380 13512
rect 30374 13472 30380 13484
rect 30432 13472 30438 13524
rect 32217 13515 32275 13521
rect 32217 13481 32229 13515
rect 32263 13512 32275 13515
rect 32674 13512 32680 13524
rect 32263 13484 32680 13512
rect 32263 13481 32275 13484
rect 32217 13475 32275 13481
rect 32674 13472 32680 13484
rect 32732 13472 32738 13524
rect 33594 13472 33600 13524
rect 33652 13512 33658 13524
rect 33689 13515 33747 13521
rect 33689 13512 33701 13515
rect 33652 13484 33701 13512
rect 33652 13472 33658 13484
rect 33689 13481 33701 13484
rect 33735 13481 33747 13515
rect 37550 13512 37556 13524
rect 37511 13484 37556 13512
rect 33689 13475 33747 13481
rect 37550 13472 37556 13484
rect 37608 13472 37614 13524
rect 40402 13472 40408 13524
rect 40460 13512 40466 13524
rect 43346 13512 43352 13524
rect 40460 13484 43352 13512
rect 40460 13472 40466 13484
rect 43346 13472 43352 13484
rect 43404 13472 43410 13524
rect 45738 13512 45744 13524
rect 45699 13484 45744 13512
rect 45738 13472 45744 13484
rect 45796 13472 45802 13524
rect 22462 13404 22468 13456
rect 22520 13444 22526 13456
rect 43364 13444 43392 13472
rect 44910 13444 44916 13456
rect 22520 13416 28120 13444
rect 22520 13404 22526 13416
rect 23109 13379 23167 13385
rect 23109 13376 23121 13379
rect 22066 13348 23121 13376
rect 23109 13345 23121 13348
rect 23155 13345 23167 13379
rect 23109 13339 23167 13345
rect 20809 13311 20867 13317
rect 20809 13277 20821 13311
rect 20855 13277 20867 13311
rect 20809 13271 20867 13277
rect 21076 13311 21134 13317
rect 21076 13277 21088 13311
rect 21122 13277 21134 13311
rect 22830 13308 22836 13320
rect 22791 13280 22836 13308
rect 21076 13271 21134 13277
rect 20714 13132 20720 13184
rect 20772 13172 20778 13184
rect 20824 13172 20852 13271
rect 20990 13200 20996 13252
rect 21048 13240 21054 13252
rect 21100 13240 21128 13271
rect 22830 13268 22836 13280
rect 22888 13268 22894 13320
rect 22922 13268 22928 13320
rect 22980 13308 22986 13320
rect 23124 13308 23152 13339
rect 23198 13336 23204 13388
rect 23256 13376 23262 13388
rect 28092 13376 28120 13416
rect 41386 13416 43300 13444
rect 43364 13416 44916 13444
rect 23256 13348 27844 13376
rect 23256 13336 23262 13348
rect 24946 13308 24952 13320
rect 22980 13280 23152 13308
rect 24907 13280 24952 13308
rect 22980 13268 22986 13280
rect 24946 13268 24952 13280
rect 25004 13268 25010 13320
rect 25225 13311 25283 13317
rect 25225 13277 25237 13311
rect 25271 13277 25283 13311
rect 25406 13308 25412 13320
rect 25367 13280 25412 13308
rect 25225 13271 25283 13277
rect 21048 13212 21128 13240
rect 21048 13200 21054 13212
rect 24854 13200 24860 13252
rect 24912 13240 24918 13252
rect 25240 13240 25268 13271
rect 25406 13268 25412 13280
rect 25464 13308 25470 13320
rect 27706 13308 27712 13320
rect 25464 13280 27712 13308
rect 25464 13268 25470 13280
rect 27706 13268 27712 13280
rect 27764 13268 27770 13320
rect 27816 13317 27844 13348
rect 28092 13348 28488 13376
rect 28092 13317 28120 13348
rect 27801 13311 27859 13317
rect 27801 13277 27813 13311
rect 27847 13277 27859 13311
rect 27801 13271 27859 13277
rect 28077 13311 28135 13317
rect 28077 13277 28089 13311
rect 28123 13277 28135 13311
rect 28258 13308 28264 13320
rect 28219 13280 28264 13308
rect 28077 13271 28135 13277
rect 28258 13268 28264 13280
rect 28316 13268 28322 13320
rect 24912 13212 25268 13240
rect 27724 13240 27752 13268
rect 28350 13240 28356 13252
rect 27724 13212 28356 13240
rect 24912 13200 24918 13212
rect 28350 13200 28356 13212
rect 28408 13200 28414 13252
rect 28460 13240 28488 13348
rect 30760 13348 31754 13376
rect 30760 13320 30788 13348
rect 30561 13311 30619 13317
rect 30561 13277 30573 13311
rect 30607 13308 30619 13311
rect 30742 13308 30748 13320
rect 30607 13280 30748 13308
rect 30607 13277 30619 13280
rect 30561 13271 30619 13277
rect 30742 13268 30748 13280
rect 30800 13268 30806 13320
rect 30837 13311 30895 13317
rect 30837 13277 30849 13311
rect 30883 13277 30895 13311
rect 31018 13308 31024 13320
rect 30979 13280 31024 13308
rect 30837 13271 30895 13277
rect 30852 13240 30880 13271
rect 31018 13268 31024 13280
rect 31076 13268 31082 13320
rect 31726 13308 31754 13348
rect 32490 13336 32496 13388
rect 32548 13376 32554 13388
rect 40034 13376 40040 13388
rect 32548 13348 40040 13376
rect 32548 13336 32554 13348
rect 40034 13336 40040 13348
rect 40092 13376 40098 13388
rect 40862 13376 40868 13388
rect 40092 13348 40172 13376
rect 40823 13348 40868 13376
rect 40092 13336 40098 13348
rect 32401 13311 32459 13317
rect 32401 13308 32413 13311
rect 31726 13280 32413 13308
rect 32401 13277 32413 13280
rect 32447 13277 32459 13311
rect 32401 13271 32459 13277
rect 32677 13311 32735 13317
rect 32677 13277 32689 13311
rect 32723 13277 32735 13311
rect 32677 13271 32735 13277
rect 32861 13311 32919 13317
rect 32861 13277 32873 13311
rect 32907 13277 32919 13311
rect 32861 13271 32919 13277
rect 31110 13240 31116 13252
rect 28460 13212 31116 13240
rect 31110 13200 31116 13212
rect 31168 13240 31174 13252
rect 32692 13240 32720 13271
rect 31168 13212 32720 13240
rect 32876 13240 32904 13271
rect 33410 13268 33416 13320
rect 33468 13308 33474 13320
rect 33505 13311 33563 13317
rect 33505 13308 33517 13311
rect 33468 13280 33517 13308
rect 33468 13268 33474 13280
rect 33505 13277 33517 13280
rect 33551 13277 33563 13311
rect 33505 13271 33563 13277
rect 33778 13268 33784 13320
rect 33836 13308 33842 13320
rect 33836 13280 33881 13308
rect 33836 13268 33842 13280
rect 36814 13268 36820 13320
rect 36872 13308 36878 13320
rect 37001 13311 37059 13317
rect 37001 13308 37013 13311
rect 36872 13280 37013 13308
rect 36872 13268 36878 13280
rect 37001 13277 37013 13280
rect 37047 13277 37059 13311
rect 37001 13271 37059 13277
rect 37090 13268 37096 13320
rect 37148 13308 37154 13320
rect 37369 13311 37427 13317
rect 37369 13308 37381 13311
rect 37148 13280 37381 13308
rect 37148 13268 37154 13280
rect 37369 13277 37381 13280
rect 37415 13277 37427 13311
rect 38010 13308 38016 13320
rect 37971 13280 38016 13308
rect 37369 13271 37427 13277
rect 38010 13268 38016 13280
rect 38068 13268 38074 13320
rect 38194 13308 38200 13320
rect 38155 13280 38200 13308
rect 38194 13268 38200 13280
rect 38252 13268 38258 13320
rect 40144 13317 40172 13348
rect 40862 13336 40868 13348
rect 40920 13376 40926 13388
rect 41386 13376 41414 13416
rect 40920 13348 41414 13376
rect 43272 13376 43300 13416
rect 44910 13404 44916 13416
rect 44968 13444 44974 13456
rect 47946 13444 47952 13456
rect 44968 13416 45232 13444
rect 44968 13404 44974 13416
rect 45094 13376 45100 13388
rect 43272 13348 45100 13376
rect 40920 13336 40926 13348
rect 45094 13336 45100 13348
rect 45152 13336 45158 13388
rect 40129 13311 40187 13317
rect 40129 13277 40141 13311
rect 40175 13277 40187 13311
rect 41506 13308 41512 13320
rect 41467 13280 41512 13308
rect 40129 13271 40187 13277
rect 41506 13268 41512 13280
rect 41564 13268 41570 13320
rect 41598 13268 41604 13320
rect 41656 13308 41662 13320
rect 41693 13311 41751 13317
rect 41693 13308 41705 13311
rect 41656 13280 41705 13308
rect 41656 13268 41662 13280
rect 41693 13277 41705 13280
rect 41739 13277 41751 13311
rect 41693 13271 41751 13277
rect 33796 13240 33824 13268
rect 32876 13212 33824 13240
rect 31168 13200 31174 13212
rect 36722 13200 36728 13252
rect 36780 13240 36786 13252
rect 37185 13243 37243 13249
rect 37185 13240 37197 13243
rect 36780 13212 37197 13240
rect 36780 13200 36786 13212
rect 37185 13209 37197 13212
rect 37231 13209 37243 13243
rect 37185 13203 37243 13209
rect 37274 13200 37280 13252
rect 37332 13240 37338 13252
rect 38028 13240 38056 13268
rect 37332 13212 38056 13240
rect 41708 13240 41736 13271
rect 41782 13268 41788 13320
rect 41840 13308 41846 13320
rect 42242 13308 42248 13320
rect 41840 13280 41885 13308
rect 42203 13280 42248 13308
rect 41840 13268 41846 13280
rect 42242 13268 42248 13280
rect 42300 13268 42306 13320
rect 42429 13311 42487 13317
rect 42429 13277 42441 13311
rect 42475 13308 42487 13311
rect 42886 13308 42892 13320
rect 42475 13280 42892 13308
rect 42475 13277 42487 13280
rect 42429 13271 42487 13277
rect 42886 13268 42892 13280
rect 42944 13268 42950 13320
rect 43530 13308 43536 13320
rect 43491 13280 43536 13308
rect 43530 13268 43536 13280
rect 43588 13268 43594 13320
rect 43714 13308 43720 13320
rect 43675 13280 43720 13308
rect 43714 13268 43720 13280
rect 43772 13268 43778 13320
rect 44174 13308 44180 13320
rect 44135 13280 44180 13308
rect 44174 13268 44180 13280
rect 44232 13268 44238 13320
rect 45204 13317 45232 13416
rect 46492 13416 47952 13444
rect 46492 13385 46520 13416
rect 47946 13404 47952 13416
rect 48004 13404 48010 13456
rect 46477 13379 46535 13385
rect 46477 13345 46489 13379
rect 46523 13345 46535 13379
rect 46477 13339 46535 13345
rect 46661 13379 46719 13385
rect 46661 13345 46673 13379
rect 46707 13376 46719 13379
rect 47118 13376 47124 13388
rect 46707 13348 47124 13376
rect 46707 13345 46719 13348
rect 46661 13339 46719 13345
rect 47118 13336 47124 13348
rect 47176 13336 47182 13388
rect 48222 13376 48228 13388
rect 48183 13348 48228 13376
rect 48222 13336 48228 13348
rect 48280 13336 48286 13388
rect 44361 13311 44419 13317
rect 44361 13277 44373 13311
rect 44407 13277 44419 13311
rect 44361 13271 44419 13277
rect 45189 13311 45247 13317
rect 45189 13277 45201 13311
rect 45235 13277 45247 13311
rect 45462 13308 45468 13320
rect 45423 13280 45468 13308
rect 45189 13271 45247 13277
rect 42337 13243 42395 13249
rect 42337 13240 42349 13243
rect 41708 13212 42349 13240
rect 37332 13200 37338 13212
rect 42337 13209 42349 13212
rect 42383 13209 42395 13243
rect 42337 13203 42395 13209
rect 43625 13243 43683 13249
rect 43625 13209 43637 13243
rect 43671 13240 43683 13243
rect 44376 13240 44404 13271
rect 45462 13268 45468 13280
rect 45520 13268 45526 13320
rect 45554 13268 45560 13320
rect 45612 13308 45618 13320
rect 45612 13280 45657 13308
rect 45612 13268 45618 13280
rect 43671 13212 44404 13240
rect 43671 13209 43683 13212
rect 43625 13203 43683 13209
rect 45002 13200 45008 13252
rect 45060 13240 45066 13252
rect 45373 13243 45431 13249
rect 45373 13240 45385 13243
rect 45060 13212 45385 13240
rect 45060 13200 45066 13212
rect 45373 13209 45385 13212
rect 45419 13209 45431 13243
rect 45373 13203 45431 13209
rect 22094 13172 22100 13184
rect 20772 13144 22100 13172
rect 20772 13132 20778 13144
rect 22094 13132 22100 13144
rect 22152 13132 22158 13184
rect 22646 13172 22652 13184
rect 22607 13144 22652 13172
rect 22646 13132 22652 13144
rect 22704 13132 22710 13184
rect 33321 13175 33379 13181
rect 33321 13141 33333 13175
rect 33367 13172 33379 13175
rect 33778 13172 33784 13184
rect 33367 13144 33784 13172
rect 33367 13141 33379 13144
rect 33321 13135 33379 13141
rect 33778 13132 33784 13144
rect 33836 13132 33842 13184
rect 37458 13132 37464 13184
rect 37516 13172 37522 13184
rect 38381 13175 38439 13181
rect 38381 13172 38393 13175
rect 37516 13144 38393 13172
rect 37516 13132 37522 13144
rect 38381 13141 38393 13144
rect 38427 13141 38439 13175
rect 38381 13135 38439 13141
rect 40310 13132 40316 13184
rect 40368 13172 40374 13184
rect 41601 13175 41659 13181
rect 41601 13172 41613 13175
rect 40368 13144 41613 13172
rect 40368 13132 40374 13144
rect 41601 13141 41613 13144
rect 41647 13141 41659 13175
rect 41601 13135 41659 13141
rect 43162 13132 43168 13184
rect 43220 13172 43226 13184
rect 43714 13172 43720 13184
rect 43220 13144 43720 13172
rect 43220 13132 43226 13144
rect 43714 13132 43720 13144
rect 43772 13172 43778 13184
rect 44269 13175 44327 13181
rect 44269 13172 44281 13175
rect 43772 13144 44281 13172
rect 43772 13132 43778 13144
rect 44269 13141 44281 13144
rect 44315 13141 44327 13175
rect 44269 13135 44327 13141
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 22005 12971 22063 12977
rect 22005 12937 22017 12971
rect 22051 12968 22063 12971
rect 22830 12968 22836 12980
rect 22051 12940 22836 12968
rect 22051 12937 22063 12940
rect 22005 12931 22063 12937
rect 22830 12928 22836 12940
rect 22888 12928 22894 12980
rect 40037 12971 40095 12977
rect 40037 12937 40049 12971
rect 40083 12968 40095 12971
rect 40126 12968 40132 12980
rect 40083 12940 40132 12968
rect 40083 12937 40095 12940
rect 40037 12931 40095 12937
rect 40126 12928 40132 12940
rect 40184 12928 40190 12980
rect 40770 12928 40776 12980
rect 40828 12968 40834 12980
rect 40828 12940 41649 12968
rect 40828 12928 40834 12940
rect 23198 12900 23204 12912
rect 22296 12872 23204 12900
rect 22186 12832 22192 12844
rect 22099 12804 22192 12832
rect 22186 12792 22192 12804
rect 22244 12832 22250 12844
rect 22296 12832 22324 12872
rect 23198 12860 23204 12872
rect 23256 12860 23262 12912
rect 32306 12860 32312 12912
rect 32364 12900 32370 12912
rect 33042 12900 33048 12912
rect 32364 12872 33048 12900
rect 32364 12860 32370 12872
rect 33042 12860 33048 12872
rect 33100 12900 33106 12912
rect 33229 12903 33287 12909
rect 33229 12900 33241 12903
rect 33100 12872 33241 12900
rect 33100 12860 33106 12872
rect 33229 12869 33241 12872
rect 33275 12900 33287 12903
rect 40310 12900 40316 12912
rect 33275 12872 33916 12900
rect 40271 12872 40316 12900
rect 33275 12869 33287 12872
rect 33229 12863 33287 12869
rect 22462 12832 22468 12844
rect 22244 12804 22324 12832
rect 22423 12804 22468 12832
rect 22244 12792 22250 12804
rect 22462 12792 22468 12804
rect 22520 12792 22526 12844
rect 22649 12835 22707 12841
rect 22649 12801 22661 12835
rect 22695 12832 22707 12835
rect 22738 12832 22744 12844
rect 22695 12804 22744 12832
rect 22695 12801 22707 12804
rect 22649 12795 22707 12801
rect 22738 12792 22744 12804
rect 22796 12792 22802 12844
rect 32490 12832 32496 12844
rect 32451 12804 32496 12832
rect 32490 12792 32496 12804
rect 32548 12792 32554 12844
rect 33888 12841 33916 12872
rect 40310 12860 40316 12872
rect 40368 12860 40374 12912
rect 41621 12900 41649 12940
rect 41690 12928 41696 12980
rect 41748 12968 41754 12980
rect 41785 12971 41843 12977
rect 41785 12968 41797 12971
rect 41748 12940 41797 12968
rect 41748 12928 41754 12940
rect 41785 12937 41797 12940
rect 41831 12937 41843 12971
rect 41785 12931 41843 12937
rect 42889 12971 42947 12977
rect 42889 12937 42901 12971
rect 42935 12937 42947 12971
rect 45002 12968 45008 12980
rect 44963 12940 45008 12968
rect 42889 12931 42947 12937
rect 42242 12900 42248 12912
rect 41621 12872 42248 12900
rect 34146 12841 34152 12844
rect 33873 12835 33931 12841
rect 33873 12801 33885 12835
rect 33919 12801 33931 12835
rect 33873 12795 33931 12801
rect 34140 12795 34152 12841
rect 34204 12832 34210 12844
rect 36354 12832 36360 12844
rect 34204 12804 34240 12832
rect 36315 12804 36360 12832
rect 34146 12792 34152 12795
rect 34204 12792 34210 12804
rect 36354 12792 36360 12804
rect 36412 12792 36418 12844
rect 37458 12832 37464 12844
rect 37419 12804 37464 12832
rect 37458 12792 37464 12804
rect 37516 12792 37522 12844
rect 37642 12832 37648 12844
rect 37603 12804 37648 12832
rect 37642 12792 37648 12804
rect 37700 12792 37706 12844
rect 40218 12832 40224 12844
rect 40179 12804 40224 12832
rect 40218 12792 40224 12804
rect 40276 12792 40282 12844
rect 40402 12832 40408 12844
rect 40363 12804 40408 12832
rect 40402 12792 40408 12804
rect 40460 12792 40466 12844
rect 40543 12835 40601 12841
rect 40543 12801 40555 12835
rect 40589 12832 40601 12835
rect 41138 12832 41144 12844
rect 40589 12804 41000 12832
rect 41099 12804 41144 12832
rect 40589 12801 40601 12804
rect 40543 12795 40601 12801
rect 36446 12764 36452 12776
rect 36359 12736 36452 12764
rect 36446 12724 36452 12736
rect 36504 12764 36510 12776
rect 36722 12764 36728 12776
rect 36504 12736 36584 12764
rect 36683 12736 36728 12764
rect 36504 12724 36510 12736
rect 36556 12696 36584 12736
rect 36722 12724 36728 12736
rect 36780 12724 36786 12776
rect 40681 12767 40739 12773
rect 40681 12733 40693 12767
rect 40727 12764 40739 12767
rect 40770 12764 40776 12776
rect 40727 12736 40776 12764
rect 40727 12733 40739 12736
rect 40681 12727 40739 12733
rect 40770 12724 40776 12736
rect 40828 12724 40834 12776
rect 37553 12699 37611 12705
rect 37553 12696 37565 12699
rect 36556 12668 37565 12696
rect 37553 12665 37565 12668
rect 37599 12665 37611 12699
rect 37553 12659 37611 12665
rect 34514 12588 34520 12640
rect 34572 12628 34578 12640
rect 35253 12631 35311 12637
rect 35253 12628 35265 12631
rect 34572 12600 35265 12628
rect 34572 12588 34578 12600
rect 35253 12597 35265 12600
rect 35299 12597 35311 12631
rect 35253 12591 35311 12597
rect 36814 12588 36820 12640
rect 36872 12628 36878 12640
rect 40402 12628 40408 12640
rect 36872 12600 40408 12628
rect 36872 12588 36878 12600
rect 40402 12588 40408 12600
rect 40460 12588 40466 12640
rect 40972 12628 41000 12804
rect 41138 12792 41144 12804
rect 41196 12792 41202 12844
rect 41230 12792 41236 12844
rect 41288 12832 41294 12844
rect 41621 12841 41649 12872
rect 42242 12860 42248 12872
rect 42300 12860 42306 12912
rect 42904 12900 42932 12931
rect 45002 12928 45008 12940
rect 45060 12928 45066 12980
rect 42904 12872 44956 12900
rect 41417 12835 41475 12841
rect 41288 12804 41333 12832
rect 41288 12792 41294 12804
rect 41417 12801 41429 12835
rect 41463 12801 41475 12835
rect 41417 12795 41475 12801
rect 41509 12835 41567 12841
rect 41509 12801 41521 12835
rect 41555 12801 41567 12835
rect 41509 12795 41567 12801
rect 41606 12835 41664 12841
rect 41606 12801 41618 12835
rect 41652 12801 41664 12835
rect 42886 12832 42892 12844
rect 42847 12804 42892 12832
rect 41606 12795 41664 12801
rect 41322 12656 41328 12708
rect 41380 12696 41386 12708
rect 41432 12696 41460 12795
rect 41524 12764 41552 12795
rect 42886 12792 42892 12804
rect 42944 12792 42950 12844
rect 42978 12792 42984 12844
rect 43036 12792 43042 12844
rect 43162 12832 43168 12844
rect 43123 12804 43168 12832
rect 43162 12792 43168 12804
rect 43220 12792 43226 12844
rect 44174 12792 44180 12844
rect 44232 12832 44238 12844
rect 44928 12841 44956 12872
rect 44269 12835 44327 12841
rect 44269 12832 44281 12835
rect 44232 12804 44281 12832
rect 44232 12792 44238 12804
rect 44269 12801 44281 12804
rect 44315 12801 44327 12835
rect 44269 12795 44327 12801
rect 44913 12835 44971 12841
rect 44913 12801 44925 12835
rect 44959 12801 44971 12835
rect 44913 12795 44971 12801
rect 45097 12835 45155 12841
rect 45097 12801 45109 12835
rect 45143 12801 45155 12835
rect 45097 12795 45155 12801
rect 47029 12835 47087 12841
rect 47029 12801 47041 12835
rect 47075 12832 47087 12835
rect 47302 12832 47308 12844
rect 47075 12804 47308 12832
rect 47075 12801 47087 12804
rect 47029 12795 47087 12801
rect 42996 12764 43024 12792
rect 44085 12767 44143 12773
rect 44085 12764 44097 12767
rect 41524 12736 43024 12764
rect 44008 12736 44097 12764
rect 41380 12668 41460 12696
rect 42981 12699 43039 12705
rect 41380 12656 41386 12668
rect 42981 12665 42993 12699
rect 43027 12696 43039 12699
rect 43254 12696 43260 12708
rect 43027 12668 43260 12696
rect 43027 12665 43039 12668
rect 42981 12659 43039 12665
rect 43254 12656 43260 12668
rect 43312 12656 43318 12708
rect 42702 12628 42708 12640
rect 40972 12600 42708 12628
rect 42702 12588 42708 12600
rect 42760 12588 42766 12640
rect 42794 12588 42800 12640
rect 42852 12628 42858 12640
rect 44008 12628 44036 12736
rect 44085 12733 44097 12736
rect 44131 12764 44143 12767
rect 44358 12764 44364 12776
rect 44131 12736 44364 12764
rect 44131 12733 44143 12736
rect 44085 12727 44143 12733
rect 44358 12724 44364 12736
rect 44416 12764 44422 12776
rect 45112 12764 45140 12795
rect 47302 12792 47308 12804
rect 47360 12832 47366 12844
rect 47486 12832 47492 12844
rect 47360 12804 47492 12832
rect 47360 12792 47366 12804
rect 47486 12792 47492 12804
rect 47544 12792 47550 12844
rect 44416 12736 45140 12764
rect 44416 12724 44422 12736
rect 42852 12600 44036 12628
rect 44453 12631 44511 12637
rect 42852 12588 42858 12600
rect 44453 12597 44465 12631
rect 44499 12628 44511 12631
rect 44726 12628 44732 12640
rect 44499 12600 44732 12628
rect 44499 12597 44511 12600
rect 44453 12591 44511 12597
rect 44726 12588 44732 12600
rect 44784 12588 44790 12640
rect 47118 12628 47124 12640
rect 47079 12600 47124 12628
rect 47118 12588 47124 12600
rect 47176 12588 47182 12640
rect 47946 12628 47952 12640
rect 47907 12600 47952 12628
rect 47946 12588 47952 12600
rect 48004 12588 48010 12640
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 26068 12396 31754 12424
rect 23014 12356 23020 12368
rect 22756 12328 23020 12356
rect 20714 12288 20720 12300
rect 20675 12260 20720 12288
rect 20714 12248 20720 12260
rect 20772 12248 20778 12300
rect 2038 12180 2044 12232
rect 2096 12220 2102 12232
rect 2225 12223 2283 12229
rect 2225 12220 2237 12223
rect 2096 12192 2237 12220
rect 2096 12180 2102 12192
rect 2225 12189 2237 12192
rect 2271 12189 2283 12223
rect 2225 12183 2283 12189
rect 20984 12223 21042 12229
rect 20984 12189 20996 12223
rect 21030 12220 21042 12223
rect 22646 12220 22652 12232
rect 21030 12192 22652 12220
rect 21030 12189 21042 12192
rect 20984 12183 21042 12189
rect 22646 12180 22652 12192
rect 22704 12180 22710 12232
rect 22756 12229 22784 12328
rect 23014 12316 23020 12328
rect 23072 12316 23078 12368
rect 24302 12248 24308 12300
rect 24360 12288 24366 12300
rect 24360 12260 25728 12288
rect 24360 12248 24366 12260
rect 22741 12223 22799 12229
rect 22741 12189 22753 12223
rect 22787 12189 22799 12223
rect 23014 12220 23020 12232
rect 22975 12192 23020 12220
rect 22741 12183 22799 12189
rect 22462 12112 22468 12164
rect 22520 12152 22526 12164
rect 22756 12152 22784 12183
rect 23014 12180 23020 12192
rect 23072 12180 23078 12232
rect 23201 12223 23259 12229
rect 23201 12189 23213 12223
rect 23247 12220 23259 12223
rect 23290 12220 23296 12232
rect 23247 12192 23296 12220
rect 23247 12189 23259 12192
rect 23201 12183 23259 12189
rect 23290 12180 23296 12192
rect 23348 12180 23354 12232
rect 24946 12180 24952 12232
rect 25004 12220 25010 12232
rect 25700 12229 25728 12260
rect 25225 12223 25283 12229
rect 25225 12220 25237 12223
rect 25004 12192 25237 12220
rect 25004 12180 25010 12192
rect 25225 12189 25237 12192
rect 25271 12189 25283 12223
rect 25225 12183 25283 12189
rect 25501 12223 25559 12229
rect 25501 12189 25513 12223
rect 25547 12189 25559 12223
rect 25501 12183 25559 12189
rect 25685 12223 25743 12229
rect 25685 12189 25697 12223
rect 25731 12220 25743 12223
rect 26068 12220 26096 12396
rect 31726 12288 31754 12396
rect 34146 12384 34152 12436
rect 34204 12424 34210 12436
rect 34333 12427 34391 12433
rect 34333 12424 34345 12427
rect 34204 12396 34345 12424
rect 34204 12384 34210 12396
rect 34333 12393 34345 12396
rect 34379 12393 34391 12427
rect 37093 12427 37151 12433
rect 37093 12424 37105 12427
rect 34333 12387 34391 12393
rect 36280 12396 37105 12424
rect 32674 12288 32680 12300
rect 31726 12260 32680 12288
rect 32674 12248 32680 12260
rect 32732 12248 32738 12300
rect 25731 12192 26096 12220
rect 25731 12189 25743 12192
rect 25685 12183 25743 12189
rect 22520 12124 22784 12152
rect 22520 12112 22526 12124
rect 24854 12112 24860 12164
rect 24912 12152 24918 12164
rect 25516 12152 25544 12183
rect 26142 12180 26148 12232
rect 26200 12220 26206 12232
rect 26513 12223 26571 12229
rect 26513 12220 26525 12223
rect 26200 12192 26525 12220
rect 26200 12180 26206 12192
rect 26513 12189 26525 12192
rect 26559 12220 26571 12223
rect 31754 12220 31760 12232
rect 26559 12192 31760 12220
rect 26559 12189 26571 12192
rect 26513 12183 26571 12189
rect 31754 12180 31760 12192
rect 31812 12180 31818 12232
rect 33778 12220 33784 12232
rect 33739 12192 33784 12220
rect 33778 12180 33784 12192
rect 33836 12180 33842 12232
rect 34149 12223 34207 12229
rect 34149 12189 34161 12223
rect 34195 12220 34207 12223
rect 35710 12220 35716 12232
rect 34195 12192 35716 12220
rect 34195 12189 34207 12192
rect 34149 12183 34207 12189
rect 35710 12180 35716 12192
rect 35768 12220 35774 12232
rect 36280 12229 36308 12396
rect 37093 12393 37105 12396
rect 37139 12424 37151 12427
rect 37642 12424 37648 12436
rect 37139 12396 37648 12424
rect 37139 12393 37151 12396
rect 37093 12387 37151 12393
rect 37642 12384 37648 12396
rect 37700 12384 37706 12436
rect 40957 12427 41015 12433
rect 40957 12393 40969 12427
rect 41003 12424 41015 12427
rect 41782 12424 41788 12436
rect 41003 12396 41788 12424
rect 41003 12393 41015 12396
rect 40957 12387 41015 12393
rect 41782 12384 41788 12396
rect 41840 12384 41846 12436
rect 42794 12424 42800 12436
rect 42755 12396 42800 12424
rect 42794 12384 42800 12396
rect 42852 12384 42858 12436
rect 42886 12384 42892 12436
rect 42944 12424 42950 12436
rect 43165 12427 43223 12433
rect 43165 12424 43177 12427
rect 42944 12396 43177 12424
rect 42944 12384 42950 12396
rect 43165 12393 43177 12396
rect 43211 12393 43223 12427
rect 43165 12387 43223 12393
rect 43901 12427 43959 12433
rect 43901 12393 43913 12427
rect 43947 12424 43959 12427
rect 44174 12424 44180 12436
rect 43947 12396 44180 12424
rect 43947 12393 43959 12396
rect 43901 12387 43959 12393
rect 44174 12384 44180 12396
rect 44232 12384 44238 12436
rect 36446 12356 36452 12368
rect 36407 12328 36452 12356
rect 36446 12316 36452 12328
rect 36504 12316 36510 12368
rect 44085 12359 44143 12365
rect 44085 12325 44097 12359
rect 44131 12325 44143 12359
rect 47946 12356 47952 12368
rect 44085 12319 44143 12325
rect 46492 12328 47952 12356
rect 36354 12248 36360 12300
rect 36412 12288 36418 12300
rect 36541 12291 36599 12297
rect 36541 12288 36553 12291
rect 36412 12260 36553 12288
rect 36412 12248 36418 12260
rect 36541 12257 36553 12260
rect 36587 12257 36599 12291
rect 37274 12288 37280 12300
rect 36541 12251 36599 12257
rect 37016 12260 37280 12288
rect 37016 12229 37044 12260
rect 37274 12248 37280 12260
rect 37332 12248 37338 12300
rect 41230 12248 41236 12300
rect 41288 12288 41294 12300
rect 44100 12288 44128 12319
rect 46492 12297 46520 12328
rect 47946 12316 47952 12328
rect 48004 12316 48010 12368
rect 41288 12260 44128 12288
rect 46477 12291 46535 12297
rect 41288 12248 41294 12260
rect 36265 12223 36323 12229
rect 35768 12192 36216 12220
rect 35768 12180 35774 12192
rect 24912 12124 25544 12152
rect 26780 12155 26838 12161
rect 24912 12112 24918 12124
rect 26780 12121 26792 12155
rect 26826 12152 26838 12155
rect 27798 12152 27804 12164
rect 26826 12124 27804 12152
rect 26826 12121 26838 12124
rect 26780 12115 26838 12121
rect 27798 12112 27804 12124
rect 27856 12112 27862 12164
rect 33962 12152 33968 12164
rect 33923 12124 33968 12152
rect 33962 12112 33968 12124
rect 34020 12112 34026 12164
rect 34057 12155 34115 12161
rect 34057 12121 34069 12155
rect 34103 12152 34115 12155
rect 34514 12152 34520 12164
rect 34103 12124 34520 12152
rect 34103 12121 34115 12124
rect 34057 12115 34115 12121
rect 34514 12112 34520 12124
rect 34572 12112 34578 12164
rect 36188 12152 36216 12192
rect 36265 12189 36277 12223
rect 36311 12189 36323 12223
rect 36265 12183 36323 12189
rect 37001 12223 37059 12229
rect 37001 12189 37013 12223
rect 37047 12189 37059 12223
rect 37001 12183 37059 12189
rect 37185 12223 37243 12229
rect 37185 12189 37197 12223
rect 37231 12220 37243 12223
rect 38746 12220 38752 12232
rect 37231 12192 38752 12220
rect 37231 12189 37243 12192
rect 37185 12183 37243 12189
rect 38746 12180 38752 12192
rect 38804 12180 38810 12232
rect 41138 12220 41144 12232
rect 41099 12192 41144 12220
rect 41138 12180 41144 12192
rect 41196 12180 41202 12232
rect 41432 12229 41460 12260
rect 46477 12257 46489 12291
rect 46523 12257 46535 12291
rect 46477 12251 46535 12257
rect 46661 12291 46719 12297
rect 46661 12257 46673 12291
rect 46707 12288 46719 12291
rect 47118 12288 47124 12300
rect 46707 12260 47124 12288
rect 46707 12257 46719 12260
rect 46661 12251 46719 12257
rect 47118 12248 47124 12260
rect 47176 12248 47182 12300
rect 48222 12288 48228 12300
rect 48183 12260 48228 12288
rect 48222 12248 48228 12260
rect 48280 12248 48286 12300
rect 41417 12223 41475 12229
rect 41417 12189 41429 12223
rect 41463 12189 41475 12223
rect 41417 12183 41475 12189
rect 42981 12223 43039 12229
rect 42981 12189 42993 12223
rect 43027 12189 43039 12223
rect 43254 12220 43260 12232
rect 43215 12192 43260 12220
rect 42981 12183 43039 12189
rect 37090 12152 37096 12164
rect 36188 12124 37096 12152
rect 37090 12112 37096 12124
rect 37148 12112 37154 12164
rect 42996 12152 43024 12183
rect 43254 12180 43260 12192
rect 43312 12180 43318 12232
rect 43714 12152 43720 12164
rect 42996 12124 43720 12152
rect 43714 12112 43720 12124
rect 43772 12112 43778 12164
rect 22094 12084 22100 12096
rect 22055 12056 22100 12084
rect 22094 12044 22100 12056
rect 22152 12044 22158 12096
rect 22554 12084 22560 12096
rect 22515 12056 22560 12084
rect 22554 12044 22560 12056
rect 22612 12044 22618 12096
rect 25041 12087 25099 12093
rect 25041 12053 25053 12087
rect 25087 12084 25099 12087
rect 25590 12084 25596 12096
rect 25087 12056 25596 12084
rect 25087 12053 25099 12056
rect 25041 12047 25099 12053
rect 25590 12044 25596 12056
rect 25648 12044 25654 12096
rect 27522 12044 27528 12096
rect 27580 12084 27586 12096
rect 27893 12087 27951 12093
rect 27893 12084 27905 12087
rect 27580 12056 27905 12084
rect 27580 12044 27586 12056
rect 27893 12053 27905 12056
rect 27939 12053 27951 12087
rect 27893 12047 27951 12053
rect 35434 12044 35440 12096
rect 35492 12084 35498 12096
rect 36081 12087 36139 12093
rect 36081 12084 36093 12087
rect 35492 12056 36093 12084
rect 35492 12044 35498 12056
rect 36081 12053 36093 12056
rect 36127 12053 36139 12087
rect 41322 12084 41328 12096
rect 41283 12056 41328 12084
rect 36081 12047 36139 12053
rect 41322 12044 41328 12056
rect 41380 12084 41386 12096
rect 42886 12084 42892 12096
rect 41380 12056 42892 12084
rect 41380 12044 41386 12056
rect 42886 12044 42892 12056
rect 42944 12044 42950 12096
rect 43927 12087 43985 12093
rect 43927 12053 43939 12087
rect 43973 12084 43985 12087
rect 45002 12084 45008 12096
rect 43973 12056 45008 12084
rect 43973 12053 43985 12056
rect 43927 12047 43985 12053
rect 45002 12044 45008 12056
rect 45060 12044 45066 12096
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 22094 11840 22100 11892
rect 22152 11880 22158 11892
rect 22738 11880 22744 11892
rect 22152 11852 22744 11880
rect 22152 11840 22158 11852
rect 22738 11840 22744 11852
rect 22796 11880 22802 11892
rect 22796 11852 27752 11880
rect 22796 11840 22802 11852
rect 23014 11812 23020 11824
rect 22756 11784 23020 11812
rect 2038 11744 2044 11756
rect 1999 11716 2044 11744
rect 2038 11704 2044 11716
rect 2096 11704 2102 11756
rect 22462 11744 22468 11756
rect 22423 11716 22468 11744
rect 22462 11704 22468 11716
rect 22520 11704 22526 11756
rect 22756 11753 22784 11784
rect 23014 11772 23020 11784
rect 23072 11812 23078 11824
rect 24854 11812 24860 11824
rect 23072 11784 24860 11812
rect 23072 11772 23078 11784
rect 22741 11747 22799 11753
rect 22741 11713 22753 11747
rect 22787 11713 22799 11747
rect 22922 11744 22928 11756
rect 22883 11716 22928 11744
rect 22741 11707 22799 11713
rect 22922 11704 22928 11716
rect 22980 11704 22986 11756
rect 24780 11753 24808 11784
rect 24854 11772 24860 11784
rect 24912 11772 24918 11824
rect 25866 11812 25872 11824
rect 25148 11784 25872 11812
rect 25148 11756 25176 11784
rect 25866 11772 25872 11784
rect 25924 11772 25930 11824
rect 27522 11812 27528 11824
rect 27448 11784 27528 11812
rect 24489 11747 24547 11753
rect 24489 11713 24501 11747
rect 24535 11713 24547 11747
rect 24489 11707 24547 11713
rect 24765 11747 24823 11753
rect 24765 11713 24777 11747
rect 24811 11713 24823 11747
rect 24765 11707 24823 11713
rect 24949 11747 25007 11753
rect 24949 11713 24961 11747
rect 24995 11744 25007 11747
rect 25130 11744 25136 11756
rect 24995 11716 25136 11744
rect 24995 11713 25007 11716
rect 24949 11707 25007 11713
rect 2225 11679 2283 11685
rect 2225 11645 2237 11679
rect 2271 11676 2283 11679
rect 2314 11676 2320 11688
rect 2271 11648 2320 11676
rect 2271 11645 2283 11648
rect 2225 11639 2283 11645
rect 2314 11636 2320 11648
rect 2372 11636 2378 11688
rect 2774 11676 2780 11688
rect 2735 11648 2780 11676
rect 2774 11636 2780 11648
rect 2832 11636 2838 11688
rect 22480 11676 22508 11704
rect 24504 11676 24532 11707
rect 25130 11704 25136 11716
rect 25188 11704 25194 11756
rect 25590 11744 25596 11756
rect 25551 11716 25596 11744
rect 25590 11704 25596 11716
rect 25648 11704 25654 11756
rect 27154 11744 27160 11756
rect 27115 11716 27160 11744
rect 27154 11704 27160 11716
rect 27212 11704 27218 11756
rect 27246 11704 27252 11756
rect 27304 11742 27310 11756
rect 27448 11753 27476 11784
rect 27522 11772 27528 11784
rect 27580 11772 27586 11824
rect 27724 11753 27752 11852
rect 27982 11840 27988 11892
rect 28040 11880 28046 11892
rect 29917 11883 29975 11889
rect 28040 11852 29868 11880
rect 28040 11840 28046 11852
rect 29840 11812 29868 11852
rect 29917 11849 29929 11883
rect 29963 11880 29975 11883
rect 30006 11880 30012 11892
rect 29963 11852 30012 11880
rect 29963 11849 29975 11852
rect 29917 11843 29975 11849
rect 30006 11840 30012 11852
rect 30064 11880 30070 11892
rect 30837 11883 30895 11889
rect 30837 11880 30849 11883
rect 30064 11852 30849 11880
rect 30064 11840 30070 11852
rect 30837 11849 30849 11852
rect 30883 11880 30895 11883
rect 31938 11880 31944 11892
rect 30883 11852 31944 11880
rect 30883 11849 30895 11852
rect 30837 11843 30895 11849
rect 31938 11840 31944 11852
rect 31996 11840 32002 11892
rect 33962 11880 33968 11892
rect 33923 11852 33968 11880
rect 33962 11840 33968 11852
rect 34020 11840 34026 11892
rect 37274 11840 37280 11892
rect 37332 11880 37338 11892
rect 37332 11852 38424 11880
rect 37332 11840 37338 11852
rect 33594 11812 33600 11824
rect 29840 11784 30972 11812
rect 27341 11747 27399 11753
rect 27341 11742 27353 11747
rect 27304 11714 27353 11742
rect 27304 11704 27310 11714
rect 27341 11713 27353 11714
rect 27387 11713 27399 11747
rect 27341 11707 27399 11713
rect 27433 11747 27491 11753
rect 27433 11713 27445 11747
rect 27479 11713 27491 11747
rect 27433 11707 27491 11713
rect 27709 11747 27767 11753
rect 27709 11713 27721 11747
rect 27755 11713 27767 11747
rect 27709 11707 27767 11713
rect 27798 11704 27804 11756
rect 27856 11744 27862 11756
rect 27893 11747 27951 11753
rect 27893 11744 27905 11747
rect 27856 11716 27905 11744
rect 27856 11704 27862 11716
rect 27893 11713 27905 11716
rect 27939 11713 27951 11747
rect 28626 11744 28632 11756
rect 28587 11716 28632 11744
rect 27893 11707 27951 11713
rect 28626 11704 28632 11716
rect 28684 11704 28690 11756
rect 28810 11744 28816 11756
rect 28771 11716 28816 11744
rect 28810 11704 28816 11716
rect 28868 11704 28874 11756
rect 28994 11744 29000 11756
rect 28955 11716 29000 11744
rect 28994 11704 29000 11716
rect 29052 11704 29058 11756
rect 29086 11704 29092 11756
rect 29144 11744 29150 11756
rect 29549 11747 29607 11753
rect 29549 11744 29561 11747
rect 29144 11716 29561 11744
rect 29144 11704 29150 11716
rect 29549 11713 29561 11716
rect 29595 11713 29607 11747
rect 29730 11744 29736 11756
rect 29691 11716 29736 11744
rect 29549 11707 29607 11713
rect 29730 11704 29736 11716
rect 29788 11704 29794 11756
rect 29840 11744 29868 11784
rect 29914 11744 29920 11756
rect 29840 11716 29920 11744
rect 29914 11704 29920 11716
rect 29972 11744 29978 11756
rect 30009 11747 30067 11753
rect 30009 11744 30021 11747
rect 29972 11716 30021 11744
rect 29972 11704 29978 11716
rect 30009 11713 30021 11716
rect 30055 11713 30067 11747
rect 30650 11744 30656 11756
rect 30611 11716 30656 11744
rect 30009 11707 30067 11713
rect 30650 11704 30656 11716
rect 30708 11704 30714 11756
rect 30944 11753 30972 11784
rect 31726 11784 33600 11812
rect 30929 11747 30987 11753
rect 30929 11713 30941 11747
rect 30975 11713 30987 11747
rect 30929 11707 30987 11713
rect 24854 11676 24860 11688
rect 22480 11648 24860 11676
rect 24854 11636 24860 11648
rect 24912 11636 24918 11688
rect 25869 11679 25927 11685
rect 25869 11645 25881 11679
rect 25915 11645 25927 11679
rect 25869 11639 25927 11645
rect 27525 11679 27583 11685
rect 27525 11645 27537 11679
rect 27571 11676 27583 11679
rect 31726 11676 31754 11784
rect 33594 11772 33600 11784
rect 33652 11812 33658 11824
rect 33652 11784 34008 11812
rect 33652 11772 33658 11784
rect 32030 11704 32036 11756
rect 32088 11744 32094 11756
rect 32769 11747 32827 11753
rect 32769 11744 32781 11747
rect 32088 11716 32781 11744
rect 32088 11704 32094 11716
rect 32769 11713 32781 11716
rect 32815 11713 32827 11747
rect 33778 11744 33784 11756
rect 33739 11716 33784 11744
rect 32769 11707 32827 11713
rect 33778 11704 33784 11716
rect 33836 11704 33842 11756
rect 33980 11753 34008 11784
rect 36354 11772 36360 11824
rect 36412 11812 36418 11824
rect 37645 11815 37703 11821
rect 37645 11812 37657 11815
rect 36412 11784 37657 11812
rect 36412 11772 36418 11784
rect 37645 11781 37657 11784
rect 37691 11781 37703 11815
rect 37645 11775 37703 11781
rect 38396 11756 38424 11852
rect 41138 11840 41144 11892
rect 41196 11880 41202 11892
rect 43073 11883 43131 11889
rect 43073 11880 43085 11883
rect 41196 11852 43085 11880
rect 41196 11840 41202 11852
rect 43073 11849 43085 11852
rect 43119 11849 43131 11883
rect 43073 11843 43131 11849
rect 44726 11812 44732 11824
rect 43732 11784 44732 11812
rect 33965 11747 34023 11753
rect 33965 11713 33977 11747
rect 34011 11713 34023 11747
rect 33965 11707 34023 11713
rect 35894 11704 35900 11756
rect 35952 11744 35958 11756
rect 36449 11747 36507 11753
rect 36449 11744 36461 11747
rect 35952 11716 36461 11744
rect 35952 11704 35958 11716
rect 36449 11713 36461 11716
rect 36495 11713 36507 11747
rect 37461 11747 37519 11753
rect 37461 11744 37473 11747
rect 36449 11707 36507 11713
rect 36924 11716 37473 11744
rect 27571 11648 31754 11676
rect 27571 11645 27583 11648
rect 27525 11639 27583 11645
rect 25038 11568 25044 11620
rect 25096 11608 25102 11620
rect 25884 11608 25912 11639
rect 31846 11636 31852 11688
rect 31904 11676 31910 11688
rect 32493 11679 32551 11685
rect 32493 11676 32505 11679
rect 31904 11648 32505 11676
rect 31904 11636 31910 11648
rect 32493 11645 32505 11648
rect 32539 11645 32551 11679
rect 32493 11639 32551 11645
rect 32585 11679 32643 11685
rect 32585 11645 32597 11679
rect 32631 11645 32643 11679
rect 32585 11639 32643 11645
rect 32677 11679 32735 11685
rect 32677 11645 32689 11679
rect 32723 11676 32735 11679
rect 36722 11676 36728 11688
rect 32723 11648 36728 11676
rect 32723 11645 32735 11648
rect 32677 11639 32735 11645
rect 25958 11608 25964 11620
rect 25096 11580 25820 11608
rect 25871 11580 25964 11608
rect 25096 11568 25102 11580
rect 25792 11552 25820 11580
rect 25958 11568 25964 11580
rect 26016 11608 26022 11620
rect 32398 11608 32404 11620
rect 26016 11580 32404 11608
rect 26016 11568 26022 11580
rect 32398 11568 32404 11580
rect 32456 11568 32462 11620
rect 32600 11552 32628 11639
rect 36722 11636 36728 11648
rect 36780 11636 36786 11688
rect 36924 11685 36952 11716
rect 37461 11713 37473 11716
rect 37507 11744 37519 11747
rect 38010 11744 38016 11756
rect 37507 11716 38016 11744
rect 37507 11713 37519 11716
rect 37461 11707 37519 11713
rect 38010 11704 38016 11716
rect 38068 11704 38074 11756
rect 38378 11744 38384 11756
rect 38339 11716 38384 11744
rect 38378 11704 38384 11716
rect 38436 11704 38442 11756
rect 42705 11747 42763 11753
rect 42705 11713 42717 11747
rect 42751 11744 42763 11747
rect 43070 11744 43076 11756
rect 42751 11716 43076 11744
rect 42751 11713 42763 11716
rect 42705 11707 42763 11713
rect 43070 11704 43076 11716
rect 43128 11704 43134 11756
rect 43622 11744 43628 11756
rect 43535 11716 43628 11744
rect 36909 11679 36967 11685
rect 36909 11645 36921 11679
rect 36955 11645 36967 11679
rect 36909 11639 36967 11645
rect 38657 11679 38715 11685
rect 38657 11645 38669 11679
rect 38703 11676 38715 11679
rect 38930 11676 38936 11688
rect 38703 11648 38936 11676
rect 38703 11645 38715 11648
rect 38657 11639 38715 11645
rect 38930 11636 38936 11648
rect 38988 11636 38994 11688
rect 42794 11676 42800 11688
rect 42755 11648 42800 11676
rect 42794 11636 42800 11648
rect 42852 11676 42858 11688
rect 43254 11676 43260 11688
rect 42852 11648 43260 11676
rect 42852 11636 42858 11648
rect 43254 11636 43260 11648
rect 43312 11636 43318 11688
rect 43548 11608 43576 11716
rect 43622 11704 43628 11716
rect 43680 11704 43686 11756
rect 43732 11753 43760 11784
rect 44726 11772 44732 11784
rect 44784 11772 44790 11824
rect 43717 11747 43775 11753
rect 43717 11713 43729 11747
rect 43763 11713 43775 11747
rect 43717 11707 43775 11713
rect 44450 11704 44456 11756
rect 44508 11744 44514 11756
rect 44545 11747 44603 11753
rect 44545 11744 44557 11747
rect 44508 11716 44557 11744
rect 44508 11704 44514 11716
rect 44545 11713 44557 11716
rect 44591 11713 44603 11747
rect 44545 11707 44603 11713
rect 44821 11747 44879 11753
rect 44821 11713 44833 11747
rect 44867 11744 44879 11747
rect 44910 11744 44916 11756
rect 44867 11716 44916 11744
rect 44867 11713 44879 11716
rect 44821 11707 44879 11713
rect 44910 11704 44916 11716
rect 44968 11704 44974 11756
rect 43901 11679 43959 11685
rect 43901 11645 43913 11679
rect 43947 11676 43959 11679
rect 44468 11676 44496 11704
rect 43947 11648 44496 11676
rect 43947 11645 43959 11648
rect 43901 11639 43959 11645
rect 44637 11611 44695 11617
rect 44637 11608 44649 11611
rect 42904 11580 44649 11608
rect 22281 11543 22339 11549
rect 22281 11509 22293 11543
rect 22327 11540 22339 11543
rect 22646 11540 22652 11552
rect 22327 11512 22652 11540
rect 22327 11509 22339 11512
rect 22281 11503 22339 11509
rect 22646 11500 22652 11512
rect 22704 11500 22710 11552
rect 24305 11543 24363 11549
rect 24305 11509 24317 11543
rect 24351 11540 24363 11543
rect 24762 11540 24768 11552
rect 24351 11512 24768 11540
rect 24351 11509 24363 11512
rect 24305 11503 24363 11509
rect 24762 11500 24768 11512
rect 24820 11500 24826 11552
rect 25406 11540 25412 11552
rect 25367 11512 25412 11540
rect 25406 11500 25412 11512
rect 25464 11500 25470 11552
rect 25774 11540 25780 11552
rect 25735 11512 25780 11540
rect 25774 11500 25780 11512
rect 25832 11500 25838 11552
rect 25866 11500 25872 11552
rect 25924 11540 25930 11552
rect 27706 11540 27712 11552
rect 25924 11512 27712 11540
rect 25924 11500 25930 11512
rect 27706 11500 27712 11512
rect 27764 11500 27770 11552
rect 30469 11543 30527 11549
rect 30469 11509 30481 11543
rect 30515 11540 30527 11543
rect 32122 11540 32128 11552
rect 30515 11512 32128 11540
rect 30515 11509 30527 11512
rect 30469 11503 30527 11509
rect 32122 11500 32128 11512
rect 32180 11500 32186 11552
rect 32306 11540 32312 11552
rect 32267 11512 32312 11540
rect 32306 11500 32312 11512
rect 32364 11500 32370 11552
rect 32582 11500 32588 11552
rect 32640 11500 32646 11552
rect 36446 11500 36452 11552
rect 36504 11540 36510 11552
rect 36541 11543 36599 11549
rect 36541 11540 36553 11543
rect 36504 11512 36553 11540
rect 36504 11500 36510 11512
rect 36541 11509 36553 11512
rect 36587 11509 36599 11543
rect 37826 11540 37832 11552
rect 37787 11512 37832 11540
rect 36541 11503 36599 11509
rect 37826 11500 37832 11512
rect 37884 11500 37890 11552
rect 38286 11500 38292 11552
rect 38344 11540 38350 11552
rect 38473 11543 38531 11549
rect 38473 11540 38485 11543
rect 38344 11512 38485 11540
rect 38344 11500 38350 11512
rect 38473 11509 38485 11512
rect 38519 11509 38531 11543
rect 38473 11503 38531 11509
rect 38562 11500 38568 11552
rect 38620 11540 38626 11552
rect 42904 11549 42932 11580
rect 44637 11577 44649 11580
rect 44683 11577 44695 11611
rect 44637 11571 44695 11577
rect 44726 11568 44732 11620
rect 44784 11608 44790 11620
rect 44784 11580 44829 11608
rect 44784 11568 44790 11580
rect 42889 11543 42947 11549
rect 38620 11512 38665 11540
rect 38620 11500 38626 11512
rect 42889 11509 42901 11543
rect 42935 11509 42947 11543
rect 42889 11503 42947 11509
rect 43809 11543 43867 11549
rect 43809 11509 43821 11543
rect 43855 11540 43867 11543
rect 44174 11540 44180 11552
rect 43855 11512 44180 11540
rect 43855 11509 43867 11512
rect 43809 11503 43867 11509
rect 44174 11500 44180 11512
rect 44232 11500 44238 11552
rect 44361 11543 44419 11549
rect 44361 11509 44373 11543
rect 44407 11540 44419 11543
rect 45094 11540 45100 11552
rect 44407 11512 45100 11540
rect 44407 11509 44419 11512
rect 44361 11503 44419 11509
rect 45094 11500 45100 11512
rect 45152 11500 45158 11552
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 2314 11336 2320 11348
rect 2275 11308 2320 11336
rect 2314 11296 2320 11308
rect 2372 11296 2378 11348
rect 23290 11296 23296 11348
rect 23348 11336 23354 11348
rect 23348 11308 27660 11336
rect 23348 11296 23354 11308
rect 25958 11228 25964 11280
rect 26016 11268 26022 11280
rect 26053 11271 26111 11277
rect 26053 11268 26065 11271
rect 26016 11240 26065 11268
rect 26016 11228 26022 11240
rect 26053 11237 26065 11240
rect 26099 11237 26111 11271
rect 26053 11231 26111 11237
rect 20714 11160 20720 11212
rect 20772 11200 20778 11212
rect 21818 11200 21824 11212
rect 20772 11172 21824 11200
rect 20772 11160 20778 11172
rect 21818 11160 21824 11172
rect 21876 11200 21882 11212
rect 21913 11203 21971 11209
rect 21913 11200 21925 11203
rect 21876 11172 21925 11200
rect 21876 11160 21882 11172
rect 21913 11169 21925 11172
rect 21959 11169 21971 11203
rect 21913 11163 21971 11169
rect 2222 11132 2228 11144
rect 2183 11104 2228 11132
rect 2222 11092 2228 11104
rect 2280 11092 2286 11144
rect 3050 11132 3056 11144
rect 3011 11104 3056 11132
rect 3050 11092 3056 11104
rect 3108 11092 3114 11144
rect 3786 11092 3792 11144
rect 3844 11132 3850 11144
rect 3973 11135 4031 11141
rect 3973 11132 3985 11135
rect 3844 11104 3985 11132
rect 3844 11092 3850 11104
rect 3973 11101 3985 11104
rect 4019 11132 4031 11135
rect 12529 11135 12587 11141
rect 4019 11104 6914 11132
rect 4019 11101 4031 11104
rect 3973 11095 4031 11101
rect 6886 11064 6914 11104
rect 12529 11101 12541 11135
rect 12575 11132 12587 11135
rect 12618 11132 12624 11144
rect 12575 11104 12624 11132
rect 12575 11101 12587 11104
rect 12529 11095 12587 11101
rect 12618 11092 12624 11104
rect 12676 11092 12682 11144
rect 12989 11135 13047 11141
rect 12989 11101 13001 11135
rect 13035 11101 13047 11135
rect 12989 11095 13047 11101
rect 24673 11135 24731 11141
rect 24673 11101 24685 11135
rect 24719 11132 24731 11135
rect 26142 11132 26148 11144
rect 24719 11104 26148 11132
rect 24719 11101 24731 11104
rect 24673 11095 24731 11101
rect 13004 11064 13032 11095
rect 26142 11092 26148 11104
rect 26200 11092 26206 11144
rect 27522 11132 27528 11144
rect 27483 11104 27528 11132
rect 27522 11092 27528 11104
rect 27580 11092 27586 11144
rect 27632 11132 27660 11308
rect 28994 11296 29000 11348
rect 29052 11336 29058 11348
rect 29825 11339 29883 11345
rect 29825 11336 29837 11339
rect 29052 11308 29837 11336
rect 29052 11296 29058 11308
rect 29825 11305 29837 11308
rect 29871 11305 29883 11339
rect 29825 11299 29883 11305
rect 31662 11296 31668 11348
rect 31720 11336 31726 11348
rect 32401 11339 32459 11345
rect 32401 11336 32413 11339
rect 31720 11308 32413 11336
rect 31720 11296 31726 11308
rect 32401 11305 32413 11308
rect 32447 11305 32459 11339
rect 32401 11299 32459 11305
rect 36354 11296 36360 11348
rect 36412 11336 36418 11348
rect 36909 11339 36967 11345
rect 36909 11336 36921 11339
rect 36412 11308 36921 11336
rect 36412 11296 36418 11308
rect 36909 11305 36921 11308
rect 36955 11305 36967 11339
rect 39114 11336 39120 11348
rect 36909 11299 36967 11305
rect 37752 11308 39120 11336
rect 32122 11228 32128 11280
rect 32180 11268 32186 11280
rect 32180 11240 35296 11268
rect 32180 11228 32186 11240
rect 28718 11200 28724 11212
rect 28460 11172 28724 11200
rect 27709 11135 27767 11141
rect 27709 11132 27721 11135
rect 27632 11104 27721 11132
rect 27709 11101 27721 11104
rect 27755 11132 27767 11135
rect 28353 11135 28411 11141
rect 28353 11132 28365 11135
rect 27755 11104 28365 11132
rect 27755 11101 27767 11104
rect 27709 11095 27767 11101
rect 28353 11101 28365 11104
rect 28399 11101 28411 11135
rect 28353 11095 28411 11101
rect 6886 11036 13032 11064
rect 22180 11067 22238 11073
rect 22180 11033 22192 11067
rect 22226 11064 22238 11067
rect 22462 11064 22468 11076
rect 22226 11036 22468 11064
rect 22226 11033 22238 11036
rect 22180 11027 22238 11033
rect 22462 11024 22468 11036
rect 22520 11024 22526 11076
rect 24940 11067 24998 11073
rect 24940 11033 24952 11067
rect 24986 11064 24998 11067
rect 25406 11064 25412 11076
rect 24986 11036 25412 11064
rect 24986 11033 24998 11036
rect 24940 11027 24998 11033
rect 25406 11024 25412 11036
rect 25464 11024 25470 11076
rect 27540 11064 27568 11092
rect 28169 11067 28227 11073
rect 28169 11064 28181 11067
rect 27540 11036 28181 11064
rect 28169 11033 28181 11036
rect 28215 11033 28227 11067
rect 28169 11027 28227 11033
rect 2866 10956 2872 11008
rect 2924 10996 2930 11008
rect 4065 10999 4123 11005
rect 4065 10996 4077 10999
rect 2924 10968 4077 10996
rect 2924 10956 2930 10968
rect 4065 10965 4077 10968
rect 4111 10965 4123 10999
rect 4065 10959 4123 10965
rect 12526 10956 12532 11008
rect 12584 10996 12590 11008
rect 13081 10999 13139 11005
rect 13081 10996 13093 10999
rect 12584 10968 13093 10996
rect 12584 10956 12590 10968
rect 13081 10965 13093 10968
rect 13127 10965 13139 10999
rect 23290 10996 23296 11008
rect 23251 10968 23296 10996
rect 13081 10959 13139 10965
rect 23290 10956 23296 10968
rect 23348 10956 23354 11008
rect 27709 10999 27767 11005
rect 27709 10965 27721 10999
rect 27755 10996 27767 10999
rect 28460 10996 28488 11172
rect 28718 11160 28724 11172
rect 28776 11200 28782 11212
rect 34514 11200 34520 11212
rect 28776 11172 29224 11200
rect 28776 11160 28782 11172
rect 29196 11144 29224 11172
rect 33152 11172 34520 11200
rect 28537 11135 28595 11141
rect 28537 11101 28549 11135
rect 28583 11132 28595 11135
rect 28997 11135 29055 11141
rect 28997 11132 29009 11135
rect 28583 11104 29009 11132
rect 28583 11101 28595 11104
rect 28537 11095 28595 11101
rect 28997 11101 29009 11104
rect 29043 11101 29055 11135
rect 28997 11095 29055 11101
rect 29178 11092 29184 11144
rect 29236 11132 29242 11144
rect 29730 11132 29736 11144
rect 29236 11104 29329 11132
rect 29691 11104 29736 11132
rect 29236 11092 29242 11104
rect 29730 11092 29736 11104
rect 29788 11092 29794 11144
rect 30006 11132 30012 11144
rect 29967 11104 30012 11132
rect 30006 11092 30012 11104
rect 30064 11092 30070 11144
rect 31021 11135 31079 11141
rect 31021 11101 31033 11135
rect 31067 11132 31079 11135
rect 31754 11132 31760 11144
rect 31067 11104 31760 11132
rect 31067 11101 31079 11104
rect 31021 11095 31079 11101
rect 31754 11092 31760 11104
rect 31812 11132 31818 11144
rect 32858 11132 32864 11144
rect 31812 11104 32864 11132
rect 31812 11092 31818 11104
rect 32858 11092 32864 11104
rect 32916 11092 32922 11144
rect 33152 11141 33180 11172
rect 33796 11141 33824 11172
rect 34514 11160 34520 11172
rect 34572 11160 34578 11212
rect 33137 11135 33195 11141
rect 33137 11101 33149 11135
rect 33183 11101 33195 11135
rect 33137 11095 33195 11101
rect 33321 11135 33379 11141
rect 33321 11101 33333 11135
rect 33367 11101 33379 11135
rect 33321 11095 33379 11101
rect 33781 11135 33839 11141
rect 33781 11101 33793 11135
rect 33827 11101 33839 11135
rect 33781 11095 33839 11101
rect 33965 11135 34023 11141
rect 33965 11101 33977 11135
rect 34011 11101 34023 11135
rect 33965 11095 34023 11101
rect 29089 11067 29147 11073
rect 29089 11033 29101 11067
rect 29135 11064 29147 11067
rect 29748 11064 29776 11092
rect 29914 11064 29920 11076
rect 29135 11036 29776 11064
rect 29875 11036 29920 11064
rect 29135 11033 29147 11036
rect 29089 11027 29147 11033
rect 29914 11024 29920 11036
rect 29972 11024 29978 11076
rect 31288 11067 31346 11073
rect 31288 11033 31300 11067
rect 31334 11064 31346 11067
rect 32306 11064 32312 11076
rect 31334 11036 32312 11064
rect 31334 11033 31346 11036
rect 31288 11027 31346 11033
rect 32306 11024 32312 11036
rect 32364 11024 32370 11076
rect 32398 11024 32404 11076
rect 32456 11064 32462 11076
rect 33336 11064 33364 11095
rect 33980 11064 34008 11095
rect 32456 11036 34008 11064
rect 35268 11064 35296 11240
rect 35802 11228 35808 11280
rect 35860 11268 35866 11280
rect 37752 11268 37780 11308
rect 39114 11296 39120 11308
rect 39172 11296 39178 11348
rect 43070 11336 43076 11348
rect 43031 11308 43076 11336
rect 43070 11296 43076 11308
rect 43128 11296 43134 11348
rect 44450 11296 44456 11348
rect 44508 11336 44514 11348
rect 44637 11339 44695 11345
rect 44637 11336 44649 11339
rect 44508 11308 44649 11336
rect 44508 11296 44514 11308
rect 44637 11305 44649 11308
rect 44683 11305 44695 11339
rect 44637 11299 44695 11305
rect 35860 11240 37780 11268
rect 37829 11271 37887 11277
rect 35860 11228 35866 11240
rect 35434 11200 35440 11212
rect 35395 11172 35440 11200
rect 35434 11160 35440 11172
rect 35492 11160 35498 11212
rect 35345 11135 35403 11141
rect 35345 11101 35357 11135
rect 35391 11132 35403 11135
rect 35894 11132 35900 11144
rect 35391 11104 35900 11132
rect 35391 11101 35403 11104
rect 35345 11095 35403 11101
rect 35894 11092 35900 11104
rect 35952 11092 35958 11144
rect 36740 11141 36768 11240
rect 37829 11237 37841 11271
rect 37875 11268 37887 11271
rect 41322 11268 41328 11280
rect 37875 11240 41328 11268
rect 37875 11237 37887 11240
rect 37829 11231 37887 11237
rect 41322 11228 41328 11240
rect 41380 11228 41386 11280
rect 38102 11160 38108 11212
rect 38160 11200 38166 11212
rect 40310 11200 40316 11212
rect 38160 11172 40316 11200
rect 38160 11160 38166 11172
rect 40310 11160 40316 11172
rect 40368 11200 40374 11212
rect 40862 11200 40868 11212
rect 40368 11172 40868 11200
rect 40368 11160 40374 11172
rect 40862 11160 40868 11172
rect 40920 11160 40926 11212
rect 43441 11203 43499 11209
rect 43441 11169 43453 11203
rect 43487 11200 43499 11203
rect 43898 11200 43904 11212
rect 43487 11172 43904 11200
rect 43487 11169 43499 11172
rect 43441 11163 43499 11169
rect 43898 11160 43904 11172
rect 43956 11160 43962 11212
rect 44269 11203 44327 11209
rect 44269 11169 44281 11203
rect 44315 11200 44327 11203
rect 45646 11200 45652 11212
rect 44315 11172 45652 11200
rect 44315 11169 44327 11172
rect 44269 11163 44327 11169
rect 45646 11160 45652 11172
rect 45704 11160 45710 11212
rect 36633 11135 36691 11141
rect 36633 11101 36645 11135
rect 36679 11101 36691 11135
rect 36633 11095 36691 11101
rect 36725 11135 36783 11141
rect 36725 11101 36737 11135
rect 36771 11101 36783 11135
rect 36725 11095 36783 11101
rect 37829 11135 37887 11141
rect 37829 11101 37841 11135
rect 37875 11132 37887 11135
rect 37918 11132 37924 11144
rect 37875 11104 37924 11132
rect 37875 11101 37887 11104
rect 37829 11095 37887 11101
rect 36648 11064 36676 11095
rect 37918 11092 37924 11104
rect 37976 11092 37982 11144
rect 38010 11092 38016 11144
rect 38068 11132 38074 11144
rect 38470 11132 38476 11144
rect 38068 11104 38113 11132
rect 38431 11104 38476 11132
rect 38068 11092 38074 11104
rect 38470 11092 38476 11104
rect 38528 11092 38534 11144
rect 38749 11135 38807 11141
rect 38749 11101 38761 11135
rect 38795 11101 38807 11135
rect 39114 11132 39120 11144
rect 39075 11104 39120 11132
rect 38749 11095 38807 11101
rect 38764 11064 38792 11095
rect 39114 11092 39120 11104
rect 39172 11092 39178 11144
rect 42978 11092 42984 11144
rect 43036 11132 43042 11144
rect 43257 11135 43315 11141
rect 43257 11132 43269 11135
rect 43036 11104 43269 11132
rect 43036 11092 43042 11104
rect 43257 11101 43269 11104
rect 43303 11101 43315 11135
rect 43257 11095 43315 11101
rect 43533 11135 43591 11141
rect 43533 11101 43545 11135
rect 43579 11101 43591 11135
rect 44450 11132 44456 11144
rect 44411 11104 44456 11132
rect 43533 11095 43591 11101
rect 35268 11036 38792 11064
rect 43548 11064 43576 11095
rect 44450 11092 44456 11104
rect 44508 11092 44514 11144
rect 45094 11092 45100 11144
rect 45152 11132 45158 11144
rect 45189 11135 45247 11141
rect 45189 11132 45201 11135
rect 45152 11104 45201 11132
rect 45152 11092 45158 11104
rect 45189 11101 45201 11104
rect 45235 11101 45247 11135
rect 45554 11132 45560 11144
rect 45515 11104 45560 11132
rect 45189 11095 45247 11101
rect 45554 11092 45560 11104
rect 45612 11092 45618 11144
rect 43548 11036 44128 11064
rect 32456 11024 32462 11036
rect 27755 10968 28488 10996
rect 27755 10965 27767 10968
rect 27709 10959 27767 10965
rect 30558 10956 30564 11008
rect 30616 10996 30622 11008
rect 32766 10996 32772 11008
rect 30616 10968 32772 10996
rect 30616 10956 30622 10968
rect 32766 10956 32772 10968
rect 32824 10956 32830 11008
rect 33134 10956 33140 11008
rect 33192 10996 33198 11008
rect 33229 10999 33287 11005
rect 33229 10996 33241 10999
rect 33192 10968 33241 10996
rect 33192 10956 33198 10968
rect 33229 10965 33241 10968
rect 33275 10965 33287 10999
rect 33229 10959 33287 10965
rect 33965 10999 34023 11005
rect 33965 10965 33977 10999
rect 34011 10996 34023 10999
rect 34054 10996 34060 11008
rect 34011 10968 34060 10996
rect 34011 10965 34023 10968
rect 33965 10959 34023 10965
rect 34054 10956 34060 10968
rect 34112 10956 34118 11008
rect 35526 10956 35532 11008
rect 35584 10996 35590 11008
rect 35713 10999 35771 11005
rect 35713 10996 35725 10999
rect 35584 10968 35725 10996
rect 35584 10956 35590 10968
rect 35713 10965 35725 10968
rect 35759 10965 35771 10999
rect 35713 10959 35771 10965
rect 38654 10956 38660 11008
rect 38712 10996 38718 11008
rect 42794 10996 42800 11008
rect 38712 10968 42800 10996
rect 38712 10956 38718 10968
rect 42794 10956 42800 10968
rect 42852 10956 42858 11008
rect 44100 10996 44128 11036
rect 44174 11024 44180 11076
rect 44232 11064 44238 11076
rect 45373 11067 45431 11073
rect 45373 11064 45385 11067
rect 44232 11036 45385 11064
rect 44232 11024 44238 11036
rect 45373 11033 45385 11036
rect 45419 11033 45431 11067
rect 45373 11027 45431 11033
rect 45465 11067 45523 11073
rect 45465 11033 45477 11067
rect 45511 11033 45523 11067
rect 45465 11027 45523 11033
rect 44910 10996 44916 11008
rect 44100 10968 44916 10996
rect 44910 10956 44916 10968
rect 44968 10996 44974 11008
rect 45480 10996 45508 11027
rect 45738 10996 45744 11008
rect 44968 10968 45508 10996
rect 45699 10968 45744 10996
rect 44968 10956 44974 10968
rect 45738 10956 45744 10968
rect 45796 10956 45802 11008
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 22462 10792 22468 10804
rect 22423 10764 22468 10792
rect 22462 10752 22468 10764
rect 22520 10752 22526 10804
rect 25317 10795 25375 10801
rect 25317 10761 25329 10795
rect 25363 10761 25375 10795
rect 25317 10755 25375 10761
rect 30009 10795 30067 10801
rect 30009 10761 30021 10795
rect 30055 10792 30067 10795
rect 30650 10792 30656 10804
rect 30055 10764 30656 10792
rect 30055 10761 30067 10764
rect 30009 10755 30067 10761
rect 2866 10724 2872 10736
rect 2827 10696 2872 10724
rect 2866 10684 2872 10696
rect 2924 10684 2930 10736
rect 12526 10724 12532 10736
rect 12487 10696 12532 10724
rect 12526 10684 12532 10696
rect 12584 10684 12590 10736
rect 25038 10684 25044 10736
rect 25096 10724 25102 10736
rect 25332 10724 25360 10755
rect 30650 10752 30656 10764
rect 30708 10752 30714 10804
rect 30926 10792 30932 10804
rect 30760 10764 30932 10792
rect 30760 10724 30788 10764
rect 30926 10752 30932 10764
rect 30984 10752 30990 10804
rect 33413 10795 33471 10801
rect 33413 10761 33425 10795
rect 33459 10792 33471 10795
rect 35802 10792 35808 10804
rect 33459 10764 35808 10792
rect 33459 10761 33471 10764
rect 33413 10755 33471 10761
rect 35802 10752 35808 10764
rect 35860 10752 35866 10804
rect 38105 10795 38163 10801
rect 38105 10792 38117 10795
rect 36556 10764 38117 10792
rect 31389 10727 31447 10733
rect 31389 10724 31401 10727
rect 25096 10696 30788 10724
rect 30852 10696 31401 10724
rect 25096 10684 25102 10696
rect 22646 10656 22652 10668
rect 22607 10628 22652 10656
rect 22646 10616 22652 10628
rect 22704 10616 22710 10668
rect 23937 10659 23995 10665
rect 23937 10656 23949 10659
rect 22848 10628 23949 10656
rect 2685 10591 2743 10597
rect 2685 10557 2697 10591
rect 2731 10588 2743 10591
rect 3050 10588 3056 10600
rect 2731 10560 3056 10588
rect 2731 10557 2743 10560
rect 2685 10551 2743 10557
rect 3050 10548 3056 10560
rect 3108 10548 3114 10600
rect 3142 10548 3148 10600
rect 3200 10588 3206 10600
rect 12345 10591 12403 10597
rect 3200 10560 3245 10588
rect 3200 10548 3206 10560
rect 12345 10557 12357 10591
rect 12391 10588 12403 10591
rect 12618 10588 12624 10600
rect 12391 10560 12624 10588
rect 12391 10557 12403 10560
rect 12345 10551 12403 10557
rect 12618 10548 12624 10560
rect 12676 10548 12682 10600
rect 14182 10588 14188 10600
rect 14143 10560 14188 10588
rect 14182 10548 14188 10560
rect 14240 10548 14246 10600
rect 21818 10548 21824 10600
rect 21876 10588 21882 10600
rect 22848 10588 22876 10628
rect 23937 10625 23949 10628
rect 23983 10625 23995 10659
rect 23937 10619 23995 10625
rect 24204 10659 24262 10665
rect 24204 10625 24216 10659
rect 24250 10656 24262 10659
rect 24578 10656 24584 10668
rect 24250 10628 24584 10656
rect 24250 10625 24262 10628
rect 24204 10619 24262 10625
rect 24578 10616 24584 10628
rect 24636 10616 24642 10668
rect 26510 10616 26516 10668
rect 26568 10656 26574 10668
rect 27157 10659 27215 10665
rect 27157 10656 27169 10659
rect 26568 10628 27169 10656
rect 26568 10616 26574 10628
rect 27157 10625 27169 10628
rect 27203 10625 27215 10659
rect 27157 10619 27215 10625
rect 27341 10659 27399 10665
rect 27341 10625 27353 10659
rect 27387 10625 27399 10659
rect 27522 10656 27528 10668
rect 27483 10628 27528 10656
rect 27341 10619 27399 10625
rect 21876 10560 22876 10588
rect 22925 10591 22983 10597
rect 21876 10548 21882 10560
rect 22925 10557 22937 10591
rect 22971 10588 22983 10591
rect 23290 10588 23296 10600
rect 22971 10560 23296 10588
rect 22971 10557 22983 10560
rect 22925 10551 22983 10557
rect 23290 10548 23296 10560
rect 23348 10548 23354 10600
rect 27356 10520 27384 10619
rect 27522 10616 27528 10628
rect 27580 10616 27586 10668
rect 27706 10656 27712 10668
rect 27667 10628 27712 10656
rect 27706 10616 27712 10628
rect 27764 10616 27770 10668
rect 28905 10659 28963 10665
rect 28905 10625 28917 10659
rect 28951 10656 28963 10659
rect 28994 10656 29000 10668
rect 28951 10628 29000 10656
rect 28951 10625 28963 10628
rect 28905 10619 28963 10625
rect 28994 10616 29000 10628
rect 29052 10616 29058 10668
rect 29089 10659 29147 10665
rect 29089 10625 29101 10659
rect 29135 10656 29147 10659
rect 29178 10656 29184 10668
rect 29135 10628 29184 10656
rect 29135 10625 29147 10628
rect 29089 10619 29147 10625
rect 29178 10616 29184 10628
rect 29236 10616 29242 10668
rect 29641 10659 29699 10665
rect 29641 10625 29653 10659
rect 29687 10656 29699 10659
rect 30558 10656 30564 10668
rect 29687 10628 30564 10656
rect 29687 10625 29699 10628
rect 29641 10619 29699 10625
rect 30558 10616 30564 10628
rect 30616 10616 30622 10668
rect 30745 10659 30803 10665
rect 30745 10625 30757 10659
rect 30791 10656 30803 10659
rect 30852 10656 30880 10696
rect 31389 10693 31401 10696
rect 31435 10724 31447 10727
rect 31478 10724 31484 10736
rect 31435 10696 31484 10724
rect 31435 10693 31447 10696
rect 31389 10687 31447 10693
rect 31478 10684 31484 10696
rect 31536 10684 31542 10736
rect 34054 10724 34060 10736
rect 32692 10696 34060 10724
rect 30791 10628 30880 10656
rect 30791 10625 30803 10628
rect 30745 10619 30803 10625
rect 30926 10616 30932 10668
rect 30984 10656 30990 10668
rect 32692 10665 32720 10696
rect 34054 10684 34060 10696
rect 34112 10684 34118 10736
rect 35526 10724 35532 10736
rect 35487 10696 35532 10724
rect 35526 10684 35532 10696
rect 35584 10684 35590 10736
rect 31573 10659 31631 10665
rect 31573 10656 31585 10659
rect 30984 10628 31585 10656
rect 30984 10616 30990 10628
rect 31573 10625 31585 10628
rect 31619 10625 31631 10659
rect 31573 10619 31631 10625
rect 32677 10659 32735 10665
rect 32677 10625 32689 10659
rect 32723 10625 32735 10659
rect 32677 10619 32735 10625
rect 32766 10616 32772 10668
rect 32824 10656 32830 10668
rect 32861 10659 32919 10665
rect 32861 10656 32873 10659
rect 32824 10628 32873 10656
rect 32824 10616 32830 10628
rect 32861 10625 32873 10628
rect 32907 10625 32919 10659
rect 32861 10619 32919 10625
rect 33045 10659 33103 10665
rect 33045 10625 33057 10659
rect 33091 10656 33103 10659
rect 33134 10656 33140 10668
rect 33091 10628 33140 10656
rect 33091 10625 33103 10628
rect 33045 10619 33103 10625
rect 33134 10616 33140 10628
rect 33192 10616 33198 10668
rect 33229 10659 33287 10665
rect 33229 10625 33241 10659
rect 33275 10625 33287 10659
rect 33229 10619 33287 10625
rect 35345 10659 35403 10665
rect 35345 10625 35357 10659
rect 35391 10625 35403 10659
rect 35618 10656 35624 10668
rect 35579 10628 35624 10656
rect 35345 10619 35403 10625
rect 27433 10591 27491 10597
rect 27433 10557 27445 10591
rect 27479 10588 27491 10591
rect 28810 10588 28816 10600
rect 27479 10560 28816 10588
rect 27479 10557 27491 10560
rect 27433 10551 27491 10557
rect 28810 10548 28816 10560
rect 28868 10548 28874 10600
rect 29730 10588 29736 10600
rect 29691 10560 29736 10588
rect 29730 10548 29736 10560
rect 29788 10548 29794 10600
rect 29914 10548 29920 10600
rect 29972 10588 29978 10600
rect 32953 10591 33011 10597
rect 32953 10588 32965 10591
rect 29972 10560 32965 10588
rect 29972 10548 29978 10560
rect 32953 10557 32965 10560
rect 32999 10557 33011 10591
rect 32953 10551 33011 10557
rect 28902 10520 28908 10532
rect 27356 10492 28908 10520
rect 28902 10480 28908 10492
rect 28960 10480 28966 10532
rect 30837 10523 30895 10529
rect 30837 10489 30849 10523
rect 30883 10520 30895 10523
rect 31938 10520 31944 10532
rect 30883 10492 31944 10520
rect 30883 10489 30895 10492
rect 30837 10483 30895 10489
rect 31938 10480 31944 10492
rect 31996 10520 32002 10532
rect 33244 10520 33272 10619
rect 35360 10588 35388 10619
rect 35618 10616 35624 10628
rect 35676 10616 35682 10668
rect 35710 10616 35716 10668
rect 35768 10656 35774 10668
rect 36556 10656 36584 10764
rect 38105 10761 38117 10764
rect 38151 10792 38163 10795
rect 38562 10792 38568 10804
rect 38151 10764 38568 10792
rect 38151 10761 38163 10764
rect 38105 10755 38163 10761
rect 38562 10752 38568 10764
rect 38620 10752 38626 10804
rect 38654 10752 38660 10804
rect 38712 10792 38718 10804
rect 38712 10764 38757 10792
rect 38856 10764 39436 10792
rect 38712 10752 38718 10764
rect 36633 10727 36691 10733
rect 36633 10693 36645 10727
rect 36679 10724 36691 10727
rect 37826 10724 37832 10736
rect 36679 10696 37832 10724
rect 36679 10693 36691 10696
rect 36633 10687 36691 10693
rect 37826 10684 37832 10696
rect 37884 10724 37890 10736
rect 37884 10696 38240 10724
rect 37884 10684 37890 10696
rect 38212 10665 38240 10696
rect 38378 10684 38384 10736
rect 38436 10724 38442 10736
rect 38856 10724 38884 10764
rect 38436 10696 38884 10724
rect 38436 10684 38442 10696
rect 36817 10659 36875 10665
rect 36817 10656 36829 10659
rect 35768 10628 35813 10656
rect 36556 10628 36829 10656
rect 35768 10616 35774 10628
rect 36817 10625 36829 10628
rect 36863 10625 36875 10659
rect 36817 10619 36875 10625
rect 36909 10659 36967 10665
rect 36909 10625 36921 10659
rect 36955 10656 36967 10659
rect 37921 10659 37979 10665
rect 37921 10656 37933 10659
rect 36955 10628 37933 10656
rect 36955 10625 36967 10628
rect 36909 10619 36967 10625
rect 37921 10625 37933 10628
rect 37967 10625 37979 10659
rect 37921 10619 37979 10625
rect 38197 10659 38255 10665
rect 38197 10625 38209 10659
rect 38243 10625 38255 10659
rect 38930 10656 38936 10668
rect 38891 10628 38936 10656
rect 38197 10619 38255 10625
rect 36722 10588 36728 10600
rect 35360 10560 36728 10588
rect 36722 10548 36728 10560
rect 36780 10548 36786 10600
rect 37936 10588 37964 10619
rect 38930 10616 38936 10628
rect 38988 10616 38994 10668
rect 39408 10665 39436 10764
rect 40126 10752 40132 10804
rect 40184 10792 40190 10804
rect 40497 10795 40555 10801
rect 40497 10792 40509 10795
rect 40184 10764 40509 10792
rect 40184 10752 40190 10764
rect 40497 10761 40509 10764
rect 40543 10792 40555 10795
rect 41046 10792 41052 10804
rect 40543 10764 41052 10792
rect 40543 10761 40555 10764
rect 40497 10755 40555 10761
rect 41046 10752 41052 10764
rect 41104 10752 41110 10804
rect 41598 10792 41604 10804
rect 41248 10764 41604 10792
rect 41248 10724 41276 10764
rect 41598 10752 41604 10764
rect 41656 10752 41662 10804
rect 44910 10752 44916 10804
rect 44968 10792 44974 10804
rect 47029 10795 47087 10801
rect 47029 10792 47041 10795
rect 44968 10764 47041 10792
rect 44968 10752 44974 10764
rect 47029 10761 47041 10764
rect 47075 10761 47087 10795
rect 47029 10755 47087 10761
rect 39776 10696 41276 10724
rect 39025 10659 39083 10665
rect 39025 10625 39037 10659
rect 39071 10656 39083 10659
rect 39393 10659 39451 10665
rect 39071 10628 39344 10656
rect 39071 10625 39083 10628
rect 39025 10619 39083 10625
rect 38470 10588 38476 10600
rect 37936 10560 38476 10588
rect 38470 10548 38476 10560
rect 38528 10548 38534 10600
rect 39117 10591 39175 10597
rect 39117 10557 39129 10591
rect 39163 10588 39175 10591
rect 39206 10588 39212 10600
rect 39163 10560 39212 10588
rect 39163 10557 39175 10560
rect 39117 10551 39175 10557
rect 39206 10548 39212 10560
rect 39264 10548 39270 10600
rect 39316 10588 39344 10628
rect 39393 10625 39405 10659
rect 39439 10625 39451 10659
rect 39393 10619 39451 10625
rect 39776 10588 39804 10696
rect 44634 10684 44640 10736
rect 44692 10724 44698 10736
rect 45370 10724 45376 10736
rect 44692 10696 45376 10724
rect 44692 10684 44698 10696
rect 40310 10656 40316 10668
rect 40271 10628 40316 10656
rect 40310 10616 40316 10628
rect 40368 10616 40374 10668
rect 40589 10659 40647 10665
rect 40589 10625 40601 10659
rect 40635 10656 40647 10659
rect 40635 10628 40715 10656
rect 40635 10625 40647 10628
rect 40589 10619 40647 10625
rect 39316 10560 39804 10588
rect 31996 10492 33272 10520
rect 37737 10523 37795 10529
rect 31996 10480 32002 10492
rect 37737 10489 37749 10523
rect 37783 10520 37795 10523
rect 38194 10520 38200 10532
rect 37783 10492 38200 10520
rect 37783 10489 37795 10492
rect 37737 10483 37795 10489
rect 38194 10480 38200 10492
rect 38252 10520 38258 10532
rect 40687 10520 40715 10628
rect 40862 10616 40868 10668
rect 40920 10656 40926 10668
rect 41049 10659 41107 10665
rect 41049 10656 41061 10659
rect 40920 10628 41061 10656
rect 40920 10616 40926 10628
rect 41049 10625 41061 10628
rect 41095 10625 41107 10659
rect 41049 10619 41107 10625
rect 41233 10659 41291 10665
rect 41233 10625 41245 10659
rect 41279 10625 41291 10659
rect 41233 10619 41291 10625
rect 41337 10659 41395 10665
rect 41337 10625 41349 10659
rect 41383 10656 41395 10659
rect 44174 10656 44180 10668
rect 41383 10625 41414 10656
rect 44135 10628 44180 10656
rect 41337 10619 41414 10625
rect 41248 10588 41276 10619
rect 40972 10560 41276 10588
rect 40972 10520 41000 10560
rect 38252 10492 41000 10520
rect 38252 10480 38258 10492
rect 41046 10480 41052 10532
rect 41104 10520 41110 10532
rect 41386 10520 41414 10619
rect 44174 10616 44180 10628
rect 44232 10616 44238 10668
rect 44361 10659 44419 10665
rect 44361 10625 44373 10659
rect 44407 10656 44419 10659
rect 44542 10656 44548 10668
rect 44407 10628 44548 10656
rect 44407 10625 44419 10628
rect 44361 10619 44419 10625
rect 44542 10616 44548 10628
rect 44600 10616 44606 10668
rect 44910 10656 44916 10668
rect 44871 10628 44916 10656
rect 44910 10616 44916 10628
rect 44968 10616 44974 10668
rect 45112 10665 45140 10696
rect 45370 10684 45376 10696
rect 45428 10684 45434 10736
rect 45738 10684 45744 10736
rect 45796 10724 45802 10736
rect 45894 10727 45952 10733
rect 45894 10724 45906 10727
rect 45796 10696 45906 10724
rect 45796 10684 45802 10696
rect 45894 10693 45906 10696
rect 45940 10693 45952 10727
rect 45894 10687 45952 10693
rect 45097 10659 45155 10665
rect 45097 10625 45109 10659
rect 45143 10625 45155 10659
rect 45097 10619 45155 10625
rect 45186 10616 45192 10668
rect 45244 10656 45250 10668
rect 45649 10659 45707 10665
rect 45649 10656 45661 10659
rect 45244 10628 45661 10656
rect 45244 10616 45250 10628
rect 45649 10625 45661 10628
rect 45695 10625 45707 10659
rect 45649 10619 45707 10625
rect 44082 10588 44088 10600
rect 44043 10560 44088 10588
rect 44082 10548 44088 10560
rect 44140 10548 44146 10600
rect 44269 10591 44327 10597
rect 44269 10557 44281 10591
rect 44315 10588 44327 10591
rect 44450 10588 44456 10600
rect 44315 10560 44456 10588
rect 44315 10557 44327 10560
rect 44269 10551 44327 10557
rect 44450 10548 44456 10560
rect 44508 10588 44514 10600
rect 44818 10588 44824 10600
rect 44508 10560 44824 10588
rect 44508 10548 44514 10560
rect 44818 10548 44824 10560
rect 44876 10548 44882 10600
rect 41104 10492 41414 10520
rect 41104 10480 41110 10492
rect 42610 10480 42616 10532
rect 42668 10520 42674 10532
rect 45204 10520 45232 10616
rect 42668 10492 45232 10520
rect 42668 10480 42674 10492
rect 22738 10412 22744 10464
rect 22796 10452 22802 10464
rect 22833 10455 22891 10461
rect 22833 10452 22845 10455
rect 22796 10424 22845 10452
rect 22796 10412 22802 10424
rect 22833 10421 22845 10424
rect 22879 10421 22891 10455
rect 27890 10452 27896 10464
rect 27851 10424 27896 10452
rect 22833 10415 22891 10421
rect 27890 10412 27896 10424
rect 27948 10412 27954 10464
rect 28994 10452 29000 10464
rect 28955 10424 29000 10452
rect 28994 10412 29000 10424
rect 29052 10412 29058 10464
rect 29822 10452 29828 10464
rect 29783 10424 29828 10452
rect 29822 10412 29828 10424
rect 29880 10412 29886 10464
rect 31757 10455 31815 10461
rect 31757 10421 31769 10455
rect 31803 10452 31815 10455
rect 32122 10452 32128 10464
rect 31803 10424 32128 10452
rect 31803 10421 31815 10424
rect 31757 10415 31815 10421
rect 32122 10412 32128 10424
rect 32180 10412 32186 10464
rect 35894 10452 35900 10464
rect 35855 10424 35900 10452
rect 35894 10412 35900 10424
rect 35952 10412 35958 10464
rect 36906 10452 36912 10464
rect 36867 10424 36912 10452
rect 36906 10412 36912 10424
rect 36964 10412 36970 10464
rect 38286 10412 38292 10464
rect 38344 10452 38350 10464
rect 39209 10455 39267 10461
rect 39209 10452 39221 10455
rect 38344 10424 39221 10452
rect 38344 10412 38350 10424
rect 39209 10421 39221 10424
rect 39255 10421 39267 10455
rect 39209 10415 39267 10421
rect 40129 10455 40187 10461
rect 40129 10421 40141 10455
rect 40175 10452 40187 10455
rect 40402 10452 40408 10464
rect 40175 10424 40408 10452
rect 40175 10421 40187 10424
rect 40129 10415 40187 10421
rect 40402 10412 40408 10424
rect 40460 10412 40466 10464
rect 41138 10452 41144 10464
rect 41099 10424 41144 10452
rect 41138 10412 41144 10424
rect 41196 10412 41202 10464
rect 43530 10412 43536 10464
rect 43588 10452 43594 10464
rect 43901 10455 43959 10461
rect 43901 10452 43913 10455
rect 43588 10424 43913 10452
rect 43588 10412 43594 10424
rect 43901 10421 43913 10424
rect 43947 10421 43959 10455
rect 43901 10415 43959 10421
rect 44818 10412 44824 10464
rect 44876 10452 44882 10464
rect 45005 10455 45063 10461
rect 45005 10452 45017 10455
rect 44876 10424 45017 10452
rect 44876 10412 44882 10424
rect 45005 10421 45017 10424
rect 45051 10421 45063 10455
rect 45005 10415 45063 10421
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 24578 10248 24584 10260
rect 24539 10220 24584 10248
rect 24578 10208 24584 10220
rect 24636 10208 24642 10260
rect 27525 10251 27583 10257
rect 27525 10217 27537 10251
rect 27571 10248 27583 10251
rect 27706 10248 27712 10260
rect 27571 10220 27712 10248
rect 27571 10217 27583 10220
rect 27525 10211 27583 10217
rect 27706 10208 27712 10220
rect 27764 10208 27770 10260
rect 28997 10251 29055 10257
rect 28997 10217 29009 10251
rect 29043 10248 29055 10251
rect 29086 10248 29092 10260
rect 29043 10220 29092 10248
rect 29043 10217 29055 10220
rect 28997 10211 29055 10217
rect 29086 10208 29092 10220
rect 29144 10208 29150 10260
rect 29733 10251 29791 10257
rect 29733 10217 29745 10251
rect 29779 10248 29791 10251
rect 29914 10248 29920 10260
rect 29779 10220 29920 10248
rect 29779 10217 29791 10220
rect 29733 10211 29791 10217
rect 29914 10208 29920 10220
rect 29972 10208 29978 10260
rect 30929 10251 30987 10257
rect 30929 10217 30941 10251
rect 30975 10248 30987 10251
rect 32582 10248 32588 10260
rect 30975 10220 32588 10248
rect 30975 10217 30987 10220
rect 30929 10211 30987 10217
rect 32582 10208 32588 10220
rect 32640 10208 32646 10260
rect 33321 10251 33379 10257
rect 33321 10217 33333 10251
rect 33367 10248 33379 10251
rect 33778 10248 33784 10260
rect 33367 10220 33784 10248
rect 33367 10217 33379 10220
rect 33321 10211 33379 10217
rect 33778 10208 33784 10220
rect 33836 10208 33842 10260
rect 35618 10208 35624 10260
rect 35676 10248 35682 10260
rect 36265 10251 36323 10257
rect 36265 10248 36277 10251
rect 35676 10220 36277 10248
rect 35676 10208 35682 10220
rect 36265 10217 36277 10220
rect 36311 10248 36323 10251
rect 38286 10248 38292 10260
rect 36311 10220 38292 10248
rect 36311 10217 36323 10220
rect 36265 10211 36323 10217
rect 38286 10208 38292 10220
rect 38344 10208 38350 10260
rect 40862 10208 40868 10260
rect 40920 10248 40926 10260
rect 42153 10251 42211 10257
rect 42153 10248 42165 10251
rect 40920 10220 42165 10248
rect 40920 10208 40926 10220
rect 42153 10217 42165 10220
rect 42199 10217 42211 10251
rect 42153 10211 42211 10217
rect 45557 10251 45615 10257
rect 45557 10217 45569 10251
rect 45603 10248 45615 10251
rect 45646 10248 45652 10260
rect 45603 10220 45652 10248
rect 45603 10217 45615 10220
rect 45557 10211 45615 10217
rect 45646 10208 45652 10220
rect 45704 10208 45710 10260
rect 22830 10140 22836 10192
rect 22888 10180 22894 10192
rect 24949 10183 25007 10189
rect 24949 10180 24961 10183
rect 22888 10152 24961 10180
rect 22888 10140 22894 10152
rect 24949 10149 24961 10152
rect 24995 10180 25007 10183
rect 25774 10180 25780 10192
rect 24995 10152 25780 10180
rect 24995 10149 25007 10152
rect 24949 10143 25007 10149
rect 25774 10140 25780 10152
rect 25832 10140 25838 10192
rect 21818 10112 21824 10124
rect 21779 10084 21824 10112
rect 21818 10072 21824 10084
rect 21876 10072 21882 10124
rect 25038 10112 25044 10124
rect 24999 10084 25044 10112
rect 25038 10072 25044 10084
rect 25096 10072 25102 10124
rect 26142 10112 26148 10124
rect 26103 10084 26148 10112
rect 26142 10072 26148 10084
rect 26200 10072 26206 10124
rect 27724 10112 27752 10208
rect 29181 10183 29239 10189
rect 29181 10149 29193 10183
rect 29227 10180 29239 10183
rect 30834 10180 30840 10192
rect 29227 10152 30840 10180
rect 29227 10149 29239 10152
rect 29181 10143 29239 10149
rect 30834 10140 30840 10152
rect 30892 10140 30898 10192
rect 31849 10183 31907 10189
rect 31849 10180 31861 10183
rect 31036 10152 31861 10180
rect 28077 10115 28135 10121
rect 27724 10084 28028 10112
rect 2038 10004 2044 10056
rect 2096 10044 2102 10056
rect 2317 10047 2375 10053
rect 2317 10044 2329 10047
rect 2096 10016 2329 10044
rect 2096 10004 2102 10016
rect 2317 10013 2329 10016
rect 2363 10013 2375 10047
rect 24762 10044 24768 10056
rect 24723 10016 24768 10044
rect 2317 10007 2375 10013
rect 24762 10004 24768 10016
rect 24820 10004 24826 10056
rect 26412 10047 26470 10053
rect 26412 10013 26424 10047
rect 26458 10044 26470 10047
rect 27890 10044 27896 10056
rect 26458 10016 27896 10044
rect 26458 10013 26470 10016
rect 26412 10007 26470 10013
rect 27890 10004 27896 10016
rect 27948 10004 27954 10056
rect 28000 10053 28028 10084
rect 28077 10081 28089 10115
rect 28123 10112 28135 10115
rect 29730 10112 29736 10124
rect 28123 10084 29736 10112
rect 28123 10081 28135 10084
rect 28077 10075 28135 10081
rect 29730 10072 29736 10084
rect 29788 10112 29794 10124
rect 31036 10121 31064 10152
rect 31849 10149 31861 10152
rect 31895 10180 31907 10183
rect 32030 10180 32036 10192
rect 31895 10152 32036 10180
rect 31895 10149 31907 10152
rect 31849 10143 31907 10149
rect 32030 10140 32036 10152
rect 32088 10140 32094 10192
rect 32858 10140 32864 10192
rect 32916 10180 32922 10192
rect 34054 10180 34060 10192
rect 32916 10152 33456 10180
rect 34015 10152 34060 10180
rect 32916 10140 32922 10152
rect 31021 10115 31079 10121
rect 29788 10084 30788 10112
rect 29788 10072 29794 10084
rect 27985 10047 28043 10053
rect 27985 10013 27997 10047
rect 28031 10013 28043 10047
rect 28166 10044 28172 10056
rect 28127 10016 28172 10044
rect 27985 10007 28043 10013
rect 28166 10004 28172 10016
rect 28224 10004 28230 10056
rect 29932 10053 29960 10084
rect 29917 10047 29975 10053
rect 29917 10013 29929 10047
rect 29963 10013 29975 10047
rect 30190 10044 30196 10056
rect 30151 10016 30196 10044
rect 29917 10007 29975 10013
rect 30190 10004 30196 10016
rect 30248 10004 30254 10056
rect 30760 10053 30788 10084
rect 31021 10081 31033 10115
rect 31067 10081 31079 10115
rect 31021 10075 31079 10081
rect 31481 10115 31539 10121
rect 31481 10081 31493 10115
rect 31527 10112 31539 10115
rect 33045 10115 33103 10121
rect 33045 10112 33057 10115
rect 31527 10084 33057 10112
rect 31527 10081 31539 10084
rect 31481 10075 31539 10081
rect 33045 10081 33057 10084
rect 33091 10081 33103 10115
rect 33428 10112 33456 10152
rect 34054 10140 34060 10152
rect 34112 10140 34118 10192
rect 41598 10180 41604 10192
rect 41559 10152 41604 10180
rect 41598 10140 41604 10152
rect 41656 10140 41662 10192
rect 44361 10183 44419 10189
rect 44361 10180 44373 10183
rect 43456 10152 44373 10180
rect 34885 10115 34943 10121
rect 34885 10112 34897 10115
rect 33428 10084 34897 10112
rect 33045 10075 33103 10081
rect 34885 10081 34897 10084
rect 34931 10081 34943 10115
rect 34885 10075 34943 10081
rect 36906 10072 36912 10124
rect 36964 10112 36970 10124
rect 42610 10112 42616 10124
rect 36964 10084 38332 10112
rect 36964 10072 36970 10084
rect 30745 10047 30803 10053
rect 30745 10013 30757 10047
rect 30791 10044 30803 10047
rect 31665 10047 31723 10053
rect 31665 10044 31677 10047
rect 30791 10016 31677 10044
rect 30791 10013 30803 10016
rect 30745 10007 30803 10013
rect 31665 10013 31677 10016
rect 31711 10013 31723 10047
rect 31665 10007 31723 10013
rect 31757 10047 31815 10053
rect 31757 10013 31769 10047
rect 31803 10013 31815 10047
rect 31938 10044 31944 10056
rect 31899 10016 31944 10044
rect 31757 10007 31815 10013
rect 22088 9979 22146 9985
rect 22088 9945 22100 9979
rect 22134 9976 22146 9979
rect 22370 9976 22376 9988
rect 22134 9948 22376 9976
rect 22134 9945 22146 9948
rect 22088 9939 22146 9945
rect 22370 9936 22376 9948
rect 22428 9936 22434 9988
rect 28718 9936 28724 9988
rect 28776 9976 28782 9988
rect 28813 9979 28871 9985
rect 28813 9976 28825 9979
rect 28776 9948 28825 9976
rect 28776 9936 28782 9948
rect 28813 9945 28825 9948
rect 28859 9945 28871 9979
rect 28813 9939 28871 9945
rect 29029 9979 29087 9985
rect 29029 9945 29041 9979
rect 29075 9976 29087 9979
rect 29178 9976 29184 9988
rect 29075 9948 29184 9976
rect 29075 9945 29087 9948
rect 29029 9939 29087 9945
rect 23198 9908 23204 9920
rect 23159 9880 23204 9908
rect 23198 9868 23204 9880
rect 23256 9868 23262 9920
rect 28828 9908 28856 9939
rect 29178 9936 29184 9948
rect 29236 9936 29242 9988
rect 30101 9979 30159 9985
rect 30101 9945 30113 9979
rect 30147 9945 30159 9979
rect 30101 9939 30159 9945
rect 30116 9908 30144 9939
rect 30834 9936 30840 9988
rect 30892 9976 30898 9988
rect 31386 9976 31392 9988
rect 30892 9948 31392 9976
rect 30892 9936 30898 9948
rect 31386 9936 31392 9948
rect 31444 9976 31450 9988
rect 31772 9976 31800 10007
rect 31938 10004 31944 10016
rect 31996 10004 32002 10056
rect 32953 10047 33011 10053
rect 32953 10013 32965 10047
rect 32999 10013 33011 10047
rect 32953 10007 33011 10013
rect 31444 9948 31800 9976
rect 31444 9936 31450 9948
rect 28828 9880 30144 9908
rect 32398 9868 32404 9920
rect 32456 9908 32462 9920
rect 32968 9908 32996 10007
rect 33134 10004 33140 10056
rect 33192 10044 33198 10056
rect 33781 10047 33839 10053
rect 33781 10044 33793 10047
rect 33192 10016 33793 10044
rect 33192 10004 33198 10016
rect 33781 10013 33793 10016
rect 33827 10013 33839 10047
rect 33781 10007 33839 10013
rect 35152 10047 35210 10053
rect 35152 10013 35164 10047
rect 35198 10044 35210 10047
rect 35894 10044 35900 10056
rect 35198 10016 35900 10044
rect 35198 10013 35210 10016
rect 35152 10007 35210 10013
rect 35894 10004 35900 10016
rect 35952 10004 35958 10056
rect 38194 10044 38200 10056
rect 38155 10016 38200 10044
rect 38194 10004 38200 10016
rect 38252 10004 38258 10056
rect 38304 10053 38332 10084
rect 38396 10084 39804 10112
rect 38396 10053 38424 10084
rect 38562 10054 38568 10056
rect 38289 10047 38347 10053
rect 38289 10013 38301 10047
rect 38335 10013 38347 10047
rect 38289 10007 38347 10013
rect 38381 10047 38439 10053
rect 38381 10013 38393 10047
rect 38427 10013 38439 10047
rect 38514 10047 38568 10054
rect 38514 10016 38531 10047
rect 38381 10007 38439 10013
rect 38519 10013 38531 10016
rect 38565 10013 38568 10047
rect 38519 10007 38568 10013
rect 38562 10004 38568 10007
rect 38620 10004 38626 10056
rect 38657 10047 38715 10053
rect 38657 10013 38669 10047
rect 38703 10013 38715 10047
rect 38657 10007 38715 10013
rect 38672 9976 38700 10007
rect 38746 10004 38752 10056
rect 38804 10044 38810 10056
rect 39301 10047 39359 10053
rect 39301 10044 39313 10047
rect 38804 10016 39313 10044
rect 38804 10004 38810 10016
rect 39301 10013 39313 10016
rect 39347 10013 39359 10047
rect 39301 10007 39359 10013
rect 39117 9979 39175 9985
rect 39117 9976 39129 9979
rect 38672 9948 39129 9976
rect 39117 9945 39129 9948
rect 39163 9976 39175 9979
rect 39206 9976 39212 9988
rect 39163 9948 39212 9976
rect 39163 9945 39175 9948
rect 39117 9939 39175 9945
rect 39206 9936 39212 9948
rect 39264 9936 39270 9988
rect 34241 9911 34299 9917
rect 34241 9908 34253 9911
rect 32456 9880 34253 9908
rect 32456 9868 32462 9880
rect 34241 9877 34253 9880
rect 34287 9877 34299 9911
rect 38010 9908 38016 9920
rect 37971 9880 38016 9908
rect 34241 9871 34299 9877
rect 38010 9868 38016 9880
rect 38068 9868 38074 9920
rect 39390 9868 39396 9920
rect 39448 9908 39454 9920
rect 39485 9911 39543 9917
rect 39485 9908 39497 9911
rect 39448 9880 39497 9908
rect 39448 9868 39454 9880
rect 39485 9877 39497 9880
rect 39531 9877 39543 9911
rect 39776 9908 39804 10084
rect 41386 10084 42616 10112
rect 40218 10044 40224 10056
rect 40179 10016 40224 10044
rect 40218 10004 40224 10016
rect 40276 10044 40282 10056
rect 41386 10044 41414 10084
rect 42610 10072 42616 10084
rect 42668 10072 42674 10124
rect 43456 10121 43484 10152
rect 44361 10149 44373 10152
rect 44407 10149 44419 10183
rect 44361 10143 44419 10149
rect 43441 10115 43499 10121
rect 43441 10081 43453 10115
rect 43487 10081 43499 10115
rect 43898 10112 43904 10124
rect 43859 10084 43904 10112
rect 43441 10075 43499 10081
rect 43898 10072 43904 10084
rect 43956 10072 43962 10124
rect 44174 10072 44180 10124
rect 44232 10112 44238 10124
rect 44232 10084 44680 10112
rect 44232 10072 44238 10084
rect 42058 10044 42064 10056
rect 40276 10016 41414 10044
rect 42019 10016 42064 10044
rect 40276 10004 40282 10016
rect 42058 10004 42064 10016
rect 42116 10004 42122 10056
rect 43530 10004 43536 10056
rect 43588 10044 43594 10056
rect 43806 10044 43812 10056
rect 43588 10016 43633 10044
rect 43767 10016 43812 10044
rect 43588 10004 43594 10016
rect 43806 10004 43812 10016
rect 43864 10004 43870 10056
rect 44082 10004 44088 10056
rect 44140 10044 44146 10056
rect 44652 10053 44680 10084
rect 44361 10047 44419 10053
rect 44361 10044 44373 10047
rect 44140 10016 44373 10044
rect 44140 10004 44146 10016
rect 44361 10013 44373 10016
rect 44407 10013 44419 10047
rect 44361 10007 44419 10013
rect 44637 10047 44695 10053
rect 44637 10013 44649 10047
rect 44683 10013 44695 10047
rect 44637 10007 44695 10013
rect 44910 10004 44916 10056
rect 44968 10044 44974 10056
rect 45189 10047 45247 10053
rect 45189 10044 45201 10047
rect 44968 10016 45201 10044
rect 44968 10004 44974 10016
rect 45189 10013 45201 10016
rect 45235 10013 45247 10047
rect 45189 10007 45247 10013
rect 40310 9936 40316 9988
rect 40368 9976 40374 9988
rect 40466 9979 40524 9985
rect 40466 9976 40478 9979
rect 40368 9948 40478 9976
rect 40368 9936 40374 9948
rect 40466 9945 40478 9948
rect 40512 9945 40524 9979
rect 45370 9976 45376 9988
rect 45331 9948 45376 9976
rect 40466 9939 40524 9945
rect 45370 9936 45376 9948
rect 45428 9936 45434 9988
rect 40586 9908 40592 9920
rect 39776 9880 40592 9908
rect 39485 9871 39543 9877
rect 40586 9868 40592 9880
rect 40644 9868 40650 9920
rect 43254 9908 43260 9920
rect 43215 9880 43260 9908
rect 43254 9868 43260 9880
rect 43312 9868 43318 9920
rect 44545 9911 44603 9917
rect 44545 9877 44557 9911
rect 44591 9908 44603 9911
rect 44818 9908 44824 9920
rect 44591 9880 44824 9908
rect 44591 9877 44603 9880
rect 44545 9871 44603 9877
rect 44818 9868 44824 9880
rect 44876 9868 44882 9920
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 22370 9704 22376 9716
rect 22331 9676 22376 9704
rect 22370 9664 22376 9676
rect 22428 9664 22434 9716
rect 23198 9664 23204 9716
rect 23256 9704 23262 9716
rect 28166 9704 28172 9716
rect 23256 9676 28172 9704
rect 23256 9664 23262 9676
rect 2038 9568 2044 9580
rect 1999 9540 2044 9568
rect 2038 9528 2044 9540
rect 2096 9528 2102 9580
rect 22554 9568 22560 9580
rect 22515 9540 22560 9568
rect 22554 9528 22560 9540
rect 22612 9528 22618 9580
rect 22738 9568 22744 9580
rect 22699 9540 22744 9568
rect 22738 9528 22744 9540
rect 22796 9528 22802 9580
rect 22833 9571 22891 9577
rect 22833 9537 22845 9571
rect 22879 9568 22891 9571
rect 23198 9568 23204 9580
rect 22879 9540 23204 9568
rect 22879 9537 22891 9540
rect 22833 9531 22891 9537
rect 23198 9528 23204 9540
rect 23256 9528 23262 9580
rect 27706 9528 27712 9580
rect 27764 9568 27770 9580
rect 28092 9577 28120 9676
rect 28166 9664 28172 9676
rect 28224 9664 28230 9716
rect 29822 9664 29828 9716
rect 29880 9704 29886 9716
rect 30009 9707 30067 9713
rect 30009 9704 30021 9707
rect 29880 9676 30021 9704
rect 29880 9664 29886 9676
rect 30009 9673 30021 9676
rect 30055 9673 30067 9707
rect 30009 9667 30067 9673
rect 32766 9664 32772 9716
rect 32824 9704 32830 9716
rect 32861 9707 32919 9713
rect 32861 9704 32873 9707
rect 32824 9676 32873 9704
rect 32824 9664 32830 9676
rect 32861 9673 32873 9676
rect 32907 9673 32919 9707
rect 32861 9667 32919 9673
rect 35710 9664 35716 9716
rect 35768 9704 35774 9716
rect 38562 9704 38568 9716
rect 35768 9676 38568 9704
rect 35768 9664 35774 9676
rect 38562 9664 38568 9676
rect 38620 9704 38626 9716
rect 40678 9704 40684 9716
rect 38620 9676 40684 9704
rect 38620 9664 38626 9676
rect 40678 9664 40684 9676
rect 40736 9704 40742 9716
rect 43806 9704 43812 9716
rect 40736 9676 41736 9704
rect 40736 9664 40742 9676
rect 29086 9636 29092 9648
rect 28644 9608 29092 9636
rect 27893 9571 27951 9577
rect 27893 9568 27905 9571
rect 27764 9540 27905 9568
rect 27764 9528 27770 9540
rect 27893 9537 27905 9540
rect 27939 9537 27951 9571
rect 27893 9531 27951 9537
rect 28077 9571 28135 9577
rect 28077 9537 28089 9571
rect 28123 9537 28135 9571
rect 28077 9531 28135 9537
rect 2225 9503 2283 9509
rect 2225 9469 2237 9503
rect 2271 9500 2283 9503
rect 2314 9500 2320 9512
rect 2271 9472 2320 9500
rect 2271 9469 2283 9472
rect 2225 9463 2283 9469
rect 2314 9460 2320 9472
rect 2372 9460 2378 9512
rect 2774 9500 2780 9512
rect 2735 9472 2780 9500
rect 2774 9460 2780 9472
rect 2832 9460 2838 9512
rect 27985 9503 28043 9509
rect 27985 9469 27997 9503
rect 28031 9500 28043 9503
rect 28644 9500 28672 9608
rect 29086 9596 29092 9608
rect 29144 9636 29150 9648
rect 30190 9636 30196 9648
rect 29144 9608 30196 9636
rect 29144 9596 29150 9608
rect 28721 9571 28779 9577
rect 28721 9537 28733 9571
rect 28767 9568 28779 9571
rect 28994 9568 29000 9580
rect 28767 9540 29000 9568
rect 28767 9537 28779 9540
rect 28721 9531 28779 9537
rect 28994 9528 29000 9540
rect 29052 9528 29058 9580
rect 29564 9577 29592 9608
rect 30190 9596 30196 9608
rect 30248 9596 30254 9648
rect 40218 9636 40224 9648
rect 37476 9608 40224 9636
rect 29549 9571 29607 9577
rect 29549 9537 29561 9571
rect 29595 9537 29607 9571
rect 29549 9531 29607 9537
rect 31389 9571 31447 9577
rect 31389 9537 31401 9571
rect 31435 9568 31447 9571
rect 32030 9568 32036 9580
rect 31435 9540 32036 9568
rect 31435 9537 31447 9540
rect 31389 9531 31447 9537
rect 32030 9528 32036 9540
rect 32088 9528 32094 9580
rect 32398 9568 32404 9580
rect 32359 9540 32404 9568
rect 32398 9528 32404 9540
rect 32456 9528 32462 9580
rect 37476 9577 37504 9608
rect 40218 9596 40224 9608
rect 40276 9596 40282 9648
rect 40497 9639 40555 9645
rect 40497 9605 40509 9639
rect 40543 9636 40555 9639
rect 41138 9636 41144 9648
rect 40543 9608 41144 9636
rect 40543 9605 40555 9608
rect 40497 9599 40555 9605
rect 41138 9596 41144 9608
rect 41196 9596 41202 9648
rect 41598 9636 41604 9648
rect 41386 9608 41604 9636
rect 35621 9571 35679 9577
rect 35621 9537 35633 9571
rect 35667 9568 35679 9571
rect 37461 9571 37519 9577
rect 35667 9540 37412 9568
rect 35667 9537 35679 9540
rect 35621 9531 35679 9537
rect 28031 9472 28672 9500
rect 28813 9503 28871 9509
rect 28031 9469 28043 9472
rect 27985 9463 28043 9469
rect 28813 9469 28825 9503
rect 28859 9500 28871 9503
rect 29822 9500 29828 9512
rect 28859 9472 29828 9500
rect 28859 9469 28871 9472
rect 28813 9463 28871 9469
rect 29822 9460 29828 9472
rect 29880 9460 29886 9512
rect 31481 9503 31539 9509
rect 31481 9469 31493 9503
rect 31527 9469 31539 9503
rect 31481 9463 31539 9469
rect 35713 9503 35771 9509
rect 35713 9469 35725 9503
rect 35759 9469 35771 9503
rect 35986 9500 35992 9512
rect 35947 9472 35992 9500
rect 35713 9463 35771 9469
rect 31496 9432 31524 9463
rect 29748 9404 31524 9432
rect 31757 9435 31815 9441
rect 29748 9376 29776 9404
rect 31757 9401 31769 9435
rect 31803 9432 31815 9435
rect 31846 9432 31852 9444
rect 31803 9404 31852 9432
rect 31803 9401 31815 9404
rect 31757 9395 31815 9401
rect 31846 9392 31852 9404
rect 31904 9392 31910 9444
rect 35618 9392 35624 9444
rect 35676 9432 35682 9444
rect 35728 9432 35756 9463
rect 35986 9460 35992 9472
rect 36044 9460 36050 9512
rect 35676 9404 35756 9432
rect 35676 9392 35682 9404
rect 28902 9324 28908 9376
rect 28960 9364 28966 9376
rect 28997 9367 29055 9373
rect 28997 9364 29009 9367
rect 28960 9336 29009 9364
rect 28960 9324 28966 9336
rect 28997 9333 29009 9336
rect 29043 9333 29055 9367
rect 29730 9364 29736 9376
rect 29691 9336 29736 9364
rect 28997 9327 29055 9333
rect 29730 9324 29736 9336
rect 29788 9324 29794 9376
rect 31386 9364 31392 9376
rect 31347 9336 31392 9364
rect 31386 9324 31392 9336
rect 31444 9324 31450 9376
rect 32030 9324 32036 9376
rect 32088 9364 32094 9376
rect 32493 9367 32551 9373
rect 32493 9364 32505 9367
rect 32088 9336 32505 9364
rect 32088 9324 32094 9336
rect 32493 9333 32505 9336
rect 32539 9333 32551 9367
rect 37384 9364 37412 9540
rect 37461 9537 37473 9571
rect 37507 9537 37519 9571
rect 37461 9531 37519 9537
rect 37728 9571 37786 9577
rect 37728 9537 37740 9571
rect 37774 9568 37786 9571
rect 38010 9568 38016 9580
rect 37774 9540 38016 9568
rect 37774 9537 37786 9540
rect 37728 9531 37786 9537
rect 38010 9528 38016 9540
rect 38068 9528 38074 9580
rect 39301 9571 39359 9577
rect 39301 9537 39313 9571
rect 39347 9568 39359 9571
rect 39390 9568 39396 9580
rect 39347 9540 39396 9568
rect 39347 9537 39359 9540
rect 39301 9531 39359 9537
rect 39390 9528 39396 9540
rect 39448 9528 39454 9580
rect 39482 9528 39488 9580
rect 39540 9568 39546 9580
rect 40126 9568 40132 9580
rect 39540 9540 40132 9568
rect 39540 9528 39546 9540
rect 40126 9528 40132 9540
rect 40184 9528 40190 9580
rect 40402 9568 40408 9580
rect 40363 9540 40408 9568
rect 40402 9528 40408 9540
rect 40460 9528 40466 9580
rect 40586 9568 40592 9580
rect 40547 9540 40592 9568
rect 40586 9528 40592 9540
rect 40644 9528 40650 9580
rect 40678 9528 40684 9580
rect 40736 9577 40742 9580
rect 40736 9571 40765 9577
rect 40753 9537 40765 9571
rect 40736 9531 40765 9537
rect 40865 9571 40923 9577
rect 40865 9537 40877 9571
rect 40911 9568 40923 9571
rect 41386 9568 41414 9608
rect 41598 9596 41604 9608
rect 41656 9596 41662 9648
rect 41708 9636 41736 9676
rect 42812 9676 43812 9704
rect 42812 9636 42840 9676
rect 43806 9664 43812 9676
rect 43864 9664 43870 9716
rect 43898 9664 43904 9716
rect 43956 9704 43962 9716
rect 43993 9707 44051 9713
rect 43993 9704 44005 9707
rect 43956 9676 44005 9704
rect 43956 9664 43962 9676
rect 43993 9673 44005 9676
rect 44039 9673 44051 9707
rect 43993 9667 44051 9673
rect 41708 9608 42840 9636
rect 42880 9639 42938 9645
rect 42880 9605 42892 9639
rect 42926 9636 42938 9639
rect 43254 9636 43260 9648
rect 42926 9608 43260 9636
rect 42926 9605 42938 9608
rect 42880 9599 42938 9605
rect 43254 9596 43260 9608
rect 43312 9596 43318 9648
rect 44821 9639 44879 9645
rect 44821 9605 44833 9639
rect 44867 9636 44879 9639
rect 45646 9636 45652 9648
rect 44867 9608 45652 9636
rect 44867 9605 44879 9608
rect 44821 9599 44879 9605
rect 45646 9596 45652 9608
rect 45704 9596 45710 9648
rect 41509 9571 41567 9577
rect 40911 9540 41460 9568
rect 40911 9537 40923 9540
rect 40865 9531 40923 9537
rect 40736 9528 40742 9531
rect 40221 9503 40279 9509
rect 40221 9469 40233 9503
rect 40267 9500 40279 9503
rect 40310 9500 40316 9512
rect 40267 9472 40316 9500
rect 40267 9469 40279 9472
rect 40221 9463 40279 9469
rect 40310 9460 40316 9472
rect 40368 9460 40374 9512
rect 41432 9509 41460 9540
rect 41509 9537 41521 9571
rect 41555 9537 41567 9571
rect 42610 9568 42616 9580
rect 42571 9540 42616 9568
rect 41509 9531 41567 9537
rect 41417 9503 41475 9509
rect 41417 9469 41429 9503
rect 41463 9469 41475 9503
rect 41417 9463 41475 9469
rect 38470 9392 38476 9444
rect 38528 9432 38534 9444
rect 39393 9435 39451 9441
rect 39393 9432 39405 9435
rect 38528 9404 39405 9432
rect 38528 9392 38534 9404
rect 39393 9401 39405 9404
rect 39439 9401 39451 9435
rect 39393 9395 39451 9401
rect 41322 9392 41328 9444
rect 41380 9432 41386 9444
rect 41524 9432 41552 9531
rect 42610 9528 42616 9540
rect 42668 9528 42674 9580
rect 44082 9528 44088 9580
rect 44140 9568 44146 9580
rect 44453 9571 44511 9577
rect 44453 9568 44465 9571
rect 44140 9540 44465 9568
rect 44140 9528 44146 9540
rect 44453 9537 44465 9540
rect 44499 9537 44511 9571
rect 44453 9531 44511 9537
rect 41877 9503 41935 9509
rect 41877 9469 41889 9503
rect 41923 9500 41935 9503
rect 42058 9500 42064 9512
rect 41923 9472 42064 9500
rect 41923 9469 41935 9472
rect 41877 9463 41935 9469
rect 42058 9460 42064 9472
rect 42116 9460 42122 9512
rect 45002 9432 45008 9444
rect 41380 9404 41552 9432
rect 44963 9404 45008 9432
rect 41380 9392 41386 9404
rect 45002 9392 45008 9404
rect 45060 9392 45066 9444
rect 38746 9364 38752 9376
rect 37384 9336 38752 9364
rect 32493 9327 32551 9333
rect 38746 9324 38752 9336
rect 38804 9324 38810 9376
rect 38841 9367 38899 9373
rect 38841 9333 38853 9367
rect 38887 9364 38899 9367
rect 39206 9364 39212 9376
rect 38887 9336 39212 9364
rect 38887 9333 38899 9336
rect 38841 9327 38899 9333
rect 39206 9324 39212 9336
rect 39264 9324 39270 9376
rect 44818 9364 44824 9376
rect 44779 9336 44824 9364
rect 44818 9324 44824 9336
rect 44876 9324 44882 9376
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 2314 9160 2320 9172
rect 2275 9132 2320 9160
rect 2314 9120 2320 9132
rect 2372 9120 2378 9172
rect 32030 9160 32036 9172
rect 31991 9132 32036 9160
rect 32030 9120 32036 9132
rect 32088 9120 32094 9172
rect 39301 9163 39359 9169
rect 39301 9129 39313 9163
rect 39347 9160 39359 9163
rect 39482 9160 39488 9172
rect 39347 9132 39488 9160
rect 39347 9129 39359 9132
rect 39301 9123 39359 9129
rect 39482 9120 39488 9132
rect 39540 9120 39546 9172
rect 39666 9120 39672 9172
rect 39724 9160 39730 9172
rect 48041 9163 48099 9169
rect 48041 9160 48053 9163
rect 39724 9132 48053 9160
rect 39724 9120 39730 9132
rect 48041 9129 48053 9132
rect 48087 9129 48099 9163
rect 48041 9123 48099 9129
rect 44082 9092 44088 9104
rect 44043 9064 44088 9092
rect 44082 9052 44088 9064
rect 44140 9052 44146 9104
rect 38746 8984 38752 9036
rect 38804 9024 38810 9036
rect 43809 9027 43867 9033
rect 38804 8996 39436 9024
rect 38804 8984 38810 8996
rect 2222 8956 2228 8968
rect 2183 8928 2228 8956
rect 2222 8916 2228 8928
rect 2280 8956 2286 8968
rect 8294 8956 8300 8968
rect 2280 8928 8300 8956
rect 2280 8916 2286 8928
rect 8294 8916 8300 8928
rect 8352 8916 8358 8968
rect 31938 8956 31944 8968
rect 31899 8928 31944 8956
rect 31938 8916 31944 8928
rect 31996 8916 32002 8968
rect 32122 8956 32128 8968
rect 32083 8928 32128 8956
rect 32122 8916 32128 8928
rect 32180 8916 32186 8968
rect 39206 8956 39212 8968
rect 39167 8928 39212 8956
rect 39206 8916 39212 8928
rect 39264 8916 39270 8968
rect 39408 8965 39436 8996
rect 43809 8993 43821 9027
rect 43855 9024 43867 9027
rect 43898 9024 43904 9036
rect 43855 8996 43904 9024
rect 43855 8993 43867 8996
rect 43809 8987 43867 8993
rect 43898 8984 43904 8996
rect 43956 8984 43962 9036
rect 39393 8959 39451 8965
rect 39393 8925 39405 8959
rect 39439 8956 39451 8959
rect 41322 8956 41328 8968
rect 39439 8928 41328 8956
rect 39439 8925 39451 8928
rect 39393 8919 39451 8925
rect 41322 8916 41328 8928
rect 41380 8956 41386 8968
rect 43717 8959 43775 8965
rect 43717 8956 43729 8959
rect 41380 8928 43729 8956
rect 41380 8916 41386 8928
rect 43717 8925 43729 8928
rect 43763 8956 43775 8959
rect 45370 8956 45376 8968
rect 43763 8928 45376 8956
rect 43763 8925 43775 8928
rect 43717 8919 43775 8925
rect 45370 8916 45376 8928
rect 45428 8916 45434 8968
rect 47946 8888 47952 8900
rect 47907 8860 47952 8888
rect 47946 8848 47952 8860
rect 48004 8848 48010 8900
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 47854 8480 47860 8492
rect 47815 8452 47860 8480
rect 47854 8440 47860 8452
rect 47912 8440 47918 8492
rect 32214 8372 32220 8424
rect 32272 8412 32278 8424
rect 48041 8415 48099 8421
rect 48041 8412 48053 8415
rect 32272 8384 48053 8412
rect 32272 8372 32278 8384
rect 48041 8381 48053 8384
rect 48087 8381 48099 8415
rect 48041 8375 48099 8381
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 2038 7828 2044 7880
rect 2096 7868 2102 7880
rect 2317 7871 2375 7877
rect 2317 7868 2329 7871
rect 2096 7840 2329 7868
rect 2096 7828 2102 7840
rect 2317 7837 2329 7840
rect 2363 7837 2375 7871
rect 2317 7831 2375 7837
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7868 2835 7871
rect 3234 7868 3240 7880
rect 2823 7840 3240 7868
rect 2823 7837 2835 7840
rect 2777 7831 2835 7837
rect 3234 7828 3240 7840
rect 3292 7868 3298 7880
rect 5626 7868 5632 7880
rect 3292 7840 5632 7868
rect 3292 7828 3298 7840
rect 5626 7828 5632 7840
rect 5684 7828 5690 7880
rect 2222 7692 2228 7744
rect 2280 7732 2286 7744
rect 2869 7735 2927 7741
rect 2869 7732 2881 7735
rect 2280 7704 2881 7732
rect 2280 7692 2286 7704
rect 2869 7701 2881 7704
rect 2915 7701 2927 7735
rect 2869 7695 2927 7701
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 2222 7460 2228 7472
rect 2183 7432 2228 7460
rect 2222 7420 2228 7432
rect 2280 7420 2286 7472
rect 2038 7392 2044 7404
rect 1999 7364 2044 7392
rect 2038 7352 2044 7364
rect 2096 7352 2102 7404
rect 2774 7324 2780 7336
rect 2735 7296 2780 7324
rect 2774 7284 2780 7296
rect 2832 7284 2838 7336
rect 47946 7188 47952 7200
rect 47907 7160 47952 7188
rect 47946 7148 47952 7160
rect 48004 7148 48010 7200
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 2774 6848 2780 6860
rect 2735 6820 2780 6848
rect 2774 6808 2780 6820
rect 2832 6808 2838 6860
rect 46477 6851 46535 6857
rect 46477 6817 46489 6851
rect 46523 6848 46535 6851
rect 47946 6848 47952 6860
rect 46523 6820 47952 6848
rect 46523 6817 46535 6820
rect 46477 6811 46535 6817
rect 47946 6808 47952 6820
rect 48004 6808 48010 6860
rect 48222 6848 48228 6860
rect 48183 6820 48228 6848
rect 48222 6808 48228 6820
rect 48280 6808 48286 6860
rect 1578 6780 1584 6792
rect 1539 6752 1584 6780
rect 1578 6740 1584 6752
rect 1636 6740 1642 6792
rect 1762 6712 1768 6724
rect 1723 6684 1768 6712
rect 1762 6672 1768 6684
rect 1820 6672 1826 6724
rect 46661 6715 46719 6721
rect 46661 6681 46673 6715
rect 46707 6712 46719 6715
rect 47854 6712 47860 6724
rect 46707 6684 47860 6712
rect 46707 6681 46719 6684
rect 46661 6675 46719 6681
rect 47854 6672 47860 6684
rect 47912 6672 47918 6724
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 1762 6400 1768 6452
rect 1820 6440 1826 6452
rect 2869 6443 2927 6449
rect 2869 6440 2881 6443
rect 1820 6412 2881 6440
rect 1820 6400 1826 6412
rect 2869 6409 2881 6412
rect 2915 6409 2927 6443
rect 47854 6440 47860 6452
rect 47815 6412 47860 6440
rect 2869 6403 2927 6409
rect 47854 6400 47860 6412
rect 47912 6400 47918 6452
rect 41386 6344 47808 6372
rect 1578 6264 1584 6316
rect 1636 6304 1642 6316
rect 2317 6307 2375 6313
rect 2317 6304 2329 6307
rect 1636 6276 2329 6304
rect 1636 6264 1642 6276
rect 2317 6273 2329 6276
rect 2363 6273 2375 6307
rect 2317 6267 2375 6273
rect 2777 6307 2835 6313
rect 2777 6273 2789 6307
rect 2823 6304 2835 6307
rect 2866 6304 2872 6316
rect 2823 6276 2872 6304
rect 2823 6273 2835 6276
rect 2777 6267 2835 6273
rect 2866 6264 2872 6276
rect 2924 6304 2930 6316
rect 39025 6307 39083 6313
rect 39025 6304 39037 6307
rect 2924 6276 39037 6304
rect 2924 6264 2930 6276
rect 39025 6273 39037 6276
rect 39071 6304 39083 6307
rect 41386 6304 41414 6344
rect 47780 6316 47808 6344
rect 39071 6276 41414 6304
rect 46385 6307 46443 6313
rect 39071 6273 39083 6276
rect 39025 6267 39083 6273
rect 46385 6273 46397 6307
rect 46431 6304 46443 6307
rect 47026 6304 47032 6316
rect 46431 6276 47032 6304
rect 46431 6273 46443 6276
rect 46385 6267 46443 6273
rect 47026 6264 47032 6276
rect 47084 6264 47090 6316
rect 47762 6304 47768 6316
rect 47675 6276 47768 6304
rect 47762 6264 47768 6276
rect 47820 6264 47826 6316
rect 39117 6103 39175 6109
rect 39117 6069 39129 6103
rect 39163 6100 39175 6103
rect 39206 6100 39212 6112
rect 39163 6072 39212 6100
rect 39163 6069 39175 6072
rect 39117 6063 39175 6069
rect 39206 6060 39212 6072
rect 39264 6060 39270 6112
rect 43070 6060 43076 6112
rect 43128 6100 43134 6112
rect 45925 6103 45983 6109
rect 45925 6100 45937 6103
rect 43128 6072 45937 6100
rect 43128 6060 43134 6072
rect 45925 6069 45937 6072
rect 45971 6069 45983 6103
rect 46474 6100 46480 6112
rect 46435 6072 46480 6100
rect 45925 6063 45983 6069
rect 46474 6060 46480 6072
rect 46532 6060 46538 6112
rect 47210 6100 47216 6112
rect 47171 6072 47216 6100
rect 47210 6060 47216 6072
rect 47268 6060 47274 6112
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 46477 5763 46535 5769
rect 46477 5729 46489 5763
rect 46523 5760 46535 5763
rect 47210 5760 47216 5772
rect 46523 5732 47216 5760
rect 46523 5729 46535 5732
rect 46477 5723 46535 5729
rect 47210 5720 47216 5732
rect 47268 5720 47274 5772
rect 48222 5760 48228 5772
rect 48183 5732 48228 5760
rect 48222 5720 48228 5732
rect 48280 5720 48286 5772
rect 1854 5692 1860 5704
rect 1815 5664 1860 5692
rect 1854 5652 1860 5664
rect 1912 5652 1918 5704
rect 2317 5695 2375 5701
rect 2317 5661 2329 5695
rect 2363 5692 2375 5695
rect 2682 5692 2688 5704
rect 2363 5664 2688 5692
rect 2363 5661 2375 5664
rect 2317 5655 2375 5661
rect 2682 5652 2688 5664
rect 2740 5652 2746 5704
rect 3142 5692 3148 5704
rect 3103 5664 3148 5692
rect 3142 5652 3148 5664
rect 3200 5652 3206 5704
rect 9766 5692 9772 5704
rect 9727 5664 9772 5692
rect 9766 5652 9772 5664
rect 9824 5652 9830 5704
rect 10229 5695 10287 5701
rect 10229 5661 10241 5695
rect 10275 5692 10287 5695
rect 16114 5692 16120 5704
rect 10275 5664 16120 5692
rect 10275 5661 10287 5664
rect 10229 5655 10287 5661
rect 16114 5652 16120 5664
rect 16172 5652 16178 5704
rect 39022 5652 39028 5704
rect 39080 5692 39086 5704
rect 39209 5695 39267 5701
rect 39209 5692 39221 5695
rect 39080 5664 39221 5692
rect 39080 5652 39086 5664
rect 39209 5661 39221 5664
rect 39255 5661 39267 5695
rect 46014 5692 46020 5704
rect 45975 5664 46020 5692
rect 39209 5655 39267 5661
rect 46014 5652 46020 5664
rect 46072 5652 46078 5704
rect 46661 5627 46719 5633
rect 46661 5593 46673 5627
rect 46707 5624 46719 5627
rect 47578 5624 47584 5636
rect 46707 5596 47584 5624
rect 46707 5593 46719 5596
rect 46661 5587 46719 5593
rect 47578 5584 47584 5596
rect 47636 5584 47642 5636
rect 1762 5516 1768 5568
rect 1820 5556 1826 5568
rect 2409 5559 2467 5565
rect 2409 5556 2421 5559
rect 1820 5528 2421 5556
rect 1820 5516 1826 5528
rect 2409 5525 2421 5528
rect 2455 5525 2467 5559
rect 2409 5519 2467 5525
rect 10042 5516 10048 5568
rect 10100 5556 10106 5568
rect 10321 5559 10379 5565
rect 10321 5556 10333 5559
rect 10100 5528 10333 5556
rect 10100 5516 10106 5528
rect 10321 5525 10333 5528
rect 10367 5525 10379 5559
rect 10321 5519 10379 5525
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 47486 5352 47492 5364
rect 44744 5324 47492 5352
rect 39206 5284 39212 5296
rect 39167 5256 39212 5284
rect 39206 5244 39212 5256
rect 39264 5244 39270 5296
rect 39022 5216 39028 5228
rect 38983 5188 39028 5216
rect 39022 5176 39028 5188
rect 39080 5176 39086 5228
rect 44744 5225 44772 5324
rect 47486 5312 47492 5324
rect 47544 5312 47550 5364
rect 45557 5287 45615 5293
rect 45557 5253 45569 5287
rect 45603 5284 45615 5287
rect 47857 5287 47915 5293
rect 47857 5284 47869 5287
rect 45603 5256 47869 5284
rect 45603 5253 45615 5256
rect 45557 5247 45615 5253
rect 47857 5253 47869 5256
rect 47903 5253 47915 5287
rect 47857 5247 47915 5253
rect 44729 5219 44787 5225
rect 44729 5185 44741 5219
rect 44775 5185 44787 5219
rect 47762 5216 47768 5228
rect 47723 5188 47768 5216
rect 44729 5179 44787 5185
rect 47762 5176 47768 5188
rect 47820 5176 47826 5228
rect 1765 5151 1823 5157
rect 1765 5117 1777 5151
rect 1811 5148 1823 5151
rect 2225 5151 2283 5157
rect 2225 5148 2237 5151
rect 1811 5120 2237 5148
rect 1811 5117 1823 5120
rect 1765 5111 1823 5117
rect 2225 5117 2237 5120
rect 2271 5117 2283 5151
rect 2225 5111 2283 5117
rect 2409 5151 2467 5157
rect 2409 5117 2421 5151
rect 2455 5148 2467 5151
rect 2866 5148 2872 5160
rect 2455 5120 2872 5148
rect 2455 5117 2467 5120
rect 2409 5111 2467 5117
rect 2866 5108 2872 5120
rect 2924 5108 2930 5160
rect 2958 5108 2964 5160
rect 3016 5148 3022 5160
rect 40034 5148 40040 5160
rect 3016 5120 3061 5148
rect 39995 5120 40040 5148
rect 3016 5108 3022 5120
rect 40034 5108 40040 5120
rect 40092 5108 40098 5160
rect 45373 5151 45431 5157
rect 45373 5117 45385 5151
rect 45419 5148 45431 5151
rect 46014 5148 46020 5160
rect 45419 5120 46020 5148
rect 45419 5117 45431 5120
rect 45373 5111 45431 5117
rect 46014 5108 46020 5120
rect 46072 5108 46078 5160
rect 47210 5148 47216 5160
rect 47171 5120 47216 5148
rect 47210 5108 47216 5120
rect 47268 5108 47274 5160
rect 44266 5012 44272 5024
rect 44227 4984 44272 5012
rect 44266 4972 44272 4984
rect 44324 4972 44330 5024
rect 44821 5015 44879 5021
rect 44821 4981 44833 5015
rect 44867 5012 44879 5015
rect 45370 5012 45376 5024
rect 44867 4984 45376 5012
rect 44867 4981 44879 4984
rect 44821 4975 44879 4981
rect 45370 4972 45376 4984
rect 45428 4972 45434 5024
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 47578 4808 47584 4820
rect 47539 4780 47584 4808
rect 47578 4768 47584 4780
rect 47636 4768 47642 4820
rect 3142 4740 3148 4752
rect 1596 4712 3148 4740
rect 1596 4681 1624 4712
rect 3142 4700 3148 4712
rect 3200 4700 3206 4752
rect 47670 4740 47676 4752
rect 6886 4712 10364 4740
rect 1581 4675 1639 4681
rect 1581 4641 1593 4675
rect 1627 4641 1639 4675
rect 1762 4672 1768 4684
rect 1723 4644 1768 4672
rect 1581 4635 1639 4641
rect 1762 4632 1768 4644
rect 1820 4632 1826 4684
rect 2774 4672 2780 4684
rect 2735 4644 2780 4672
rect 2774 4632 2780 4644
rect 2832 4632 2838 4684
rect 3510 4632 3516 4684
rect 3568 4672 3574 4684
rect 6886 4672 6914 4712
rect 3568 4644 6914 4672
rect 3568 4632 3574 4644
rect 9766 4632 9772 4684
rect 9824 4672 9830 4684
rect 9861 4675 9919 4681
rect 9861 4672 9873 4675
rect 9824 4644 9873 4672
rect 9824 4632 9830 4644
rect 9861 4641 9873 4644
rect 9907 4641 9919 4675
rect 10042 4672 10048 4684
rect 10003 4644 10048 4672
rect 9861 4635 9919 4641
rect 10042 4632 10048 4644
rect 10100 4632 10106 4684
rect 10336 4681 10364 4712
rect 43824 4712 47676 4740
rect 10321 4675 10379 4681
rect 10321 4641 10333 4675
rect 10367 4641 10379 4675
rect 10321 4635 10379 4641
rect 4157 4607 4215 4613
rect 4157 4573 4169 4607
rect 4203 4604 4215 4607
rect 4614 4604 4620 4616
rect 4203 4576 4620 4604
rect 4203 4573 4215 4576
rect 4157 4567 4215 4573
rect 4614 4564 4620 4576
rect 4672 4564 4678 4616
rect 4982 4604 4988 4616
rect 4943 4576 4988 4604
rect 4982 4564 4988 4576
rect 5040 4564 5046 4616
rect 5534 4604 5540 4616
rect 5495 4576 5540 4604
rect 5534 4564 5540 4576
rect 5592 4564 5598 4616
rect 43824 4613 43852 4712
rect 47670 4700 47676 4712
rect 47728 4700 47734 4752
rect 44266 4632 44272 4684
rect 44324 4672 44330 4684
rect 45189 4675 45247 4681
rect 45189 4672 45201 4675
rect 44324 4644 45201 4672
rect 44324 4632 44330 4644
rect 45189 4641 45201 4644
rect 45235 4641 45247 4675
rect 45370 4672 45376 4684
rect 45331 4644 45376 4672
rect 45189 4635 45247 4641
rect 45370 4632 45376 4644
rect 45428 4632 45434 4684
rect 45646 4672 45652 4684
rect 45607 4644 45652 4672
rect 45646 4632 45652 4644
rect 45704 4632 45710 4684
rect 43809 4607 43867 4613
rect 43809 4573 43821 4607
rect 43855 4573 43867 4607
rect 44634 4604 44640 4616
rect 44595 4576 44640 4604
rect 43809 4567 43867 4573
rect 44634 4564 44640 4576
rect 44692 4564 44698 4616
rect 47486 4604 47492 4616
rect 47447 4576 47492 4604
rect 47486 4564 47492 4576
rect 47544 4564 47550 4616
rect 48130 4604 48136 4616
rect 48091 4576 48136 4604
rect 48130 4564 48136 4576
rect 48188 4564 48194 4616
rect 6270 4536 6276 4548
rect 6231 4508 6276 4536
rect 6270 4496 6276 4508
rect 6328 4536 6334 4548
rect 6328 4508 6914 4536
rect 6328 4496 6334 4508
rect 6886 4468 6914 4508
rect 39942 4468 39948 4480
rect 6886 4440 39948 4468
rect 39942 4428 39948 4440
rect 40000 4428 40006 4480
rect 43254 4428 43260 4480
rect 43312 4468 43318 4480
rect 43901 4471 43959 4477
rect 43901 4468 43913 4471
rect 43312 4440 43913 4468
rect 43312 4428 43318 4440
rect 43901 4437 43913 4440
rect 43947 4437 43959 4471
rect 43901 4431 43959 4437
rect 46934 4428 46940 4480
rect 46992 4468 46998 4480
rect 48225 4471 48283 4477
rect 48225 4468 48237 4471
rect 46992 4440 48237 4468
rect 46992 4428 46998 4440
rect 48225 4437 48237 4440
rect 48271 4437 48283 4471
rect 48225 4431 48283 4437
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 48130 4264 48136 4276
rect 45296 4236 48136 4264
rect 43254 4196 43260 4208
rect 2792 4168 3096 4196
rect 2792 4137 2820 4168
rect 2133 4131 2191 4137
rect 2133 4097 2145 4131
rect 2179 4097 2191 4131
rect 2133 4091 2191 4097
rect 2777 4131 2835 4137
rect 2777 4097 2789 4131
rect 2823 4097 2835 4131
rect 2777 4091 2835 4097
rect 2148 3992 2176 4091
rect 2866 4088 2872 4140
rect 2924 4128 2930 4140
rect 3068 4128 3096 4168
rect 3804 4168 5212 4196
rect 43215 4168 43260 4196
rect 3804 4128 3832 4168
rect 2924 4100 2969 4128
rect 3068 4100 3832 4128
rect 2924 4088 2930 4100
rect 2958 4020 2964 4072
rect 3016 4060 3022 4072
rect 3789 4063 3847 4069
rect 3789 4060 3801 4063
rect 3016 4032 3801 4060
rect 3016 4020 3022 4032
rect 3789 4029 3801 4032
rect 3835 4029 3847 4063
rect 3970 4060 3976 4072
rect 3931 4032 3976 4060
rect 3789 4023 3847 4029
rect 3970 4020 3976 4032
rect 4028 4020 4034 4072
rect 4249 4063 4307 4069
rect 4249 4029 4261 4063
rect 4295 4029 4307 4063
rect 5184 4060 5212 4168
rect 43254 4156 43260 4168
rect 43312 4156 43318 4208
rect 45296 4196 45324 4236
rect 48130 4224 48136 4236
rect 48188 4224 48194 4276
rect 45204 4168 45324 4196
rect 45388 4168 46796 4196
rect 5534 4088 5540 4140
rect 5592 4128 5598 4140
rect 6641 4131 6699 4137
rect 6641 4128 6653 4131
rect 5592 4100 6653 4128
rect 5592 4088 5598 4100
rect 6641 4097 6653 4100
rect 6687 4097 6699 4131
rect 6641 4091 6699 4097
rect 6546 4060 6552 4072
rect 5184 4032 6552 4060
rect 4249 4023 4307 4029
rect 2148 3964 3188 3992
rect 2038 3884 2044 3936
rect 2096 3924 2102 3936
rect 2225 3927 2283 3933
rect 2225 3924 2237 3927
rect 2096 3896 2237 3924
rect 2096 3884 2102 3896
rect 2225 3893 2237 3896
rect 2271 3893 2283 3927
rect 3160 3924 3188 3964
rect 3234 3952 3240 4004
rect 3292 3992 3298 4004
rect 4264 3992 4292 4023
rect 6546 4020 6552 4032
rect 6604 4020 6610 4072
rect 6656 4060 6684 4091
rect 9858 4088 9864 4140
rect 9916 4128 9922 4140
rect 10505 4131 10563 4137
rect 10505 4128 10517 4131
rect 9916 4100 10517 4128
rect 9916 4088 9922 4100
rect 10505 4097 10517 4100
rect 10551 4128 10563 4131
rect 19337 4131 19395 4137
rect 10551 4100 16574 4128
rect 10551 4097 10563 4100
rect 10505 4091 10563 4097
rect 13262 4060 13268 4072
rect 6656 4032 13268 4060
rect 13262 4020 13268 4032
rect 13320 4020 13326 4072
rect 16546 4060 16574 4100
rect 19337 4097 19349 4131
rect 19383 4128 19395 4131
rect 19426 4128 19432 4140
rect 19383 4100 19432 4128
rect 19383 4097 19395 4100
rect 19337 4091 19395 4097
rect 19426 4088 19432 4100
rect 19484 4088 19490 4140
rect 39942 4128 39948 4140
rect 39903 4100 39948 4128
rect 39942 4088 39948 4100
rect 40000 4088 40006 4140
rect 41417 4131 41475 4137
rect 41417 4097 41429 4131
rect 41463 4097 41475 4131
rect 43070 4128 43076 4140
rect 43031 4100 43076 4128
rect 41417 4091 41475 4097
rect 17126 4060 17132 4072
rect 16546 4032 17132 4060
rect 17126 4020 17132 4032
rect 17184 4020 17190 4072
rect 19702 4020 19708 4072
rect 19760 4060 19766 4072
rect 20809 4063 20867 4069
rect 20809 4060 20821 4063
rect 19760 4032 20821 4060
rect 19760 4020 19766 4032
rect 20809 4029 20821 4032
rect 20855 4029 20867 4063
rect 20809 4023 20867 4029
rect 22005 4063 22063 4069
rect 22005 4029 22017 4063
rect 22051 4029 22063 4063
rect 22186 4060 22192 4072
rect 22147 4032 22192 4060
rect 22005 4023 22063 4029
rect 3292 3964 4292 3992
rect 3292 3952 3298 3964
rect 10134 3952 10140 4004
rect 10192 3992 10198 4004
rect 22020 3992 22048 4023
rect 22186 4020 22192 4032
rect 22244 4020 22250 4072
rect 22554 4060 22560 4072
rect 22515 4032 22560 4060
rect 22554 4020 22560 4032
rect 22612 4020 22618 4072
rect 10192 3964 22048 3992
rect 39960 3992 39988 4088
rect 41432 4060 41460 4091
rect 43070 4088 43076 4100
rect 43128 4088 43134 4140
rect 45204 4128 45232 4168
rect 45388 4128 45416 4168
rect 44468 4100 45232 4128
rect 45296 4100 45416 4128
rect 46768 4128 46796 4168
rect 47394 4128 47400 4140
rect 46768 4100 47400 4128
rect 41598 4060 41604 4072
rect 41432 4032 41604 4060
rect 41598 4020 41604 4032
rect 41656 4060 41662 4072
rect 44468 4060 44496 4100
rect 44910 4060 44916 4072
rect 41656 4032 44496 4060
rect 44871 4032 44916 4060
rect 41656 4020 41662 4032
rect 44910 4020 44916 4032
rect 44968 4020 44974 4072
rect 45296 3992 45324 4100
rect 47394 4088 47400 4100
rect 47452 4128 47458 4140
rect 47765 4131 47823 4137
rect 47765 4128 47777 4131
rect 47452 4100 47777 4128
rect 47452 4088 47458 4100
rect 47765 4097 47777 4100
rect 47811 4097 47823 4131
rect 47765 4091 47823 4097
rect 45373 4063 45431 4069
rect 45373 4029 45385 4063
rect 45419 4029 45431 4063
rect 45373 4023 45431 4029
rect 45557 4063 45615 4069
rect 45557 4029 45569 4063
rect 45603 4060 45615 4063
rect 46934 4060 46940 4072
rect 45603 4032 46940 4060
rect 45603 4029 45615 4032
rect 45557 4023 45615 4029
rect 39960 3964 45324 3992
rect 45388 3992 45416 4023
rect 46934 4020 46940 4032
rect 46992 4020 46998 4072
rect 47213 4063 47271 4069
rect 47213 4029 47225 4063
rect 47259 4060 47271 4063
rect 47670 4060 47676 4072
rect 47259 4032 47676 4060
rect 47259 4029 47271 4032
rect 47213 4023 47271 4029
rect 47670 4020 47676 4032
rect 47728 4020 47734 4072
rect 47946 3992 47952 4004
rect 45388 3964 47952 3992
rect 10192 3952 10198 3964
rect 47946 3952 47952 3964
rect 48004 3952 48010 4004
rect 5626 3924 5632 3936
rect 3160 3896 5632 3924
rect 2225 3887 2283 3893
rect 5626 3884 5632 3896
rect 5684 3924 5690 3936
rect 6270 3924 6276 3936
rect 5684 3896 6276 3924
rect 5684 3884 5690 3896
rect 6270 3884 6276 3896
rect 6328 3884 6334 3936
rect 6730 3924 6736 3936
rect 6691 3896 6736 3924
rect 6730 3884 6736 3896
rect 6788 3884 6794 3936
rect 7282 3884 7288 3936
rect 7340 3924 7346 3936
rect 7469 3927 7527 3933
rect 7469 3924 7481 3927
rect 7340 3896 7481 3924
rect 7340 3884 7346 3896
rect 7469 3893 7481 3896
rect 7515 3893 7527 3927
rect 7469 3887 7527 3893
rect 10597 3927 10655 3933
rect 10597 3893 10609 3927
rect 10643 3924 10655 3927
rect 10686 3924 10692 3936
rect 10643 3896 10692 3924
rect 10643 3893 10655 3896
rect 10597 3887 10655 3893
rect 10686 3884 10692 3896
rect 10744 3884 10750 3936
rect 12986 3884 12992 3936
rect 13044 3924 13050 3936
rect 13173 3927 13231 3933
rect 13173 3924 13185 3927
rect 13044 3896 13185 3924
rect 13044 3884 13050 3896
rect 13173 3893 13185 3896
rect 13219 3893 13231 3927
rect 13173 3887 13231 3893
rect 16758 3884 16764 3936
rect 16816 3924 16822 3936
rect 17037 3927 17095 3933
rect 17037 3924 17049 3927
rect 16816 3896 17049 3924
rect 16816 3884 16822 3896
rect 17037 3893 17049 3896
rect 17083 3893 17095 3927
rect 17037 3887 17095 3893
rect 17310 3884 17316 3936
rect 17368 3924 17374 3936
rect 18601 3927 18659 3933
rect 18601 3924 18613 3927
rect 17368 3896 18613 3924
rect 17368 3884 17374 3896
rect 18601 3893 18613 3896
rect 18647 3893 18659 3927
rect 18601 3887 18659 3893
rect 19429 3927 19487 3933
rect 19429 3893 19441 3927
rect 19475 3924 19487 3927
rect 19886 3924 19892 3936
rect 19475 3896 19892 3924
rect 19475 3893 19487 3896
rect 19429 3887 19487 3893
rect 19886 3884 19892 3896
rect 19944 3884 19950 3936
rect 20162 3924 20168 3936
rect 20123 3896 20168 3924
rect 20162 3884 20168 3896
rect 20220 3884 20226 3936
rect 24762 3884 24768 3936
rect 24820 3924 24826 3936
rect 25409 3927 25467 3933
rect 25409 3924 25421 3927
rect 24820 3896 25421 3924
rect 24820 3884 24826 3896
rect 25409 3893 25421 3896
rect 25455 3893 25467 3927
rect 25409 3887 25467 3893
rect 25958 3884 25964 3936
rect 26016 3924 26022 3936
rect 26237 3927 26295 3933
rect 26237 3924 26249 3927
rect 26016 3896 26249 3924
rect 26016 3884 26022 3896
rect 26237 3893 26249 3896
rect 26283 3893 26295 3927
rect 26237 3887 26295 3893
rect 27154 3884 27160 3936
rect 27212 3924 27218 3936
rect 27433 3927 27491 3933
rect 27433 3924 27445 3927
rect 27212 3896 27445 3924
rect 27212 3884 27218 3896
rect 27433 3893 27445 3896
rect 27479 3893 27491 3927
rect 27433 3887 27491 3893
rect 40037 3927 40095 3933
rect 40037 3893 40049 3927
rect 40083 3924 40095 3927
rect 40126 3924 40132 3936
rect 40083 3896 40132 3924
rect 40083 3893 40095 3896
rect 40037 3887 40095 3893
rect 40126 3884 40132 3896
rect 40184 3884 40190 3936
rect 40770 3884 40776 3936
rect 40828 3924 40834 3936
rect 40957 3927 41015 3933
rect 40957 3924 40969 3927
rect 40828 3896 40969 3924
rect 40828 3884 40834 3896
rect 40957 3893 40969 3896
rect 41003 3893 41015 3927
rect 40957 3887 41015 3893
rect 41414 3884 41420 3936
rect 41472 3924 41478 3936
rect 41509 3927 41567 3933
rect 41509 3924 41521 3927
rect 41472 3896 41521 3924
rect 41472 3884 41478 3896
rect 41509 3893 41521 3896
rect 41555 3893 41567 3927
rect 41509 3887 41567 3893
rect 46106 3884 46112 3936
rect 46164 3924 46170 3936
rect 47857 3927 47915 3933
rect 47857 3924 47869 3927
rect 46164 3896 47869 3924
rect 46164 3884 46170 3896
rect 47857 3893 47869 3896
rect 47903 3893 47915 3927
rect 47857 3887 47915 3893
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 2777 3723 2835 3729
rect 2777 3689 2789 3723
rect 2823 3720 2835 3723
rect 2958 3720 2964 3732
rect 2823 3692 2964 3720
rect 2823 3689 2835 3692
rect 2777 3683 2835 3689
rect 2958 3680 2964 3692
rect 3016 3680 3022 3732
rect 3329 3723 3387 3729
rect 3329 3689 3341 3723
rect 3375 3720 3387 3723
rect 3970 3720 3976 3732
rect 3375 3692 3976 3720
rect 3375 3689 3387 3692
rect 3329 3683 3387 3689
rect 3970 3680 3976 3692
rect 4028 3680 4034 3732
rect 9582 3720 9588 3732
rect 5092 3692 9588 3720
rect 5092 3652 5120 3692
rect 9582 3680 9588 3692
rect 9640 3680 9646 3732
rect 12894 3680 12900 3732
rect 12952 3720 12958 3732
rect 14182 3720 14188 3732
rect 12952 3692 14188 3720
rect 12952 3680 12958 3692
rect 14182 3680 14188 3692
rect 14240 3680 14246 3732
rect 22002 3720 22008 3732
rect 14292 3692 22008 3720
rect 3252 3624 5120 3652
rect 1946 3516 1952 3528
rect 1907 3488 1952 3516
rect 1946 3476 1952 3488
rect 2004 3476 2010 3528
rect 3252 3525 3280 3624
rect 5166 3612 5172 3664
rect 5224 3652 5230 3664
rect 9858 3652 9864 3664
rect 5224 3624 9864 3652
rect 5224 3612 5230 3624
rect 9858 3612 9864 3624
rect 9916 3612 9922 3664
rect 9968 3624 13032 3652
rect 5442 3584 5448 3596
rect 4080 3556 5448 3584
rect 4080 3525 4108 3556
rect 5442 3544 5448 3556
rect 5500 3544 5506 3596
rect 6454 3584 6460 3596
rect 6415 3556 6460 3584
rect 6454 3544 6460 3556
rect 6512 3544 6518 3596
rect 6546 3544 6552 3596
rect 6604 3584 6610 3596
rect 9968 3584 9996 3624
rect 10686 3584 10692 3596
rect 6604 3556 9996 3584
rect 10647 3556 10692 3584
rect 6604 3544 6610 3556
rect 10686 3544 10692 3556
rect 10744 3544 10750 3596
rect 10962 3584 10968 3596
rect 10923 3556 10968 3584
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 3237 3519 3295 3525
rect 3237 3485 3249 3519
rect 3283 3485 3295 3519
rect 3237 3479 3295 3485
rect 4065 3519 4123 3525
rect 4065 3485 4077 3519
rect 4111 3485 4123 3519
rect 4065 3479 4123 3485
rect 4154 3476 4160 3528
rect 4212 3476 4218 3528
rect 4709 3519 4767 3525
rect 4709 3485 4721 3519
rect 4755 3485 4767 3519
rect 4709 3479 4767 3485
rect 5537 3519 5595 3525
rect 5537 3485 5549 3519
rect 5583 3516 5595 3519
rect 5997 3519 6055 3525
rect 5997 3516 6009 3519
rect 5583 3488 6009 3516
rect 5583 3485 5595 3488
rect 5537 3479 5595 3485
rect 5997 3485 6009 3488
rect 6043 3485 6055 3519
rect 8294 3516 8300 3528
rect 8255 3488 8300 3516
rect 5997 3479 6055 3485
rect 2041 3451 2099 3457
rect 2041 3417 2053 3451
rect 2087 3448 2099 3451
rect 4172 3448 4200 3476
rect 2087 3420 4200 3448
rect 2087 3417 2099 3420
rect 2041 3411 2099 3417
rect 4157 3383 4215 3389
rect 4157 3349 4169 3383
rect 4203 3380 4215 3383
rect 4338 3380 4344 3392
rect 4203 3352 4344 3380
rect 4203 3349 4215 3352
rect 4157 3343 4215 3349
rect 4338 3340 4344 3352
rect 4396 3340 4402 3392
rect 4724 3380 4752 3479
rect 8294 3476 8300 3488
rect 8352 3476 8358 3528
rect 10502 3516 10508 3528
rect 10463 3488 10508 3516
rect 10502 3476 10508 3488
rect 10560 3476 10566 3528
rect 13004 3525 13032 3624
rect 12989 3519 13047 3525
rect 12989 3485 13001 3519
rect 13035 3485 13047 3519
rect 12989 3479 13047 3485
rect 4801 3451 4859 3457
rect 4801 3417 4813 3451
rect 4847 3448 4859 3451
rect 6181 3451 6239 3457
rect 6181 3448 6193 3451
rect 4847 3420 6193 3448
rect 4847 3417 4859 3420
rect 4801 3411 4859 3417
rect 6181 3417 6193 3420
rect 6227 3417 6239 3451
rect 6181 3411 6239 3417
rect 9582 3408 9588 3460
rect 9640 3448 9646 3460
rect 14292 3448 14320 3692
rect 22002 3680 22008 3692
rect 22060 3680 22066 3732
rect 22186 3720 22192 3732
rect 22147 3692 22192 3720
rect 22186 3680 22192 3692
rect 22244 3680 22250 3732
rect 22278 3680 22284 3732
rect 22336 3720 22342 3732
rect 22336 3692 43944 3720
rect 22336 3680 22342 3692
rect 16114 3612 16120 3664
rect 16172 3652 16178 3664
rect 16172 3624 28304 3652
rect 16172 3612 16178 3624
rect 16758 3584 16764 3596
rect 16719 3556 16764 3584
rect 16758 3544 16764 3556
rect 16816 3544 16822 3596
rect 17402 3584 17408 3596
rect 17363 3556 17408 3584
rect 17402 3544 17408 3556
rect 17460 3544 17466 3596
rect 19702 3584 19708 3596
rect 19663 3556 19708 3584
rect 19702 3544 19708 3556
rect 19760 3544 19766 3596
rect 19886 3584 19892 3596
rect 19847 3556 19892 3584
rect 19886 3544 19892 3556
rect 19944 3544 19950 3596
rect 20622 3584 20628 3596
rect 20583 3556 20628 3584
rect 20622 3544 20628 3556
rect 20680 3544 20686 3596
rect 25958 3584 25964 3596
rect 25919 3556 25964 3584
rect 25958 3544 25964 3556
rect 26016 3544 26022 3596
rect 26418 3584 26424 3596
rect 26379 3556 26424 3584
rect 26418 3544 26424 3556
rect 26476 3544 26482 3596
rect 16114 3516 16120 3528
rect 16075 3488 16120 3516
rect 16114 3476 16120 3488
rect 16172 3476 16178 3528
rect 22002 3476 22008 3528
rect 22060 3516 22066 3528
rect 22097 3519 22155 3525
rect 22097 3516 22109 3519
rect 22060 3488 22109 3516
rect 22060 3476 22066 3488
rect 22097 3485 22109 3488
rect 22143 3485 22155 3519
rect 22097 3479 22155 3485
rect 24673 3519 24731 3525
rect 24673 3485 24685 3519
rect 24719 3485 24731 3519
rect 25314 3516 25320 3528
rect 25275 3488 25320 3516
rect 24673 3479 24731 3485
rect 9640 3420 14320 3448
rect 16209 3451 16267 3457
rect 9640 3408 9646 3420
rect 16209 3417 16221 3451
rect 16255 3448 16267 3451
rect 16945 3451 17003 3457
rect 16945 3448 16957 3451
rect 16255 3420 16957 3448
rect 16255 3417 16267 3420
rect 16209 3411 16267 3417
rect 16945 3417 16957 3420
rect 16991 3417 17003 3451
rect 16945 3411 17003 3417
rect 17126 3408 17132 3460
rect 17184 3448 17190 3460
rect 24688 3448 24716 3479
rect 25314 3476 25320 3488
rect 25372 3476 25378 3528
rect 28276 3525 28304 3624
rect 39298 3612 39304 3664
rect 39356 3652 39362 3664
rect 40034 3652 40040 3664
rect 39356 3624 40040 3652
rect 39356 3612 39362 3624
rect 40034 3612 40040 3624
rect 40092 3612 40098 3664
rect 41230 3612 41236 3664
rect 41288 3652 41294 3664
rect 41288 3624 41552 3652
rect 41288 3612 41294 3624
rect 40770 3584 40776 3596
rect 40731 3556 40776 3584
rect 40770 3544 40776 3556
rect 40828 3544 40834 3596
rect 40957 3587 41015 3593
rect 40957 3553 40969 3587
rect 41003 3584 41015 3587
rect 41414 3584 41420 3596
rect 41003 3556 41420 3584
rect 41003 3553 41015 3556
rect 40957 3547 41015 3553
rect 41414 3544 41420 3556
rect 41472 3544 41478 3596
rect 41524 3593 41552 3624
rect 41509 3587 41567 3593
rect 41509 3553 41521 3587
rect 41555 3553 41567 3587
rect 41509 3547 41567 3553
rect 28261 3519 28319 3525
rect 28261 3485 28273 3519
rect 28307 3516 28319 3519
rect 32033 3519 32091 3525
rect 28307 3488 31754 3516
rect 28307 3485 28319 3488
rect 28261 3479 28319 3485
rect 17184 3420 24716 3448
rect 25409 3451 25467 3457
rect 17184 3408 17190 3420
rect 25409 3417 25421 3451
rect 25455 3448 25467 3451
rect 26145 3451 26203 3457
rect 26145 3448 26157 3451
rect 25455 3420 26157 3448
rect 25455 3417 25467 3420
rect 25409 3411 25467 3417
rect 26145 3417 26157 3420
rect 26191 3417 26203 3451
rect 31726 3448 31754 3488
rect 32033 3485 32045 3519
rect 32079 3516 32091 3519
rect 32306 3516 32312 3528
rect 32079 3488 32312 3516
rect 32079 3485 32091 3488
rect 32033 3479 32091 3485
rect 32306 3476 32312 3488
rect 32364 3476 32370 3528
rect 32493 3519 32551 3525
rect 32493 3485 32505 3519
rect 32539 3485 32551 3519
rect 32493 3479 32551 3485
rect 32508 3448 32536 3479
rect 39942 3476 39948 3528
rect 40000 3516 40006 3528
rect 40221 3519 40279 3525
rect 40221 3516 40233 3519
rect 40000 3488 40233 3516
rect 40000 3476 40006 3488
rect 40221 3485 40233 3488
rect 40267 3485 40279 3519
rect 40221 3479 40279 3485
rect 42610 3476 42616 3528
rect 42668 3516 42674 3528
rect 43257 3519 43315 3525
rect 43257 3516 43269 3519
rect 42668 3488 43269 3516
rect 42668 3476 42674 3488
rect 43257 3485 43269 3488
rect 43303 3485 43315 3519
rect 43257 3479 43315 3485
rect 40954 3448 40960 3460
rect 31726 3420 40960 3448
rect 26145 3411 26203 3417
rect 40954 3408 40960 3420
rect 41012 3408 41018 3460
rect 43916 3448 43944 3692
rect 44910 3680 44916 3732
rect 44968 3720 44974 3732
rect 48314 3720 48320 3732
rect 44968 3692 48320 3720
rect 44968 3680 44974 3692
rect 48314 3680 48320 3692
rect 48372 3680 48378 3732
rect 43993 3587 44051 3593
rect 43993 3553 44005 3587
rect 44039 3584 44051 3587
rect 45925 3587 45983 3593
rect 45925 3584 45937 3587
rect 44039 3556 45937 3584
rect 44039 3553 44051 3556
rect 43993 3547 44051 3553
rect 45925 3553 45937 3556
rect 45971 3553 45983 3587
rect 46106 3584 46112 3596
rect 46067 3556 46112 3584
rect 45925 3547 45983 3553
rect 46106 3544 46112 3556
rect 46164 3544 46170 3596
rect 47026 3584 47032 3596
rect 46987 3556 47032 3584
rect 47026 3544 47032 3556
rect 47084 3544 47090 3596
rect 44637 3519 44695 3525
rect 44637 3485 44649 3519
rect 44683 3516 44695 3519
rect 44910 3516 44916 3528
rect 44683 3488 44916 3516
rect 44683 3485 44695 3488
rect 44637 3479 44695 3485
rect 44910 3476 44916 3488
rect 44968 3476 44974 3528
rect 45189 3519 45247 3525
rect 45189 3485 45201 3519
rect 45235 3485 45247 3519
rect 45189 3479 45247 3485
rect 45204 3448 45232 3479
rect 46566 3448 46572 3460
rect 43916 3420 46572 3448
rect 46566 3408 46572 3420
rect 46624 3408 46630 3460
rect 5534 3380 5540 3392
rect 4724 3352 5540 3380
rect 5534 3340 5540 3352
rect 5592 3340 5598 3392
rect 7466 3340 7472 3392
rect 7524 3380 7530 3392
rect 8389 3383 8447 3389
rect 8389 3380 8401 3383
rect 7524 3352 8401 3380
rect 7524 3340 7530 3352
rect 8389 3349 8401 3352
rect 8435 3349 8447 3383
rect 8389 3343 8447 3349
rect 13081 3383 13139 3389
rect 13081 3349 13093 3383
rect 13127 3380 13139 3383
rect 13170 3380 13176 3392
rect 13127 3352 13176 3380
rect 13127 3349 13139 3352
rect 13081 3343 13139 3349
rect 13170 3340 13176 3352
rect 13228 3340 13234 3392
rect 13262 3340 13268 3392
rect 13320 3380 13326 3392
rect 18414 3380 18420 3392
rect 13320 3352 18420 3380
rect 13320 3340 13326 3352
rect 18414 3340 18420 3352
rect 18472 3340 18478 3392
rect 24765 3383 24823 3389
rect 24765 3349 24777 3383
rect 24811 3380 24823 3383
rect 24946 3380 24952 3392
rect 24811 3352 24952 3380
rect 24811 3349 24823 3352
rect 24765 3343 24823 3349
rect 24946 3340 24952 3352
rect 25004 3340 25010 3392
rect 27338 3340 27344 3392
rect 27396 3380 27402 3392
rect 28353 3383 28411 3389
rect 28353 3380 28365 3383
rect 27396 3352 28365 3380
rect 27396 3340 27402 3352
rect 28353 3349 28365 3352
rect 28399 3349 28411 3383
rect 28353 3343 28411 3349
rect 32490 3340 32496 3392
rect 32548 3380 32554 3392
rect 32585 3383 32643 3389
rect 32585 3380 32597 3383
rect 32548 3352 32597 3380
rect 32548 3340 32554 3352
rect 32585 3349 32597 3352
rect 32631 3349 32643 3383
rect 32585 3343 32643 3349
rect 45094 3340 45100 3392
rect 45152 3380 45158 3392
rect 45281 3383 45339 3389
rect 45281 3380 45293 3383
rect 45152 3352 45293 3380
rect 45152 3340 45158 3352
rect 45281 3349 45293 3352
rect 45327 3349 45339 3383
rect 45281 3343 45339 3349
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 1946 3136 1952 3188
rect 2004 3176 2010 3188
rect 5166 3176 5172 3188
rect 2004 3148 5172 3176
rect 2004 3136 2010 3148
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 8294 3136 8300 3188
rect 8352 3176 8358 3188
rect 19426 3176 19432 3188
rect 8352 3148 19432 3176
rect 8352 3136 8358 3148
rect 19426 3136 19432 3148
rect 19484 3136 19490 3188
rect 48958 3176 48964 3188
rect 41386 3148 48964 3176
rect 2038 3108 2044 3120
rect 1999 3080 2044 3108
rect 2038 3068 2044 3080
rect 2096 3068 2102 3120
rect 4338 3108 4344 3120
rect 4299 3080 4344 3108
rect 4338 3068 4344 3080
rect 4396 3068 4402 3120
rect 7466 3108 7472 3120
rect 7427 3080 7472 3108
rect 7466 3068 7472 3080
rect 7524 3068 7530 3120
rect 13170 3108 13176 3120
rect 13131 3080 13176 3108
rect 13170 3068 13176 3080
rect 13228 3068 13234 3120
rect 20162 3108 20168 3120
rect 19628 3080 20168 3108
rect 1854 3040 1860 3052
rect 1815 3012 1860 3040
rect 1854 3000 1860 3012
rect 1912 3000 1918 3052
rect 7282 3040 7288 3052
rect 7243 3012 7288 3040
rect 7282 3000 7288 3012
rect 7340 3000 7346 3052
rect 10502 3000 10508 3052
rect 10560 3040 10566 3052
rect 10689 3043 10747 3049
rect 10689 3040 10701 3043
rect 10560 3012 10701 3040
rect 10560 3000 10566 3012
rect 10689 3009 10701 3012
rect 10735 3009 10747 3043
rect 12986 3040 12992 3052
rect 12947 3012 12992 3040
rect 10689 3003 10747 3009
rect 12986 3000 12992 3012
rect 13044 3000 13050 3052
rect 17310 3040 17316 3052
rect 17271 3012 17316 3040
rect 17310 3000 17316 3012
rect 17368 3000 17374 3052
rect 19628 3049 19656 3080
rect 20162 3068 20168 3080
rect 20220 3068 20226 3120
rect 24946 3108 24952 3120
rect 24907 3080 24952 3108
rect 24946 3068 24952 3080
rect 25004 3068 25010 3120
rect 27338 3108 27344 3120
rect 27299 3080 27344 3108
rect 27338 3068 27344 3080
rect 27396 3068 27402 3120
rect 32490 3108 32496 3120
rect 32451 3080 32496 3108
rect 32490 3068 32496 3080
rect 32548 3068 32554 3120
rect 40126 3108 40132 3120
rect 40087 3080 40132 3108
rect 40126 3068 40132 3080
rect 40184 3068 40190 3120
rect 19613 3043 19671 3049
rect 19613 3009 19625 3043
rect 19659 3009 19671 3043
rect 24762 3040 24768 3052
rect 24723 3012 24768 3040
rect 19613 3003 19671 3009
rect 24762 3000 24768 3012
rect 24820 3000 24826 3052
rect 27154 3040 27160 3052
rect 27115 3012 27160 3040
rect 27154 3000 27160 3012
rect 27212 3000 27218 3052
rect 32306 3040 32312 3052
rect 32267 3012 32312 3040
rect 32306 3000 32312 3012
rect 32364 3000 32370 3052
rect 39942 3040 39948 3052
rect 39903 3012 39948 3040
rect 39942 3000 39948 3012
rect 40000 3000 40006 3052
rect 2774 2972 2780 2984
rect 2735 2944 2780 2972
rect 2774 2932 2780 2944
rect 2832 2932 2838 2984
rect 4157 2975 4215 2981
rect 4157 2941 4169 2975
rect 4203 2972 4215 2975
rect 4982 2972 4988 2984
rect 4203 2944 4988 2972
rect 4203 2941 4215 2944
rect 4157 2935 4215 2941
rect 4982 2932 4988 2944
rect 5040 2932 5046 2984
rect 5166 2972 5172 2984
rect 5127 2944 5172 2972
rect 5166 2932 5172 2944
rect 5224 2932 5230 2984
rect 7742 2972 7748 2984
rect 7703 2944 7748 2972
rect 7742 2932 7748 2944
rect 7800 2932 7806 2984
rect 13538 2972 13544 2984
rect 13499 2944 13544 2972
rect 13538 2932 13544 2944
rect 13596 2932 13602 2984
rect 17497 2975 17555 2981
rect 17497 2941 17509 2975
rect 17543 2972 17555 2975
rect 18506 2972 18512 2984
rect 17543 2944 18512 2972
rect 17543 2941 17555 2944
rect 17497 2935 17555 2941
rect 18506 2932 18512 2944
rect 18564 2932 18570 2984
rect 19153 2975 19211 2981
rect 19153 2941 19165 2975
rect 19199 2972 19211 2975
rect 19334 2972 19340 2984
rect 19199 2944 19340 2972
rect 19199 2941 19211 2944
rect 19153 2935 19211 2941
rect 19334 2932 19340 2944
rect 19392 2932 19398 2984
rect 19794 2972 19800 2984
rect 19755 2944 19800 2972
rect 19794 2932 19800 2944
rect 19852 2932 19858 2984
rect 21453 2975 21511 2981
rect 21453 2941 21465 2975
rect 21499 2941 21511 2975
rect 25774 2972 25780 2984
rect 25735 2944 25780 2972
rect 21453 2935 21511 2941
rect 21468 2904 21496 2935
rect 25774 2932 25780 2944
rect 25832 2932 25838 2984
rect 27706 2972 27712 2984
rect 27667 2944 27712 2972
rect 27706 2932 27712 2944
rect 27764 2932 27770 2984
rect 32214 2932 32220 2984
rect 32272 2972 32278 2984
rect 32769 2975 32827 2981
rect 32769 2972 32781 2975
rect 32272 2944 32781 2972
rect 32272 2932 32278 2944
rect 32769 2941 32781 2944
rect 32815 2941 32827 2975
rect 40586 2972 40592 2984
rect 40547 2944 40592 2972
rect 32769 2935 32827 2941
rect 40586 2932 40592 2944
rect 40644 2932 40650 2984
rect 41386 2904 41414 3148
rect 48958 3136 48964 3148
rect 49016 3136 49022 3188
rect 45094 3108 45100 3120
rect 45055 3080 45100 3108
rect 45094 3068 45100 3080
rect 45152 3068 45158 3120
rect 42610 3040 42616 3052
rect 42571 3012 42616 3040
rect 42610 3000 42616 3012
rect 42668 3000 42674 3052
rect 44910 3040 44916 3052
rect 44871 3012 44916 3040
rect 44910 3000 44916 3012
rect 44968 3000 44974 3052
rect 48038 3040 48044 3052
rect 47999 3012 48044 3040
rect 48038 3000 48044 3012
rect 48096 3000 48102 3052
rect 42797 2975 42855 2981
rect 42797 2941 42809 2975
rect 42843 2972 42855 2975
rect 42886 2972 42892 2984
rect 42843 2944 42892 2972
rect 42843 2941 42855 2944
rect 42797 2935 42855 2941
rect 42886 2932 42892 2944
rect 42944 2932 42950 2984
rect 43073 2975 43131 2981
rect 43073 2941 43085 2975
rect 43119 2941 43131 2975
rect 45738 2972 45744 2984
rect 45699 2944 45744 2972
rect 43073 2935 43131 2941
rect 21468 2876 41414 2904
rect 41874 2864 41880 2916
rect 41932 2904 41938 2916
rect 43088 2904 43116 2935
rect 45738 2932 45744 2944
rect 45796 2932 45802 2984
rect 41932 2876 43116 2904
rect 41932 2864 41938 2876
rect 45094 2864 45100 2916
rect 45152 2904 45158 2916
rect 45646 2904 45652 2916
rect 45152 2876 45652 2904
rect 45152 2864 45158 2876
rect 45646 2864 45652 2876
rect 45704 2864 45710 2916
rect 6822 2836 6828 2848
rect 6783 2808 6828 2836
rect 6822 2796 6828 2808
rect 6880 2796 6886 2848
rect 28350 2796 28356 2848
rect 28408 2836 28414 2848
rect 48225 2839 48283 2845
rect 48225 2836 48237 2839
rect 28408 2808 48237 2836
rect 28408 2796 28414 2808
rect 48225 2805 48237 2808
rect 48271 2805 48283 2839
rect 48225 2799 48283 2805
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 1949 2635 2007 2641
rect 1949 2601 1961 2635
rect 1995 2632 2007 2635
rect 14461 2635 14519 2641
rect 1995 2604 11744 2632
rect 1995 2601 2007 2604
rect 1949 2595 2007 2601
rect 4614 2564 4620 2576
rect 3988 2536 4620 2564
rect 3988 2505 4016 2536
rect 4614 2524 4620 2536
rect 4672 2524 4678 2576
rect 3973 2499 4031 2505
rect 3973 2465 3985 2499
rect 4019 2465 4031 2499
rect 4154 2496 4160 2508
rect 4115 2468 4160 2496
rect 3973 2459 4031 2465
rect 4154 2456 4160 2468
rect 4212 2456 4218 2508
rect 4522 2496 4528 2508
rect 4483 2468 4528 2496
rect 4522 2456 4528 2468
rect 4580 2456 4586 2508
rect 6641 2499 6699 2505
rect 6641 2465 6653 2499
rect 6687 2496 6699 2499
rect 6822 2496 6828 2508
rect 6687 2468 6828 2496
rect 6687 2465 6699 2468
rect 6641 2459 6699 2465
rect 6822 2456 6828 2468
rect 6880 2456 6886 2508
rect 7098 2496 7104 2508
rect 7059 2468 7104 2496
rect 7098 2456 7104 2468
rect 7156 2456 7162 2508
rect 11716 2496 11744 2604
rect 14461 2601 14473 2635
rect 14507 2632 14519 2635
rect 17586 2632 17592 2644
rect 14507 2604 17592 2632
rect 14507 2601 14519 2604
rect 14461 2595 14519 2601
rect 17586 2592 17592 2604
rect 17644 2592 17650 2644
rect 18506 2632 18512 2644
rect 18467 2604 18512 2632
rect 18506 2592 18512 2604
rect 18564 2592 18570 2644
rect 19521 2635 19579 2641
rect 19521 2601 19533 2635
rect 19567 2632 19579 2635
rect 19794 2632 19800 2644
rect 19567 2604 19800 2632
rect 19567 2601 19579 2604
rect 19521 2595 19579 2601
rect 19794 2592 19800 2604
rect 19852 2592 19858 2644
rect 41693 2635 41751 2641
rect 41693 2601 41705 2635
rect 41739 2632 41751 2635
rect 42886 2632 42892 2644
rect 41739 2604 42892 2632
rect 41739 2601 41751 2604
rect 41693 2595 41751 2601
rect 42886 2592 42892 2604
rect 42944 2592 42950 2644
rect 47946 2632 47952 2644
rect 47907 2604 47952 2632
rect 47946 2592 47952 2604
rect 48004 2592 48010 2644
rect 11885 2567 11943 2573
rect 11885 2533 11897 2567
rect 11931 2564 11943 2567
rect 17770 2564 17776 2576
rect 11931 2536 17776 2564
rect 11931 2533 11943 2536
rect 11885 2527 11943 2533
rect 17770 2524 17776 2536
rect 17828 2524 17834 2576
rect 25038 2564 25044 2576
rect 20272 2536 25044 2564
rect 20272 2496 20300 2536
rect 25038 2524 25044 2536
rect 25096 2524 25102 2576
rect 39574 2524 39580 2576
rect 39632 2564 39638 2576
rect 44177 2567 44235 2573
rect 44177 2564 44189 2567
rect 39632 2536 44189 2564
rect 39632 2524 39638 2536
rect 44177 2533 44189 2536
rect 44223 2533 44235 2567
rect 44177 2527 44235 2533
rect 11716 2468 20300 2496
rect 20349 2499 20407 2505
rect 20349 2465 20361 2499
rect 20395 2496 20407 2499
rect 26050 2496 26056 2508
rect 20395 2468 26056 2496
rect 20395 2465 20407 2468
rect 20349 2459 20407 2465
rect 26050 2456 26056 2468
rect 26108 2456 26114 2508
rect 44634 2456 44640 2508
rect 44692 2496 44698 2508
rect 45373 2499 45431 2505
rect 45373 2496 45385 2499
rect 44692 2468 45385 2496
rect 44692 2456 44698 2468
rect 45373 2465 45385 2468
rect 45419 2465 45431 2499
rect 45373 2459 45431 2465
rect 45557 2499 45615 2505
rect 45557 2465 45569 2499
rect 45603 2496 45615 2499
rect 46474 2496 46480 2508
rect 45603 2468 46480 2496
rect 45603 2465 45615 2468
rect 45557 2459 45615 2465
rect 46474 2456 46480 2468
rect 46532 2456 46538 2508
rect 46842 2496 46848 2508
rect 46803 2468 46848 2496
rect 46842 2456 46848 2468
rect 46900 2456 46906 2508
rect 11606 2388 11612 2440
rect 11664 2428 11670 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11664 2400 11713 2428
rect 11664 2388 11670 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 14182 2388 14188 2440
rect 14240 2428 14246 2440
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 14240 2400 14289 2428
rect 14240 2388 14246 2400
rect 14277 2397 14289 2400
rect 14323 2397 14335 2431
rect 18414 2428 18420 2440
rect 18327 2400 18420 2428
rect 14277 2391 14335 2397
rect 18414 2388 18420 2400
rect 18472 2388 18478 2440
rect 19426 2428 19432 2440
rect 19387 2400 19432 2428
rect 19426 2388 19432 2400
rect 19484 2388 19490 2440
rect 19978 2388 19984 2440
rect 20036 2428 20042 2440
rect 20073 2431 20131 2437
rect 20073 2428 20085 2431
rect 20036 2400 20085 2428
rect 20036 2388 20042 2400
rect 20073 2397 20085 2400
rect 20119 2397 20131 2431
rect 20073 2391 20131 2397
rect 38654 2388 38660 2440
rect 38712 2428 38718 2440
rect 38749 2431 38807 2437
rect 38749 2428 38761 2431
rect 38712 2400 38761 2428
rect 38712 2388 38718 2400
rect 38749 2397 38761 2400
rect 38795 2397 38807 2431
rect 41598 2428 41604 2440
rect 41559 2400 41604 2428
rect 38749 2391 38807 2397
rect 41598 2388 41604 2400
rect 41656 2388 41662 2440
rect 1302 2320 1308 2372
rect 1360 2360 1366 2372
rect 1673 2363 1731 2369
rect 1673 2360 1685 2363
rect 1360 2332 1685 2360
rect 1360 2320 1366 2332
rect 1673 2329 1685 2332
rect 1719 2329 1731 2363
rect 1673 2323 1731 2329
rect 2593 2363 2651 2369
rect 2593 2329 2605 2363
rect 2639 2360 2651 2363
rect 2774 2360 2780 2372
rect 2639 2332 2780 2360
rect 2639 2329 2651 2332
rect 2593 2323 2651 2329
rect 2774 2320 2780 2332
rect 2832 2320 2838 2372
rect 6822 2360 6828 2372
rect 6783 2332 6828 2360
rect 6822 2320 6828 2332
rect 6880 2320 6886 2372
rect 18432 2360 18460 2388
rect 25314 2360 25320 2372
rect 18432 2332 25320 2360
rect 25314 2320 25320 2332
rect 25372 2320 25378 2372
rect 28994 2320 29000 2372
rect 29052 2360 29058 2372
rect 29825 2363 29883 2369
rect 29825 2360 29837 2363
rect 29052 2332 29837 2360
rect 29052 2320 29058 2332
rect 29825 2329 29837 2332
rect 29871 2329 29883 2363
rect 29825 2323 29883 2329
rect 43806 2320 43812 2372
rect 43864 2360 43870 2372
rect 43993 2363 44051 2369
rect 43993 2360 44005 2363
rect 43864 2332 44005 2360
rect 43864 2320 43870 2332
rect 43993 2329 44005 2332
rect 44039 2329 44051 2363
rect 43993 2323 44051 2329
rect 2866 2292 2872 2304
rect 2827 2264 2872 2292
rect 2866 2252 2872 2264
rect 2924 2252 2930 2304
rect 23842 2252 23848 2304
rect 23900 2292 23906 2304
rect 29917 2295 29975 2301
rect 29917 2292 29929 2295
rect 23900 2264 29929 2292
rect 23900 2252 23906 2264
rect 29917 2261 29929 2264
rect 29963 2261 29975 2295
rect 29917 2255 29975 2261
rect 32858 2252 32864 2304
rect 32916 2292 32922 2304
rect 38933 2295 38991 2301
rect 38933 2292 38945 2295
rect 32916 2264 38945 2292
rect 32916 2252 32922 2264
rect 38933 2261 38945 2264
rect 38979 2261 38991 2295
rect 38933 2255 38991 2261
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
rect 2866 1980 2872 2032
rect 2924 2020 2930 2032
rect 17494 2020 17500 2032
rect 2924 1992 17500 2020
rect 2924 1980 2930 1992
rect 17494 1980 17500 1992
rect 17552 1980 17558 2032
rect 2866 1844 2872 1896
rect 2924 1884 2930 1896
rect 5350 1884 5356 1896
rect 2924 1856 5356 1884
rect 2924 1844 2930 1856
rect 5350 1844 5356 1856
rect 5408 1844 5414 1896
<< via1 >>
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 17960 47132 18012 47184
rect 32220 47132 32272 47184
rect 42892 47132 42944 47184
rect 4160 47064 4212 47116
rect 2136 47039 2188 47048
rect 2136 47005 2145 47039
rect 2145 47005 2179 47039
rect 2179 47005 2188 47039
rect 2136 46996 2188 47005
rect 4068 46996 4120 47048
rect 7196 47064 7248 47116
rect 9036 47064 9088 47116
rect 14188 47064 14240 47116
rect 47216 47107 47268 47116
rect 47216 47073 47225 47107
rect 47225 47073 47259 47107
rect 47259 47073 47268 47107
rect 47216 47064 47268 47073
rect 5356 46996 5408 47048
rect 6552 47039 6604 47048
rect 6552 47005 6561 47039
rect 6561 47005 6595 47039
rect 6595 47005 6604 47039
rect 6552 46996 6604 47005
rect 7380 47039 7432 47048
rect 7380 47005 7389 47039
rect 7389 47005 7423 47039
rect 7423 47005 7432 47039
rect 7380 46996 7432 47005
rect 8852 46996 8904 47048
rect 12716 47039 12768 47048
rect 12716 47005 12725 47039
rect 12725 47005 12759 47039
rect 12759 47005 12768 47039
rect 12716 46996 12768 47005
rect 17408 46996 17460 47048
rect 19340 46996 19392 47048
rect 22468 46996 22520 47048
rect 23848 46996 23900 47048
rect 25688 47039 25740 47048
rect 25688 47005 25697 47039
rect 25697 47005 25731 47039
rect 25731 47005 25740 47039
rect 25688 46996 25740 47005
rect 29736 46996 29788 47048
rect 31760 46996 31812 47048
rect 33232 47039 33284 47048
rect 33232 47005 33241 47039
rect 33241 47005 33275 47039
rect 33275 47005 33284 47039
rect 33232 46996 33284 47005
rect 39764 46996 39816 47048
rect 40224 47039 40276 47048
rect 40224 47005 40233 47039
rect 40233 47005 40267 47039
rect 40267 47005 40276 47039
rect 40224 46996 40276 47005
rect 41420 47039 41472 47048
rect 41420 47005 41429 47039
rect 41429 47005 41463 47039
rect 41463 47005 41472 47039
rect 41420 46996 41472 47005
rect 42524 46996 42576 47048
rect 45376 47039 45428 47048
rect 45376 47005 45385 47039
rect 45385 47005 45419 47039
rect 45419 47005 45428 47039
rect 45376 46996 45428 47005
rect 48964 46996 49016 47048
rect 4804 46971 4856 46980
rect 4804 46937 4813 46971
rect 4813 46937 4847 46971
rect 4847 46937 4856 46971
rect 4804 46928 4856 46937
rect 5632 46928 5684 46980
rect 13820 46928 13872 46980
rect 19708 46971 19760 46980
rect 19708 46937 19717 46971
rect 19717 46937 19751 46971
rect 19751 46937 19760 46971
rect 19708 46928 19760 46937
rect 25412 46928 25464 46980
rect 45560 46971 45612 46980
rect 45560 46937 45569 46971
rect 45569 46937 45603 46971
rect 45603 46937 45612 46971
rect 45560 46928 45612 46937
rect 5540 46903 5592 46912
rect 5540 46869 5549 46903
rect 5549 46869 5583 46903
rect 5583 46869 5592 46903
rect 5540 46860 5592 46869
rect 46388 46860 46440 46912
rect 46940 46860 46992 46912
rect 48044 46903 48096 46912
rect 48044 46869 48053 46903
rect 48053 46869 48087 46903
rect 48087 46869 48096 46903
rect 48044 46860 48096 46869
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 2596 46588 2648 46640
rect 4160 46563 4212 46572
rect 4160 46529 4169 46563
rect 4169 46529 4203 46563
rect 4203 46529 4212 46563
rect 4160 46520 4212 46529
rect 12716 46588 12768 46640
rect 22468 46563 22520 46572
rect 22468 46529 22477 46563
rect 22477 46529 22511 46563
rect 22511 46529 22520 46563
rect 22468 46520 22520 46529
rect 25688 46588 25740 46640
rect 33232 46588 33284 46640
rect 48320 46588 48372 46640
rect 39764 46563 39816 46572
rect 39764 46529 39773 46563
rect 39773 46529 39807 46563
rect 39807 46529 39816 46563
rect 39764 46520 39816 46529
rect 41420 46520 41472 46572
rect 47768 46563 47820 46572
rect 47768 46529 47777 46563
rect 47777 46529 47811 46563
rect 47811 46529 47820 46563
rect 47768 46520 47820 46529
rect 2044 46495 2096 46504
rect 2044 46461 2053 46495
rect 2053 46461 2087 46495
rect 2087 46461 2096 46495
rect 2044 46452 2096 46461
rect 2320 46495 2372 46504
rect 2320 46461 2329 46495
rect 2329 46461 2363 46495
rect 2363 46461 2372 46495
rect 2320 46452 2372 46461
rect 5908 46452 5960 46504
rect 12532 46452 12584 46504
rect 12900 46495 12952 46504
rect 12900 46461 12909 46495
rect 12909 46461 12943 46495
rect 12943 46461 12952 46495
rect 12900 46452 12952 46461
rect 14280 46495 14332 46504
rect 14280 46461 14289 46495
rect 14289 46461 14323 46495
rect 14323 46461 14332 46495
rect 14280 46452 14332 46461
rect 14464 46495 14516 46504
rect 14464 46461 14473 46495
rect 14473 46461 14507 46495
rect 14507 46461 14516 46495
rect 14464 46452 14516 46461
rect 14832 46495 14884 46504
rect 14832 46461 14841 46495
rect 14841 46461 14875 46495
rect 14875 46461 14884 46495
rect 14832 46452 14884 46461
rect 22744 46452 22796 46504
rect 23204 46495 23256 46504
rect 23204 46461 23213 46495
rect 23213 46461 23247 46495
rect 23247 46461 23256 46495
rect 23204 46452 23256 46461
rect 24952 46495 25004 46504
rect 24952 46461 24961 46495
rect 24961 46461 24995 46495
rect 24995 46461 25004 46495
rect 24952 46452 25004 46461
rect 25780 46495 25832 46504
rect 25780 46461 25789 46495
rect 25789 46461 25823 46495
rect 25823 46461 25832 46495
rect 25780 46452 25832 46461
rect 29184 46495 29236 46504
rect 29184 46461 29193 46495
rect 29193 46461 29227 46495
rect 29227 46461 29236 46495
rect 29184 46452 29236 46461
rect 29644 46495 29696 46504
rect 29644 46461 29653 46495
rect 29653 46461 29687 46495
rect 29687 46461 29696 46495
rect 29644 46452 29696 46461
rect 33140 46452 33192 46504
rect 33508 46495 33560 46504
rect 33508 46461 33517 46495
rect 33517 46461 33551 46495
rect 33551 46461 33560 46495
rect 33508 46452 33560 46461
rect 37648 46495 37700 46504
rect 37648 46461 37657 46495
rect 37657 46461 37691 46495
rect 37691 46461 37700 46495
rect 37648 46452 37700 46461
rect 39948 46495 40000 46504
rect 36728 46384 36780 46436
rect 39948 46461 39957 46495
rect 39957 46461 39991 46495
rect 39991 46461 40000 46495
rect 39948 46452 40000 46461
rect 42800 46495 42852 46504
rect 38660 46384 38712 46436
rect 42800 46461 42809 46495
rect 42809 46461 42843 46495
rect 42843 46461 42852 46495
rect 42800 46452 42852 46461
rect 45376 46495 45428 46504
rect 41880 46384 41932 46436
rect 45376 46461 45385 46495
rect 45385 46461 45419 46495
rect 45419 46461 45428 46495
rect 45376 46452 45428 46461
rect 47032 46452 47084 46504
rect 5264 46316 5316 46368
rect 8024 46359 8076 46368
rect 8024 46325 8033 46359
rect 8033 46325 8067 46359
rect 8067 46325 8076 46359
rect 8024 46316 8076 46325
rect 15016 46316 15068 46368
rect 35440 46316 35492 46368
rect 46664 46316 46716 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 2044 46112 2096 46164
rect 12532 46155 12584 46164
rect 12532 46121 12541 46155
rect 12541 46121 12575 46155
rect 12575 46121 12584 46155
rect 12532 46112 12584 46121
rect 13820 46112 13872 46164
rect 14464 46155 14516 46164
rect 14464 46121 14473 46155
rect 14473 46121 14507 46155
rect 14507 46121 14516 46155
rect 14464 46112 14516 46121
rect 22744 46155 22796 46164
rect 22744 46121 22753 46155
rect 22753 46121 22787 46155
rect 22787 46121 22796 46155
rect 22744 46112 22796 46121
rect 29184 46112 29236 46164
rect 33140 46155 33192 46164
rect 33140 46121 33149 46155
rect 33149 46121 33183 46155
rect 33183 46121 33192 46155
rect 33140 46112 33192 46121
rect 39948 46112 40000 46164
rect 45376 46155 45428 46164
rect 45376 46121 45385 46155
rect 45385 46121 45419 46155
rect 45419 46121 45428 46155
rect 45376 46112 45428 46121
rect 45560 46112 45612 46164
rect 8024 46044 8076 46096
rect 2780 46019 2832 46028
rect 2780 45985 2789 46019
rect 2789 45985 2823 46019
rect 2823 45985 2832 46019
rect 2780 45976 2832 45985
rect 5264 46019 5316 46028
rect 5264 45985 5273 46019
rect 5273 45985 5307 46019
rect 5307 45985 5316 46019
rect 5264 45976 5316 45985
rect 5540 45976 5592 46028
rect 5816 46019 5868 46028
rect 5816 45985 5825 46019
rect 5825 45985 5859 46019
rect 5859 45985 5868 46019
rect 5816 45976 5868 45985
rect 41328 46044 41380 46096
rect 15016 46019 15068 46028
rect 15016 45985 15025 46019
rect 15025 45985 15059 46019
rect 15059 45985 15068 46019
rect 15016 45976 15068 45985
rect 15476 46019 15528 46028
rect 15476 45985 15485 46019
rect 15485 45985 15519 46019
rect 15519 45985 15528 46019
rect 15476 45976 15528 45985
rect 19064 45976 19116 46028
rect 35440 46019 35492 46028
rect 4068 45951 4120 45960
rect 4068 45917 4077 45951
rect 4077 45917 4111 45951
rect 4111 45917 4120 45951
rect 4068 45908 4120 45917
rect 6920 45908 6972 45960
rect 4620 45883 4672 45892
rect 4620 45849 4629 45883
rect 4629 45849 4663 45883
rect 4663 45849 4672 45883
rect 4620 45840 4672 45849
rect 4896 45840 4948 45892
rect 5540 45840 5592 45892
rect 12440 45951 12492 45960
rect 12440 45917 12449 45951
rect 12449 45917 12483 45951
rect 12483 45917 12492 45951
rect 12440 45908 12492 45917
rect 22652 45951 22704 45960
rect 7288 45772 7340 45824
rect 22652 45917 22661 45951
rect 22661 45917 22695 45951
rect 22695 45917 22704 45951
rect 22652 45908 22704 45917
rect 29184 45908 29236 45960
rect 29736 45951 29788 45960
rect 29736 45917 29745 45951
rect 29745 45917 29779 45951
rect 29779 45917 29788 45951
rect 29736 45908 29788 45917
rect 32956 45908 33008 45960
rect 15200 45883 15252 45892
rect 15200 45849 15209 45883
rect 15209 45849 15243 45883
rect 15243 45849 15252 45883
rect 15200 45840 15252 45849
rect 24860 45883 24912 45892
rect 24860 45849 24869 45883
rect 24869 45849 24903 45883
rect 24903 45849 24912 45883
rect 24860 45840 24912 45849
rect 25136 45840 25188 45892
rect 29920 45883 29972 45892
rect 29920 45849 29929 45883
rect 29929 45849 29963 45883
rect 29963 45849 29972 45883
rect 29920 45840 29972 45849
rect 30288 45840 30340 45892
rect 34520 45772 34572 45824
rect 35440 45985 35449 46019
rect 35449 45985 35483 46019
rect 35483 45985 35492 46019
rect 35440 45976 35492 45985
rect 36084 46019 36136 46028
rect 36084 45985 36093 46019
rect 36093 45985 36127 46019
rect 36127 45985 36136 46019
rect 36084 45976 36136 45985
rect 40224 45976 40276 46028
rect 40592 46019 40644 46028
rect 40592 45985 40601 46019
rect 40601 45985 40635 46019
rect 40635 45985 40644 46019
rect 40592 45976 40644 45985
rect 46664 46019 46716 46028
rect 46664 45985 46673 46019
rect 46673 45985 46707 46019
rect 46707 45985 46716 46019
rect 46664 45976 46716 45985
rect 48228 46019 48280 46028
rect 48228 45985 48237 46019
rect 48237 45985 48271 46019
rect 48271 45985 48280 46019
rect 48228 45976 48280 45985
rect 38660 45908 38712 45960
rect 39948 45908 40000 45960
rect 45836 45951 45888 45960
rect 45836 45917 45845 45951
rect 45845 45917 45879 45951
rect 45879 45917 45888 45951
rect 45836 45908 45888 45917
rect 46480 45951 46532 45960
rect 46480 45917 46489 45951
rect 46489 45917 46523 45951
rect 46523 45917 46532 45951
rect 46480 45908 46532 45917
rect 35624 45883 35676 45892
rect 35624 45849 35633 45883
rect 35633 45849 35667 45883
rect 35667 45849 35676 45883
rect 35624 45840 35676 45849
rect 40224 45883 40276 45892
rect 40224 45849 40233 45883
rect 40233 45849 40267 45883
rect 40267 45849 40276 45883
rect 40224 45840 40276 45849
rect 46572 45772 46624 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 4620 45568 4672 45620
rect 10048 45568 10100 45620
rect 15200 45568 15252 45620
rect 5632 45500 5684 45552
rect 5908 45500 5960 45552
rect 7288 45543 7340 45552
rect 7288 45509 7297 45543
rect 7297 45509 7331 45543
rect 7331 45509 7340 45543
rect 7288 45500 7340 45509
rect 22652 45568 22704 45620
rect 24860 45611 24912 45620
rect 24860 45577 24869 45611
rect 24869 45577 24903 45611
rect 24903 45577 24912 45611
rect 24860 45568 24912 45577
rect 24952 45568 25004 45620
rect 29920 45568 29972 45620
rect 32956 45568 33008 45620
rect 35624 45568 35676 45620
rect 40224 45568 40276 45620
rect 4896 45432 4948 45484
rect 7196 45475 7248 45484
rect 2964 45407 3016 45416
rect 2964 45373 2973 45407
rect 2973 45373 3007 45407
rect 3007 45373 3016 45407
rect 2964 45364 3016 45373
rect 5448 45407 5500 45416
rect 5448 45373 5457 45407
rect 5457 45373 5491 45407
rect 5491 45373 5500 45407
rect 5448 45364 5500 45373
rect 7196 45441 7205 45475
rect 7205 45441 7239 45475
rect 7239 45441 7248 45475
rect 37648 45500 37700 45552
rect 42800 45500 42852 45552
rect 45928 45500 45980 45552
rect 47032 45543 47084 45552
rect 7196 45432 7248 45441
rect 14280 45432 14332 45484
rect 15200 45475 15252 45484
rect 15200 45441 15209 45475
rect 15209 45441 15243 45475
rect 15243 45441 15252 45475
rect 15200 45432 15252 45441
rect 29184 45432 29236 45484
rect 29736 45475 29788 45484
rect 29736 45441 29745 45475
rect 29745 45441 29779 45475
rect 29779 45441 29788 45475
rect 29736 45432 29788 45441
rect 34520 45432 34572 45484
rect 35624 45432 35676 45484
rect 38660 45432 38712 45484
rect 39948 45475 40000 45484
rect 39948 45441 39957 45475
rect 39957 45441 39991 45475
rect 39991 45441 40000 45475
rect 39948 45432 40000 45441
rect 40592 45432 40644 45484
rect 41328 45475 41380 45484
rect 41328 45441 41337 45475
rect 41337 45441 41371 45475
rect 41371 45441 41380 45475
rect 41328 45432 41380 45441
rect 45468 45432 45520 45484
rect 46480 45475 46532 45484
rect 46480 45441 46489 45475
rect 46489 45441 46523 45475
rect 46523 45441 46532 45475
rect 46480 45432 46532 45441
rect 47032 45509 47041 45543
rect 47041 45509 47075 45543
rect 47075 45509 47084 45543
rect 47032 45500 47084 45509
rect 47768 45432 47820 45484
rect 7380 45296 7432 45348
rect 15200 45296 15252 45348
rect 10508 45228 10560 45280
rect 47768 45296 47820 45348
rect 46480 45228 46532 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 6828 44931 6880 44940
rect 6828 44897 6837 44931
rect 6837 44897 6871 44931
rect 6871 44897 6880 44931
rect 6828 44888 6880 44897
rect 10508 44931 10560 44940
rect 10508 44897 10517 44931
rect 10517 44897 10551 44931
rect 10551 44897 10560 44931
rect 10508 44888 10560 44897
rect 11060 44931 11112 44940
rect 11060 44897 11069 44931
rect 11069 44897 11103 44931
rect 11103 44897 11112 44931
rect 11060 44888 11112 44897
rect 40592 44931 40644 44940
rect 40592 44897 40601 44931
rect 40601 44897 40635 44931
rect 40635 44897 40644 44931
rect 40592 44888 40644 44897
rect 46480 44931 46532 44940
rect 46480 44897 46489 44931
rect 46489 44897 46523 44931
rect 46523 44897 46532 44931
rect 46480 44888 46532 44897
rect 48228 44931 48280 44940
rect 48228 44897 48237 44931
rect 48237 44897 48271 44931
rect 48271 44897 48280 44931
rect 48228 44888 48280 44897
rect 20 44820 72 44872
rect 4068 44820 4120 44872
rect 4896 44820 4948 44872
rect 40040 44863 40092 44872
rect 40040 44829 40049 44863
rect 40049 44829 40083 44863
rect 40083 44829 40092 44863
rect 40040 44820 40092 44829
rect 45836 44820 45888 44872
rect 3792 44752 3844 44804
rect 5356 44752 5408 44804
rect 10692 44795 10744 44804
rect 10692 44761 10701 44795
rect 10701 44761 10735 44795
rect 10735 44761 10744 44795
rect 10692 44752 10744 44761
rect 47860 44752 47912 44804
rect 1768 44727 1820 44736
rect 1768 44693 1777 44727
rect 1777 44693 1811 44727
rect 1811 44693 1820 44727
rect 1768 44684 1820 44693
rect 5264 44727 5316 44736
rect 5264 44693 5273 44727
rect 5273 44693 5307 44727
rect 5307 44693 5316 44727
rect 5264 44684 5316 44693
rect 12440 44684 12492 44736
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 10692 44480 10744 44532
rect 47860 44523 47912 44532
rect 47860 44489 47869 44523
rect 47869 44489 47903 44523
rect 47903 44489 47912 44523
rect 47860 44480 47912 44489
rect 4896 44387 4948 44396
rect 4896 44353 4905 44387
rect 4905 44353 4939 44387
rect 4939 44353 4948 44387
rect 4896 44344 4948 44353
rect 5356 44344 5408 44396
rect 10048 44344 10100 44396
rect 29736 44344 29788 44396
rect 47768 44387 47820 44396
rect 47768 44353 47777 44387
rect 47777 44353 47811 44387
rect 47811 44353 47820 44387
rect 47768 44344 47820 44353
rect 2320 44276 2372 44328
rect 2780 44319 2832 44328
rect 2780 44285 2789 44319
rect 2789 44285 2823 44319
rect 2823 44285 2832 44319
rect 2780 44276 2832 44285
rect 4804 44276 4856 44328
rect 40040 44276 40092 44328
rect 3056 44208 3108 44260
rect 20536 44140 20588 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 3884 43936 3936 43988
rect 6552 43936 6604 43988
rect 15200 43936 15252 43988
rect 29736 43911 29788 43920
rect 29736 43877 29745 43911
rect 29745 43877 29779 43911
rect 29779 43877 29788 43911
rect 29736 43868 29788 43877
rect 2780 43843 2832 43852
rect 2780 43809 2789 43843
rect 2789 43809 2823 43843
rect 2823 43809 2832 43843
rect 2780 43800 2832 43809
rect 4988 43843 5040 43852
rect 4988 43809 4997 43843
rect 4997 43809 5031 43843
rect 5031 43809 5040 43843
rect 4988 43800 5040 43809
rect 20536 43843 20588 43852
rect 20536 43809 20545 43843
rect 20545 43809 20579 43843
rect 20579 43809 20588 43843
rect 20536 43800 20588 43809
rect 27068 43800 27120 43852
rect 29828 43800 29880 43852
rect 36544 43800 36596 43852
rect 1584 43775 1636 43784
rect 1584 43741 1593 43775
rect 1593 43741 1627 43775
rect 1627 43741 1636 43775
rect 1584 43732 1636 43741
rect 3700 43732 3752 43784
rect 4896 43732 4948 43784
rect 20352 43775 20404 43784
rect 20352 43741 20361 43775
rect 20361 43741 20395 43775
rect 20395 43741 20404 43775
rect 20352 43732 20404 43741
rect 30104 43732 30156 43784
rect 30472 43775 30524 43784
rect 30472 43741 30481 43775
rect 30481 43741 30515 43775
rect 30515 43741 30524 43775
rect 30472 43732 30524 43741
rect 30656 43775 30708 43784
rect 30656 43741 30665 43775
rect 30665 43741 30699 43775
rect 30699 43741 30708 43775
rect 30656 43732 30708 43741
rect 2412 43664 2464 43716
rect 29828 43664 29880 43716
rect 31116 43596 31168 43648
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 2412 43435 2464 43444
rect 2412 43401 2421 43435
rect 2421 43401 2455 43435
rect 2455 43401 2464 43435
rect 2412 43392 2464 43401
rect 4712 43324 4764 43376
rect 19064 43367 19116 43376
rect 19064 43333 19073 43367
rect 19073 43333 19107 43367
rect 19107 43333 19116 43367
rect 19064 43324 19116 43333
rect 27160 43324 27212 43376
rect 30656 43392 30708 43444
rect 32312 43392 32364 43444
rect 30472 43324 30524 43376
rect 31484 43324 31536 43376
rect 1584 43256 1636 43308
rect 2688 43256 2740 43308
rect 3700 43299 3752 43308
rect 3700 43265 3709 43299
rect 3709 43265 3743 43299
rect 3743 43265 3752 43299
rect 3700 43256 3752 43265
rect 25504 43299 25556 43308
rect 25504 43265 25513 43299
rect 25513 43265 25547 43299
rect 25547 43265 25556 43299
rect 25504 43256 25556 43265
rect 3148 43188 3200 43240
rect 3884 43231 3936 43240
rect 3884 43197 3893 43231
rect 3893 43197 3927 43231
rect 3927 43197 3936 43231
rect 3884 43188 3936 43197
rect 17132 43188 17184 43240
rect 17408 43231 17460 43240
rect 17408 43197 17417 43231
rect 17417 43197 17451 43231
rect 17451 43197 17460 43231
rect 17408 43188 17460 43197
rect 26240 43256 26292 43308
rect 29000 43299 29052 43308
rect 29000 43265 29009 43299
rect 29009 43265 29043 43299
rect 29043 43265 29052 43299
rect 29000 43256 29052 43265
rect 29920 43256 29972 43308
rect 30104 43299 30156 43308
rect 30104 43265 30113 43299
rect 30113 43265 30147 43299
rect 30147 43265 30156 43299
rect 30104 43256 30156 43265
rect 30564 43256 30616 43308
rect 30656 43256 30708 43308
rect 31024 43256 31076 43308
rect 31944 43256 31996 43308
rect 32496 43299 32548 43308
rect 32496 43265 32505 43299
rect 32505 43265 32539 43299
rect 32539 43265 32548 43299
rect 32496 43256 32548 43265
rect 33692 43299 33744 43308
rect 33692 43265 33701 43299
rect 33701 43265 33735 43299
rect 33735 43265 33744 43299
rect 33692 43256 33744 43265
rect 34520 43299 34572 43308
rect 34520 43265 34529 43299
rect 34529 43265 34563 43299
rect 34563 43265 34572 43299
rect 34520 43256 34572 43265
rect 36544 43256 36596 43308
rect 47400 43256 47452 43308
rect 26148 43188 26200 43240
rect 29092 43231 29144 43240
rect 29092 43197 29101 43231
rect 29101 43197 29135 43231
rect 29135 43197 29144 43231
rect 29092 43188 29144 43197
rect 29920 43120 29972 43172
rect 30288 43231 30340 43240
rect 30288 43197 30297 43231
rect 30297 43197 30331 43231
rect 30331 43197 30340 43231
rect 30288 43188 30340 43197
rect 31116 43120 31168 43172
rect 33324 43188 33376 43240
rect 34796 43231 34848 43240
rect 34796 43197 34805 43231
rect 34805 43197 34839 43231
rect 34839 43197 34848 43231
rect 34796 43188 34848 43197
rect 33508 43120 33560 43172
rect 35440 43120 35492 43172
rect 26056 43095 26108 43104
rect 26056 43061 26065 43095
rect 26065 43061 26099 43095
rect 26099 43061 26108 43095
rect 26056 43052 26108 43061
rect 30012 43052 30064 43104
rect 31300 43095 31352 43104
rect 31300 43061 31309 43095
rect 31309 43061 31343 43095
rect 31343 43061 31352 43095
rect 31300 43052 31352 43061
rect 32772 43095 32824 43104
rect 32772 43061 32781 43095
rect 32781 43061 32815 43095
rect 32815 43061 32824 43095
rect 32772 43052 32824 43061
rect 34704 43095 34756 43104
rect 34704 43061 34713 43095
rect 34713 43061 34747 43095
rect 34747 43061 34756 43095
rect 47216 43095 47268 43104
rect 34704 43052 34756 43061
rect 47216 43061 47225 43095
rect 47225 43061 47259 43095
rect 47259 43061 47268 43095
rect 47216 43052 47268 43061
rect 47860 43095 47912 43104
rect 47860 43061 47869 43095
rect 47869 43061 47903 43095
rect 47903 43061 47912 43095
rect 47860 43052 47912 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 17408 42891 17460 42900
rect 17408 42857 17417 42891
rect 17417 42857 17451 42891
rect 17451 42857 17460 42891
rect 17408 42848 17460 42857
rect 27160 42891 27212 42900
rect 27160 42857 27169 42891
rect 27169 42857 27203 42891
rect 27203 42857 27212 42891
rect 27160 42848 27212 42857
rect 29920 42848 29972 42900
rect 2320 42755 2372 42764
rect 2320 42721 2329 42755
rect 2329 42721 2363 42755
rect 2363 42721 2372 42755
rect 2320 42712 2372 42721
rect 3056 42755 3108 42764
rect 3056 42721 3065 42755
rect 3065 42721 3099 42755
rect 3099 42721 3108 42755
rect 3056 42712 3108 42721
rect 5540 42755 5592 42764
rect 5540 42721 5549 42755
rect 5549 42721 5583 42755
rect 5583 42721 5592 42755
rect 5540 42712 5592 42721
rect 29092 42780 29144 42832
rect 22560 42712 22612 42764
rect 2412 42644 2464 42696
rect 4620 42644 4672 42696
rect 2872 42576 2924 42628
rect 2136 42508 2188 42560
rect 14004 42644 14056 42696
rect 19524 42644 19576 42696
rect 20628 42644 20680 42696
rect 22836 42687 22888 42696
rect 22836 42653 22845 42687
rect 22845 42653 22879 42687
rect 22879 42653 22888 42687
rect 22836 42644 22888 42653
rect 23112 42687 23164 42696
rect 23112 42653 23147 42687
rect 23147 42653 23164 42687
rect 23112 42644 23164 42653
rect 27528 42712 27580 42764
rect 29736 42712 29788 42764
rect 30288 42712 30340 42764
rect 27068 42687 27120 42696
rect 27068 42653 27077 42687
rect 27077 42653 27111 42687
rect 27111 42653 27120 42687
rect 27252 42687 27304 42696
rect 27068 42644 27120 42653
rect 27252 42653 27261 42687
rect 27261 42653 27295 42687
rect 27295 42653 27304 42687
rect 27252 42644 27304 42653
rect 30012 42687 30064 42696
rect 30012 42653 30021 42687
rect 30021 42653 30055 42687
rect 30055 42653 30064 42687
rect 30012 42644 30064 42653
rect 5080 42619 5132 42628
rect 5080 42585 5089 42619
rect 5089 42585 5123 42619
rect 5123 42585 5132 42619
rect 5080 42576 5132 42585
rect 20352 42576 20404 42628
rect 15200 42508 15252 42560
rect 16120 42508 16172 42560
rect 19340 42508 19392 42560
rect 20168 42508 20220 42560
rect 23020 42619 23072 42628
rect 23020 42585 23029 42619
rect 23029 42585 23063 42619
rect 23063 42585 23072 42619
rect 23020 42576 23072 42585
rect 26056 42576 26108 42628
rect 24308 42508 24360 42560
rect 26148 42508 26200 42560
rect 30196 42576 30248 42628
rect 30564 42576 30616 42628
rect 32772 42712 32824 42764
rect 34520 42848 34572 42900
rect 35348 42848 35400 42900
rect 33324 42780 33376 42832
rect 31484 42687 31536 42696
rect 31484 42653 31493 42687
rect 31493 42653 31527 42687
rect 31527 42653 31536 42687
rect 31484 42644 31536 42653
rect 31944 42687 31996 42696
rect 31944 42653 31953 42687
rect 31953 42653 31987 42687
rect 31987 42653 31996 42687
rect 31944 42644 31996 42653
rect 32312 42687 32364 42696
rect 32312 42653 32321 42687
rect 32321 42653 32355 42687
rect 32355 42653 32364 42687
rect 32312 42644 32364 42653
rect 31208 42619 31260 42628
rect 31208 42585 31217 42619
rect 31217 42585 31251 42619
rect 31251 42585 31260 42619
rect 31208 42576 31260 42585
rect 31392 42576 31444 42628
rect 33416 42644 33468 42696
rect 34244 42712 34296 42764
rect 47216 42712 47268 42764
rect 48228 42755 48280 42764
rect 48228 42721 48237 42755
rect 48237 42721 48271 42755
rect 48271 42721 48280 42755
rect 48228 42712 48280 42721
rect 32496 42576 32548 42628
rect 30840 42551 30892 42560
rect 30840 42517 30849 42551
rect 30849 42517 30883 42551
rect 30883 42517 30892 42551
rect 30840 42508 30892 42517
rect 32680 42508 32732 42560
rect 34796 42644 34848 42696
rect 34428 42576 34480 42628
rect 47860 42576 47912 42628
rect 35072 42508 35124 42560
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 5080 42347 5132 42356
rect 5080 42313 5089 42347
rect 5089 42313 5123 42347
rect 5123 42313 5132 42347
rect 5080 42304 5132 42313
rect 16120 42304 16172 42356
rect 4988 42211 5040 42220
rect 4988 42177 4997 42211
rect 4997 42177 5031 42211
rect 5031 42177 5040 42211
rect 14004 42236 14056 42288
rect 4988 42168 5040 42177
rect 17132 42211 17184 42220
rect 16028 42143 16080 42152
rect 16028 42109 16037 42143
rect 16037 42109 16071 42143
rect 16071 42109 16080 42143
rect 16028 42100 16080 42109
rect 16120 42143 16172 42152
rect 16120 42109 16129 42143
rect 16129 42109 16163 42143
rect 16163 42109 16172 42143
rect 17132 42177 17141 42211
rect 17141 42177 17175 42211
rect 17175 42177 17184 42211
rect 17132 42168 17184 42177
rect 19432 42304 19484 42356
rect 19984 42304 20036 42356
rect 20352 42304 20404 42356
rect 22836 42304 22888 42356
rect 24308 42347 24360 42356
rect 24308 42313 24317 42347
rect 24317 42313 24351 42347
rect 24351 42313 24360 42347
rect 24308 42304 24360 42313
rect 25504 42304 25556 42356
rect 30472 42304 30524 42356
rect 32680 42347 32732 42356
rect 32680 42313 32689 42347
rect 32689 42313 32723 42347
rect 32723 42313 32732 42347
rect 32680 42304 32732 42313
rect 34428 42347 34480 42356
rect 34428 42313 34437 42347
rect 34437 42313 34471 42347
rect 34471 42313 34480 42347
rect 34428 42304 34480 42313
rect 19432 42168 19484 42220
rect 22100 42168 22152 42220
rect 16120 42100 16172 42109
rect 17684 42100 17736 42152
rect 22560 42143 22612 42152
rect 15476 42032 15528 42084
rect 22560 42109 22569 42143
rect 22569 42109 22603 42143
rect 22603 42109 22612 42143
rect 22560 42100 22612 42109
rect 14924 41964 14976 42016
rect 20628 42032 20680 42084
rect 23664 42211 23716 42220
rect 23664 42177 23673 42211
rect 23673 42177 23707 42211
rect 23707 42177 23716 42211
rect 23664 42168 23716 42177
rect 24216 42211 24268 42220
rect 24216 42177 24225 42211
rect 24225 42177 24259 42211
rect 24259 42177 24268 42211
rect 24216 42168 24268 42177
rect 24676 42168 24728 42220
rect 29000 42236 29052 42288
rect 30840 42236 30892 42288
rect 31944 42236 31996 42288
rect 34520 42236 34572 42288
rect 35532 42304 35584 42356
rect 26148 42143 26200 42152
rect 20996 41964 21048 42016
rect 23204 41964 23256 42016
rect 23480 42032 23532 42084
rect 26148 42109 26157 42143
rect 26157 42109 26191 42143
rect 26191 42109 26200 42143
rect 26148 42100 26200 42109
rect 27252 42168 27304 42220
rect 27528 42168 27580 42220
rect 31116 42211 31168 42220
rect 31116 42177 31125 42211
rect 31125 42177 31159 42211
rect 31159 42177 31168 42211
rect 31116 42168 31168 42177
rect 31300 42211 31352 42220
rect 31300 42177 31309 42211
rect 31309 42177 31343 42211
rect 31343 42177 31352 42211
rect 31300 42168 31352 42177
rect 31208 42100 31260 42152
rect 32128 42168 32180 42220
rect 32496 42211 32548 42220
rect 32496 42177 32505 42211
rect 32505 42177 32539 42211
rect 32539 42177 32548 42211
rect 32496 42168 32548 42177
rect 32680 42168 32732 42220
rect 33324 42168 33376 42220
rect 33416 42168 33468 42220
rect 34612 42211 34664 42220
rect 30380 42032 30432 42084
rect 31392 42032 31444 42084
rect 24216 41964 24268 42016
rect 27068 41964 27120 42016
rect 27160 41964 27212 42016
rect 31024 41964 31076 42016
rect 33692 42100 33744 42152
rect 34612 42177 34621 42211
rect 34621 42177 34655 42211
rect 34655 42177 34664 42211
rect 34612 42168 34664 42177
rect 34428 42100 34480 42152
rect 34520 42032 34572 42084
rect 34612 42032 34664 42084
rect 35072 42211 35124 42220
rect 35072 42177 35081 42211
rect 35081 42177 35115 42211
rect 35115 42177 35124 42211
rect 35072 42168 35124 42177
rect 35348 42168 35400 42220
rect 35716 42211 35768 42220
rect 35716 42177 35725 42211
rect 35725 42177 35759 42211
rect 35759 42177 35768 42211
rect 35716 42168 35768 42177
rect 47768 42211 47820 42220
rect 47768 42177 47777 42211
rect 47777 42177 47811 42211
rect 47811 42177 47820 42211
rect 47768 42168 47820 42177
rect 32036 41964 32088 42016
rect 32680 41964 32732 42016
rect 32864 42007 32916 42016
rect 32864 41973 32873 42007
rect 32873 41973 32907 42007
rect 32907 41973 32916 42007
rect 32864 41964 32916 41973
rect 34152 41964 34204 42016
rect 46480 41964 46532 42016
rect 47860 42007 47912 42016
rect 47860 41973 47869 42007
rect 47869 41973 47903 42007
rect 47903 41973 47912 42007
rect 47860 41964 47912 41973
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 17132 41760 17184 41812
rect 17500 41803 17552 41812
rect 17500 41769 17509 41803
rect 17509 41769 17543 41803
rect 17543 41769 17552 41803
rect 17500 41760 17552 41769
rect 17684 41803 17736 41812
rect 17684 41769 17693 41803
rect 17693 41769 17727 41803
rect 17727 41769 17736 41803
rect 17684 41760 17736 41769
rect 19432 41803 19484 41812
rect 19432 41769 19441 41803
rect 19441 41769 19475 41803
rect 19475 41769 19484 41803
rect 19432 41760 19484 41769
rect 22560 41760 22612 41812
rect 23204 41760 23256 41812
rect 30104 41760 30156 41812
rect 30288 41760 30340 41812
rect 31484 41760 31536 41812
rect 32312 41760 32364 41812
rect 34060 41760 34112 41812
rect 35440 41760 35492 41812
rect 17408 41692 17460 41744
rect 20168 41692 20220 41744
rect 15476 41667 15528 41676
rect 15476 41633 15485 41667
rect 15485 41633 15519 41667
rect 15519 41633 15528 41667
rect 15476 41624 15528 41633
rect 19340 41624 19392 41676
rect 20076 41667 20128 41676
rect 20076 41633 20085 41667
rect 20085 41633 20119 41667
rect 20119 41633 20128 41667
rect 20076 41624 20128 41633
rect 20352 41624 20404 41676
rect 20996 41667 21048 41676
rect 20996 41633 21005 41667
rect 21005 41633 21039 41667
rect 21039 41633 21048 41667
rect 20996 41624 21048 41633
rect 22100 41667 22152 41676
rect 22100 41633 22109 41667
rect 22109 41633 22143 41667
rect 22143 41633 22152 41667
rect 22100 41624 22152 41633
rect 2044 41556 2096 41608
rect 14924 41599 14976 41608
rect 14924 41565 14933 41599
rect 14933 41565 14967 41599
rect 14967 41565 14976 41599
rect 14924 41556 14976 41565
rect 15936 41488 15988 41540
rect 17132 41488 17184 41540
rect 14740 41463 14792 41472
rect 14740 41429 14749 41463
rect 14749 41429 14783 41463
rect 14783 41429 14792 41463
rect 14740 41420 14792 41429
rect 17408 41420 17460 41472
rect 19432 41420 19484 41472
rect 20260 41556 20312 41608
rect 20536 41556 20588 41608
rect 21824 41599 21876 41608
rect 21824 41565 21833 41599
rect 21833 41565 21867 41599
rect 21867 41565 21876 41599
rect 21824 41556 21876 41565
rect 23296 41556 23348 41608
rect 24124 41556 24176 41608
rect 32036 41692 32088 41744
rect 32128 41692 32180 41744
rect 34428 41692 34480 41744
rect 35532 41692 35584 41744
rect 26148 41624 26200 41676
rect 25780 41599 25832 41608
rect 25780 41565 25789 41599
rect 25789 41565 25823 41599
rect 25823 41565 25832 41599
rect 25780 41556 25832 41565
rect 29460 41624 29512 41676
rect 24216 41488 24268 41540
rect 24768 41531 24820 41540
rect 24768 41497 24777 41531
rect 24777 41497 24811 41531
rect 24811 41497 24820 41531
rect 24768 41488 24820 41497
rect 25964 41531 26016 41540
rect 25964 41497 25973 41531
rect 25973 41497 26007 41531
rect 26007 41497 26016 41531
rect 26976 41556 27028 41608
rect 27160 41599 27212 41608
rect 27160 41565 27169 41599
rect 27169 41565 27203 41599
rect 27203 41565 27212 41599
rect 27160 41556 27212 41565
rect 30748 41556 30800 41608
rect 31024 41599 31076 41608
rect 31024 41565 31033 41599
rect 31033 41565 31067 41599
rect 31067 41565 31076 41599
rect 31024 41556 31076 41565
rect 33416 41624 33468 41676
rect 32496 41556 32548 41608
rect 35716 41624 35768 41676
rect 46480 41667 46532 41676
rect 46480 41633 46489 41667
rect 46489 41633 46523 41667
rect 46523 41633 46532 41667
rect 46480 41624 46532 41633
rect 47860 41624 47912 41676
rect 48228 41667 48280 41676
rect 48228 41633 48237 41667
rect 48237 41633 48271 41667
rect 48271 41633 48280 41667
rect 48228 41624 48280 41633
rect 25964 41488 26016 41497
rect 27804 41488 27856 41540
rect 24308 41420 24360 41472
rect 30932 41420 30984 41472
rect 33784 41599 33836 41608
rect 33784 41565 33793 41599
rect 33793 41565 33827 41599
rect 33827 41565 33836 41599
rect 33784 41556 33836 41565
rect 34704 41556 34756 41608
rect 35348 41556 35400 41608
rect 46020 41599 46072 41608
rect 46020 41565 46029 41599
rect 46029 41565 46063 41599
rect 46063 41565 46072 41599
rect 46020 41556 46072 41565
rect 34060 41488 34112 41540
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 15200 41216 15252 41268
rect 20168 41216 20220 41268
rect 23296 41216 23348 41268
rect 24308 41216 24360 41268
rect 27068 41216 27120 41268
rect 30104 41216 30156 41268
rect 31208 41216 31260 41268
rect 14740 41148 14792 41200
rect 20076 41148 20128 41200
rect 2044 41123 2096 41132
rect 2044 41089 2053 41123
rect 2053 41089 2087 41123
rect 2087 41089 2096 41123
rect 2044 41080 2096 41089
rect 16028 41123 16080 41132
rect 16028 41089 16037 41123
rect 16037 41089 16071 41123
rect 16071 41089 16080 41123
rect 16028 41080 16080 41089
rect 17040 41123 17092 41132
rect 17040 41089 17049 41123
rect 17049 41089 17083 41123
rect 17083 41089 17092 41123
rect 17040 41080 17092 41089
rect 2320 41012 2372 41064
rect 2780 41055 2832 41064
rect 2780 41021 2789 41055
rect 2789 41021 2823 41055
rect 2823 41021 2832 41055
rect 2780 41012 2832 41021
rect 14096 41055 14148 41064
rect 14096 41021 14105 41055
rect 14105 41021 14139 41055
rect 14139 41021 14148 41055
rect 14096 41012 14148 41021
rect 17316 41123 17368 41132
rect 17316 41089 17325 41123
rect 17325 41089 17359 41123
rect 17359 41089 17368 41123
rect 17316 41080 17368 41089
rect 17500 41012 17552 41064
rect 19248 41012 19300 41064
rect 19984 41080 20036 41132
rect 20536 41148 20588 41200
rect 21824 41148 21876 41200
rect 23480 41148 23532 41200
rect 24124 41191 24176 41200
rect 20352 41123 20404 41132
rect 20352 41089 20361 41123
rect 20361 41089 20395 41123
rect 20395 41089 20404 41123
rect 20352 41080 20404 41089
rect 22100 41080 22152 41132
rect 22836 41080 22888 41132
rect 22928 41080 22980 41132
rect 24124 41157 24133 41191
rect 24133 41157 24167 41191
rect 24167 41157 24176 41191
rect 24124 41148 24176 41157
rect 25780 41148 25832 41200
rect 24308 41123 24360 41132
rect 24308 41089 24317 41123
rect 24317 41089 24351 41123
rect 24351 41089 24360 41123
rect 24308 41080 24360 41089
rect 23756 41012 23808 41064
rect 24768 41080 24820 41132
rect 26976 41080 27028 41132
rect 30932 41080 30984 41132
rect 26792 41012 26844 41064
rect 16120 40876 16172 40928
rect 20076 40876 20128 40928
rect 20444 40919 20496 40928
rect 20444 40885 20453 40919
rect 20453 40885 20487 40919
rect 20487 40885 20496 40919
rect 20444 40876 20496 40885
rect 22744 40919 22796 40928
rect 22744 40885 22753 40919
rect 22753 40885 22787 40919
rect 22787 40885 22796 40919
rect 22744 40876 22796 40885
rect 25688 40944 25740 40996
rect 25964 40944 26016 40996
rect 28448 41012 28500 41064
rect 33048 41055 33100 41064
rect 33048 41021 33057 41055
rect 33057 41021 33091 41055
rect 33091 41021 33100 41055
rect 33048 41012 33100 41021
rect 33876 41080 33928 41132
rect 34060 41055 34112 41064
rect 34060 41021 34069 41055
rect 34069 41021 34103 41055
rect 34103 41021 34112 41055
rect 34060 41012 34112 41021
rect 34612 41080 34664 41132
rect 46020 41148 46072 41200
rect 34152 40944 34204 40996
rect 24676 40876 24728 40928
rect 29460 40919 29512 40928
rect 29460 40885 29469 40919
rect 29469 40885 29503 40919
rect 29503 40885 29512 40919
rect 29460 40876 29512 40885
rect 30196 40876 30248 40928
rect 34336 40876 34388 40928
rect 34520 41055 34572 41064
rect 34520 41021 34529 41055
rect 34529 41021 34563 41055
rect 34563 41021 34572 41055
rect 34520 41012 34572 41021
rect 34796 41012 34848 41064
rect 45928 41012 45980 41064
rect 46940 41055 46992 41064
rect 46940 41021 46949 41055
rect 46949 41021 46983 41055
rect 46983 41021 46992 41055
rect 46940 41012 46992 41021
rect 46480 40876 46532 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 2320 40715 2372 40724
rect 2320 40681 2329 40715
rect 2329 40681 2363 40715
rect 2363 40681 2372 40715
rect 2320 40672 2372 40681
rect 15936 40715 15988 40724
rect 15936 40681 15945 40715
rect 15945 40681 15979 40715
rect 15979 40681 15988 40715
rect 15936 40672 15988 40681
rect 16028 40672 16080 40724
rect 21824 40672 21876 40724
rect 22928 40672 22980 40724
rect 23020 40672 23072 40724
rect 23204 40672 23256 40724
rect 23756 40672 23808 40724
rect 16948 40536 17000 40588
rect 2596 40468 2648 40520
rect 16120 40511 16172 40520
rect 16120 40477 16129 40511
rect 16129 40477 16163 40511
rect 16163 40477 16172 40511
rect 16120 40468 16172 40477
rect 17316 40536 17368 40588
rect 20076 40579 20128 40588
rect 20076 40545 20085 40579
rect 20085 40545 20119 40579
rect 20119 40545 20128 40579
rect 20076 40536 20128 40545
rect 17040 40400 17092 40452
rect 19432 40468 19484 40520
rect 20444 40468 20496 40520
rect 20628 40511 20680 40520
rect 20628 40477 20637 40511
rect 20637 40477 20671 40511
rect 20671 40477 20680 40511
rect 20628 40468 20680 40477
rect 23112 40604 23164 40656
rect 30288 40672 30340 40724
rect 33876 40715 33928 40724
rect 33876 40681 33885 40715
rect 33885 40681 33919 40715
rect 33919 40681 33928 40715
rect 33876 40672 33928 40681
rect 45928 40715 45980 40724
rect 45928 40681 45937 40715
rect 45937 40681 45971 40715
rect 45971 40681 45980 40715
rect 45928 40672 45980 40681
rect 30472 40604 30524 40656
rect 34152 40604 34204 40656
rect 22744 40536 22796 40588
rect 25780 40579 25832 40588
rect 22928 40511 22980 40520
rect 22928 40477 22963 40511
rect 22963 40477 22980 40511
rect 23112 40511 23164 40520
rect 22928 40468 22980 40477
rect 23112 40477 23121 40511
rect 23121 40477 23155 40511
rect 23155 40477 23164 40511
rect 23112 40468 23164 40477
rect 23664 40468 23716 40520
rect 25780 40545 25789 40579
rect 25789 40545 25823 40579
rect 25823 40545 25832 40579
rect 25780 40536 25832 40545
rect 26976 40536 27028 40588
rect 24676 40511 24728 40520
rect 24676 40477 24685 40511
rect 24685 40477 24719 40511
rect 24719 40477 24728 40511
rect 24676 40468 24728 40477
rect 25688 40511 25740 40520
rect 25688 40477 25697 40511
rect 25697 40477 25731 40511
rect 25731 40477 25740 40511
rect 25688 40468 25740 40477
rect 26516 40511 26568 40520
rect 26516 40477 26525 40511
rect 26525 40477 26559 40511
rect 26559 40477 26568 40511
rect 26516 40468 26568 40477
rect 26792 40468 26844 40520
rect 27068 40468 27120 40520
rect 30932 40511 30984 40520
rect 30932 40477 30941 40511
rect 30941 40477 30975 40511
rect 30975 40477 30984 40511
rect 30932 40468 30984 40477
rect 32864 40536 32916 40588
rect 34428 40536 34480 40588
rect 46480 40579 46532 40588
rect 46480 40545 46489 40579
rect 46489 40545 46523 40579
rect 46523 40545 46532 40579
rect 46480 40536 46532 40545
rect 32772 40468 32824 40520
rect 33048 40468 33100 40520
rect 20536 40400 20588 40452
rect 19432 40375 19484 40384
rect 19432 40341 19441 40375
rect 19441 40341 19475 40375
rect 19475 40341 19484 40375
rect 19432 40332 19484 40341
rect 19984 40332 20036 40384
rect 23204 40400 23256 40452
rect 26884 40400 26936 40452
rect 23480 40332 23532 40384
rect 26516 40332 26568 40384
rect 26700 40375 26752 40384
rect 26700 40341 26709 40375
rect 26709 40341 26743 40375
rect 26743 40341 26752 40375
rect 26700 40332 26752 40341
rect 27528 40400 27580 40452
rect 28448 40400 28500 40452
rect 34244 40400 34296 40452
rect 27712 40332 27764 40384
rect 28540 40375 28592 40384
rect 28540 40341 28549 40375
rect 28549 40341 28583 40375
rect 28583 40341 28592 40375
rect 28540 40332 28592 40341
rect 31116 40375 31168 40384
rect 31116 40341 31125 40375
rect 31125 40341 31159 40375
rect 31159 40341 31168 40375
rect 31116 40332 31168 40341
rect 32312 40375 32364 40384
rect 32312 40341 32321 40375
rect 32321 40341 32355 40375
rect 32355 40341 32364 40375
rect 32312 40332 32364 40341
rect 47124 40400 47176 40452
rect 48320 40443 48372 40452
rect 48320 40409 48329 40443
rect 48329 40409 48363 40443
rect 48363 40409 48372 40443
rect 48320 40400 48372 40409
rect 47032 40332 47084 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 20352 40128 20404 40180
rect 25780 40128 25832 40180
rect 27712 40171 27764 40180
rect 21824 40060 21876 40112
rect 19432 39992 19484 40044
rect 23112 40060 23164 40112
rect 22836 39992 22888 40044
rect 25688 40060 25740 40112
rect 26700 40060 26752 40112
rect 27712 40137 27721 40171
rect 27721 40137 27755 40171
rect 27755 40137 27764 40171
rect 27712 40128 27764 40137
rect 27804 40128 27856 40180
rect 28540 40060 28592 40112
rect 30472 40103 30524 40112
rect 27160 40035 27212 40044
rect 27160 40001 27169 40035
rect 27169 40001 27203 40035
rect 27203 40001 27212 40035
rect 27160 39992 27212 40001
rect 27528 40035 27580 40044
rect 27528 40001 27537 40035
rect 27537 40001 27571 40035
rect 27571 40001 27580 40035
rect 27528 39992 27580 40001
rect 30472 40069 30481 40103
rect 30481 40069 30515 40103
rect 30515 40069 30524 40103
rect 30472 40060 30524 40069
rect 32312 40060 32364 40112
rect 32864 40060 32916 40112
rect 18420 39967 18472 39976
rect 18420 39933 18429 39967
rect 18429 39933 18463 39967
rect 18463 39933 18472 39967
rect 18420 39924 18472 39933
rect 23664 39924 23716 39976
rect 26240 39924 26292 39976
rect 30196 39924 30248 39976
rect 30932 39992 30984 40044
rect 32680 40035 32732 40044
rect 32680 40001 32689 40035
rect 32689 40001 32723 40035
rect 32723 40001 32732 40035
rect 32680 39992 32732 40001
rect 47032 40035 47084 40044
rect 47032 40001 47041 40035
rect 47041 40001 47075 40035
rect 47075 40001 47084 40035
rect 47032 39992 47084 40001
rect 47124 40035 47176 40044
rect 47124 40001 47133 40035
rect 47133 40001 47167 40035
rect 47167 40001 47176 40035
rect 47124 39992 47176 40001
rect 30748 39924 30800 39976
rect 31024 39924 31076 39976
rect 25596 39856 25648 39908
rect 31116 39856 31168 39908
rect 33048 39924 33100 39976
rect 47492 39924 47544 39976
rect 28448 39788 28500 39840
rect 30380 39788 30432 39840
rect 46480 39788 46532 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 27160 39584 27212 39636
rect 30472 39584 30524 39636
rect 26516 39516 26568 39568
rect 14096 39448 14148 39500
rect 14280 39491 14332 39500
rect 14280 39457 14289 39491
rect 14289 39457 14323 39491
rect 14323 39457 14332 39491
rect 14280 39448 14332 39457
rect 18420 39448 18472 39500
rect 20628 39448 20680 39500
rect 26792 39448 26844 39500
rect 29460 39448 29512 39500
rect 26884 39423 26936 39432
rect 26884 39389 26893 39423
rect 26893 39389 26927 39423
rect 26927 39389 26936 39423
rect 27804 39423 27856 39432
rect 26884 39380 26936 39389
rect 13912 39312 13964 39364
rect 19432 39355 19484 39364
rect 19432 39321 19441 39355
rect 19441 39321 19475 39355
rect 19475 39321 19484 39355
rect 19432 39312 19484 39321
rect 15200 39244 15252 39296
rect 27804 39389 27813 39423
rect 27813 39389 27847 39423
rect 27847 39389 27856 39423
rect 27804 39380 27856 39389
rect 30472 39380 30524 39432
rect 30656 39423 30708 39432
rect 30656 39389 30665 39423
rect 30665 39389 30699 39423
rect 30699 39389 30708 39423
rect 30656 39380 30708 39389
rect 30932 39423 30984 39432
rect 30932 39389 30941 39423
rect 30941 39389 30975 39423
rect 30975 39389 30984 39423
rect 30932 39380 30984 39389
rect 34060 39516 34112 39568
rect 34152 39448 34204 39500
rect 46480 39491 46532 39500
rect 46480 39457 46489 39491
rect 46489 39457 46523 39491
rect 46523 39457 46532 39491
rect 46480 39448 46532 39457
rect 48228 39491 48280 39500
rect 48228 39457 48237 39491
rect 48237 39457 48271 39491
rect 48271 39457 48280 39491
rect 48228 39448 48280 39457
rect 32036 39423 32088 39432
rect 30564 39312 30616 39364
rect 32036 39389 32045 39423
rect 32045 39389 32079 39423
rect 32079 39389 32088 39423
rect 32036 39380 32088 39389
rect 31668 39312 31720 39364
rect 30104 39244 30156 39296
rect 30472 39287 30524 39296
rect 30472 39253 30481 39287
rect 30481 39253 30515 39287
rect 30515 39253 30524 39287
rect 30472 39244 30524 39253
rect 31484 39287 31536 39296
rect 31484 39253 31493 39287
rect 31493 39253 31527 39287
rect 31527 39253 31536 39287
rect 31484 39244 31536 39253
rect 31576 39244 31628 39296
rect 47860 39312 47912 39364
rect 32404 39287 32456 39296
rect 32404 39253 32413 39287
rect 32413 39253 32447 39287
rect 32447 39253 32456 39287
rect 32404 39244 32456 39253
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 13912 39083 13964 39092
rect 13912 39049 13921 39083
rect 13921 39049 13955 39083
rect 13955 39049 13964 39083
rect 13912 39040 13964 39049
rect 19984 39040 20036 39092
rect 21088 39040 21140 39092
rect 22376 39040 22428 39092
rect 30564 39040 30616 39092
rect 31024 39083 31076 39092
rect 31024 39049 31033 39083
rect 31033 39049 31067 39083
rect 31067 39049 31076 39083
rect 31024 39040 31076 39049
rect 1584 38947 1636 38956
rect 1584 38913 1593 38947
rect 1593 38913 1627 38947
rect 1627 38913 1636 38947
rect 1584 38904 1636 38913
rect 14096 38947 14148 38956
rect 14096 38913 14105 38947
rect 14105 38913 14139 38947
rect 14139 38913 14148 38947
rect 14096 38904 14148 38913
rect 14280 38904 14332 38956
rect 15476 38904 15528 38956
rect 18420 38972 18472 39024
rect 25412 38972 25464 39024
rect 17500 38947 17552 38956
rect 17500 38913 17534 38947
rect 17534 38913 17552 38947
rect 19616 38947 19668 38956
rect 17500 38904 17552 38913
rect 19616 38913 19625 38947
rect 19625 38913 19659 38947
rect 19659 38913 19668 38947
rect 19616 38904 19668 38913
rect 19984 38904 20036 38956
rect 20536 38904 20588 38956
rect 14372 38879 14424 38888
rect 14372 38845 14381 38879
rect 14381 38845 14415 38879
rect 14415 38845 14424 38879
rect 14372 38836 14424 38845
rect 20444 38836 20496 38888
rect 22652 38904 22704 38956
rect 24216 38947 24268 38956
rect 24216 38913 24225 38947
rect 24225 38913 24259 38947
rect 24259 38913 24268 38947
rect 24216 38904 24268 38913
rect 25044 38904 25096 38956
rect 25320 38947 25372 38956
rect 25320 38913 25329 38947
rect 25329 38913 25363 38947
rect 25363 38913 25372 38947
rect 25320 38904 25372 38913
rect 23388 38836 23440 38888
rect 24952 38879 25004 38888
rect 24952 38845 24961 38879
rect 24961 38845 24995 38879
rect 24995 38845 25004 38879
rect 24952 38836 25004 38845
rect 25136 38836 25188 38888
rect 29736 38904 29788 38956
rect 30932 38947 30984 38956
rect 30932 38913 30941 38947
rect 30941 38913 30975 38947
rect 30975 38913 30984 38947
rect 30932 38904 30984 38913
rect 31576 38904 31628 38956
rect 32680 39040 32732 39092
rect 33140 39040 33192 39092
rect 47860 39083 47912 39092
rect 47860 39049 47869 39083
rect 47869 39049 47903 39083
rect 47903 39049 47912 39083
rect 47860 39040 47912 39049
rect 32864 38972 32916 39024
rect 34060 38947 34112 38956
rect 34060 38913 34069 38947
rect 34069 38913 34103 38947
rect 34103 38913 34112 38947
rect 34060 38904 34112 38913
rect 26148 38879 26200 38888
rect 26148 38845 26157 38879
rect 26157 38845 26191 38879
rect 26191 38845 26200 38879
rect 26148 38836 26200 38845
rect 27068 38836 27120 38888
rect 30472 38836 30524 38888
rect 23480 38811 23532 38820
rect 23480 38777 23489 38811
rect 23489 38777 23523 38811
rect 23523 38777 23532 38811
rect 23480 38768 23532 38777
rect 25596 38811 25648 38820
rect 25596 38777 25605 38811
rect 25605 38777 25639 38811
rect 25639 38777 25648 38811
rect 25596 38768 25648 38777
rect 1860 38700 1912 38752
rect 15568 38700 15620 38752
rect 16120 38700 16172 38752
rect 18420 38700 18472 38752
rect 22560 38743 22612 38752
rect 22560 38709 22569 38743
rect 22569 38709 22603 38743
rect 22603 38709 22612 38743
rect 22560 38700 22612 38709
rect 22744 38743 22796 38752
rect 22744 38709 22753 38743
rect 22753 38709 22787 38743
rect 22787 38709 22796 38743
rect 22744 38700 22796 38709
rect 23572 38700 23624 38752
rect 24860 38700 24912 38752
rect 35348 38947 35400 38956
rect 35348 38913 35382 38947
rect 35382 38913 35400 38947
rect 35348 38904 35400 38913
rect 47308 38904 47360 38956
rect 34796 38836 34848 38888
rect 26148 38743 26200 38752
rect 26148 38709 26157 38743
rect 26157 38709 26191 38743
rect 26191 38709 26200 38743
rect 26148 38700 26200 38709
rect 29184 38700 29236 38752
rect 32680 38743 32732 38752
rect 32680 38709 32689 38743
rect 32689 38709 32723 38743
rect 32723 38709 32732 38743
rect 32680 38700 32732 38709
rect 34152 38700 34204 38752
rect 34704 38700 34756 38752
rect 35440 38700 35492 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 14096 38496 14148 38548
rect 17132 38496 17184 38548
rect 19616 38496 19668 38548
rect 23112 38496 23164 38548
rect 24216 38496 24268 38548
rect 24860 38539 24912 38548
rect 24860 38505 24869 38539
rect 24869 38505 24903 38539
rect 24903 38505 24912 38539
rect 24860 38496 24912 38505
rect 25044 38539 25096 38548
rect 25044 38505 25053 38539
rect 25053 38505 25087 38539
rect 25087 38505 25096 38539
rect 25044 38496 25096 38505
rect 29736 38539 29788 38548
rect 29736 38505 29745 38539
rect 29745 38505 29779 38539
rect 29779 38505 29788 38539
rect 29736 38496 29788 38505
rect 32036 38496 32088 38548
rect 32772 38539 32824 38548
rect 32772 38505 32781 38539
rect 32781 38505 32815 38539
rect 32815 38505 32824 38539
rect 32772 38496 32824 38505
rect 32864 38496 32916 38548
rect 35348 38496 35400 38548
rect 22560 38428 22612 38480
rect 23848 38428 23900 38480
rect 23940 38428 23992 38480
rect 15200 38292 15252 38344
rect 16120 38335 16172 38344
rect 16120 38301 16129 38335
rect 16129 38301 16163 38335
rect 16163 38301 16172 38335
rect 16120 38292 16172 38301
rect 16856 38335 16908 38344
rect 16856 38301 16865 38335
rect 16865 38301 16899 38335
rect 16899 38301 16908 38335
rect 16856 38292 16908 38301
rect 18420 38335 18472 38344
rect 17132 38267 17184 38276
rect 15384 38156 15436 38208
rect 17132 38233 17141 38267
rect 17141 38233 17175 38267
rect 17175 38233 17184 38267
rect 17132 38224 17184 38233
rect 17592 38224 17644 38276
rect 18420 38301 18429 38335
rect 18429 38301 18463 38335
rect 18463 38301 18472 38335
rect 18420 38292 18472 38301
rect 19984 38267 20036 38276
rect 19984 38233 19993 38267
rect 19993 38233 20027 38267
rect 20027 38233 20036 38267
rect 19984 38224 20036 38233
rect 17684 38156 17736 38208
rect 19248 38156 19300 38208
rect 20628 38360 20680 38412
rect 22560 38224 22612 38276
rect 22928 38292 22980 38344
rect 23480 38292 23532 38344
rect 26148 38428 26200 38480
rect 30564 38428 30616 38480
rect 24860 38360 24912 38412
rect 21272 38156 21324 38208
rect 22468 38156 22520 38208
rect 22836 38199 22888 38208
rect 22836 38165 22861 38199
rect 22861 38165 22888 38199
rect 23572 38224 23624 38276
rect 25964 38292 26016 38344
rect 27528 38360 27580 38412
rect 28264 38335 28316 38344
rect 25504 38224 25556 38276
rect 27252 38267 27304 38276
rect 22836 38156 22888 38165
rect 24952 38156 25004 38208
rect 27252 38233 27261 38267
rect 27261 38233 27295 38267
rect 27295 38233 27304 38267
rect 27252 38224 27304 38233
rect 27712 38224 27764 38276
rect 28264 38301 28273 38335
rect 28273 38301 28307 38335
rect 28307 38301 28316 38335
rect 28264 38292 28316 38301
rect 31484 38360 31536 38412
rect 33416 38403 33468 38412
rect 33416 38369 33425 38403
rect 33425 38369 33459 38403
rect 33459 38369 33468 38403
rect 33416 38360 33468 38369
rect 30564 38292 30616 38344
rect 31208 38292 31260 38344
rect 31668 38292 31720 38344
rect 28540 38224 28592 38276
rect 27068 38156 27120 38208
rect 27620 38199 27672 38208
rect 27620 38165 27629 38199
rect 27629 38165 27663 38199
rect 27663 38165 27672 38199
rect 27620 38156 27672 38165
rect 30104 38267 30156 38276
rect 30104 38233 30113 38267
rect 30113 38233 30147 38267
rect 30147 38233 30156 38267
rect 30104 38224 30156 38233
rect 30472 38224 30524 38276
rect 30932 38224 30984 38276
rect 32312 38267 32364 38276
rect 32312 38233 32321 38267
rect 32321 38233 32355 38267
rect 32355 38233 32364 38267
rect 32312 38224 32364 38233
rect 32956 38224 33008 38276
rect 33508 38292 33560 38344
rect 34152 38471 34204 38480
rect 34152 38437 34161 38471
rect 34161 38437 34195 38471
rect 34195 38437 34204 38471
rect 34152 38428 34204 38437
rect 34244 38360 34296 38412
rect 34704 38292 34756 38344
rect 35440 38360 35492 38412
rect 47676 38335 47728 38344
rect 34428 38224 34480 38276
rect 47676 38301 47685 38335
rect 47685 38301 47719 38335
rect 47719 38301 47728 38335
rect 47676 38292 47728 38301
rect 30380 38156 30432 38208
rect 30564 38156 30616 38208
rect 31668 38156 31720 38208
rect 33048 38156 33100 38208
rect 33876 38156 33928 38208
rect 34244 38156 34296 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 15476 37952 15528 38004
rect 17500 37995 17552 38004
rect 17500 37961 17509 37995
rect 17509 37961 17543 37995
rect 17543 37961 17552 37995
rect 17500 37952 17552 37961
rect 20260 37952 20312 38004
rect 12900 37859 12952 37868
rect 12900 37825 12909 37859
rect 12909 37825 12943 37859
rect 12943 37825 12952 37859
rect 12900 37816 12952 37825
rect 15384 37859 15436 37868
rect 15384 37825 15393 37859
rect 15393 37825 15427 37859
rect 15427 37825 15436 37859
rect 15384 37816 15436 37825
rect 15568 37859 15620 37868
rect 15568 37825 15577 37859
rect 15577 37825 15611 37859
rect 15611 37825 15620 37859
rect 17684 37859 17736 37868
rect 15568 37816 15620 37825
rect 15660 37791 15712 37800
rect 15660 37757 15669 37791
rect 15669 37757 15703 37791
rect 15703 37757 15712 37791
rect 15660 37748 15712 37757
rect 17684 37825 17693 37859
rect 17693 37825 17727 37859
rect 17727 37825 17736 37859
rect 17684 37816 17736 37825
rect 17960 37859 18012 37868
rect 17960 37825 17969 37859
rect 17969 37825 18003 37859
rect 18003 37825 18012 37859
rect 17960 37816 18012 37825
rect 18696 37816 18748 37868
rect 20168 37816 20220 37868
rect 17224 37748 17276 37800
rect 20076 37791 20128 37800
rect 20076 37757 20085 37791
rect 20085 37757 20119 37791
rect 20119 37757 20128 37791
rect 20076 37748 20128 37757
rect 22744 37884 22796 37936
rect 22284 37816 22336 37868
rect 22468 37859 22520 37868
rect 22468 37825 22477 37859
rect 22477 37825 22511 37859
rect 22511 37825 22520 37859
rect 22468 37816 22520 37825
rect 24860 37952 24912 38004
rect 25320 37995 25372 38004
rect 25320 37961 25329 37995
rect 25329 37961 25363 37995
rect 25363 37961 25372 37995
rect 25320 37952 25372 37961
rect 28540 37995 28592 38004
rect 28540 37961 28549 37995
rect 28549 37961 28583 37995
rect 28583 37961 28592 37995
rect 28540 37952 28592 37961
rect 31208 37952 31260 38004
rect 32404 37952 32456 38004
rect 33048 37952 33100 38004
rect 23848 37859 23900 37868
rect 23848 37825 23857 37859
rect 23857 37825 23891 37859
rect 23891 37825 23900 37859
rect 26056 37884 26108 37936
rect 23848 37816 23900 37825
rect 25780 37859 25832 37868
rect 25780 37825 25789 37859
rect 25789 37825 25823 37859
rect 25823 37825 25832 37859
rect 25780 37816 25832 37825
rect 26148 37816 26200 37868
rect 27620 37884 27672 37936
rect 27896 37816 27948 37868
rect 30656 37884 30708 37936
rect 30564 37859 30616 37868
rect 30564 37825 30573 37859
rect 30573 37825 30607 37859
rect 30607 37825 30616 37859
rect 30564 37816 30616 37825
rect 33416 37884 33468 37936
rect 34152 37927 34204 37936
rect 34152 37893 34161 37927
rect 34161 37893 34195 37927
rect 34195 37893 34204 37927
rect 34152 37884 34204 37893
rect 32956 37859 33008 37868
rect 32956 37825 32965 37859
rect 32965 37825 32999 37859
rect 32999 37825 33008 37859
rect 33876 37859 33928 37868
rect 32956 37816 33008 37825
rect 33876 37825 33885 37859
rect 33885 37825 33919 37859
rect 33919 37825 33928 37859
rect 33876 37816 33928 37825
rect 23480 37748 23532 37800
rect 22560 37680 22612 37732
rect 23112 37680 23164 37732
rect 23940 37791 23992 37800
rect 23940 37757 23949 37791
rect 23949 37757 23983 37791
rect 23983 37757 23992 37791
rect 23940 37748 23992 37757
rect 27068 37748 27120 37800
rect 34336 37816 34388 37868
rect 47768 37859 47820 37868
rect 47768 37825 47777 37859
rect 47777 37825 47811 37859
rect 47811 37825 47820 37859
rect 47768 37816 47820 37825
rect 12624 37612 12676 37664
rect 21732 37612 21784 37664
rect 24768 37612 24820 37664
rect 26424 37655 26476 37664
rect 26424 37621 26433 37655
rect 26433 37621 26467 37655
rect 26467 37621 26476 37655
rect 26424 37612 26476 37621
rect 32956 37612 33008 37664
rect 34704 37612 34756 37664
rect 47860 37655 47912 37664
rect 47860 37621 47869 37655
rect 47869 37621 47903 37655
rect 47903 37621 47912 37655
rect 47860 37612 47912 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 16856 37408 16908 37460
rect 19984 37408 20036 37460
rect 22652 37451 22704 37460
rect 22652 37417 22661 37451
rect 22661 37417 22695 37451
rect 22695 37417 22704 37451
rect 22652 37408 22704 37417
rect 23480 37451 23532 37460
rect 22468 37340 22520 37392
rect 1584 37247 1636 37256
rect 1584 37213 1593 37247
rect 1593 37213 1627 37247
rect 1627 37213 1636 37247
rect 1584 37204 1636 37213
rect 12348 37247 12400 37256
rect 12348 37213 12357 37247
rect 12357 37213 12391 37247
rect 12391 37213 12400 37247
rect 12348 37204 12400 37213
rect 12624 37247 12676 37256
rect 12624 37213 12658 37247
rect 12658 37213 12676 37247
rect 12624 37204 12676 37213
rect 15660 37272 15712 37324
rect 12440 37136 12492 37188
rect 17868 37247 17920 37256
rect 17868 37213 17877 37247
rect 17877 37213 17911 37247
rect 17911 37213 17920 37247
rect 17868 37204 17920 37213
rect 18696 37247 18748 37256
rect 18696 37213 18705 37247
rect 18705 37213 18739 37247
rect 18739 37213 18748 37247
rect 18696 37204 18748 37213
rect 19340 37204 19392 37256
rect 20076 37204 20128 37256
rect 21272 37247 21324 37256
rect 21272 37213 21281 37247
rect 21281 37213 21315 37247
rect 21315 37213 21324 37247
rect 21272 37204 21324 37213
rect 21548 37247 21600 37256
rect 21548 37213 21557 37247
rect 21557 37213 21591 37247
rect 21591 37213 21600 37247
rect 21548 37204 21600 37213
rect 21732 37247 21784 37256
rect 21732 37213 21741 37247
rect 21741 37213 21775 37247
rect 21775 37213 21784 37247
rect 21732 37204 21784 37213
rect 23112 37204 23164 37256
rect 23480 37417 23489 37451
rect 23489 37417 23523 37451
rect 23523 37417 23532 37451
rect 23480 37408 23532 37417
rect 27252 37408 27304 37460
rect 27896 37451 27948 37460
rect 27896 37417 27905 37451
rect 27905 37417 27939 37451
rect 27939 37417 27948 37451
rect 27896 37408 27948 37417
rect 33416 37408 33468 37460
rect 25780 37272 25832 37324
rect 26424 37272 26476 37324
rect 28264 37272 28316 37324
rect 48228 37315 48280 37324
rect 48228 37281 48237 37315
rect 48237 37281 48271 37315
rect 48271 37281 48280 37315
rect 48228 37272 48280 37281
rect 23572 37247 23624 37256
rect 23572 37213 23581 37247
rect 23581 37213 23615 37247
rect 23615 37213 23624 37247
rect 23572 37204 23624 37213
rect 24768 37204 24820 37256
rect 25872 37247 25924 37256
rect 25872 37213 25881 37247
rect 25881 37213 25915 37247
rect 25915 37213 25924 37247
rect 25872 37204 25924 37213
rect 27712 37247 27764 37256
rect 19432 37179 19484 37188
rect 13636 37068 13688 37120
rect 16948 37068 17000 37120
rect 17776 37068 17828 37120
rect 19432 37145 19441 37179
rect 19441 37145 19475 37179
rect 19475 37145 19484 37179
rect 19432 37136 19484 37145
rect 22652 37179 22704 37188
rect 20352 37068 20404 37120
rect 22652 37145 22661 37179
rect 22661 37145 22695 37179
rect 22695 37145 22704 37179
rect 22652 37136 22704 37145
rect 22836 37179 22888 37188
rect 22836 37145 22845 37179
rect 22845 37145 22879 37179
rect 22879 37145 22888 37179
rect 25044 37179 25096 37188
rect 22836 37136 22888 37145
rect 25044 37145 25053 37179
rect 25053 37145 25087 37179
rect 25087 37145 25096 37179
rect 25044 37136 25096 37145
rect 27712 37213 27721 37247
rect 27721 37213 27755 37247
rect 27755 37213 27764 37247
rect 27712 37204 27764 37213
rect 31668 37204 31720 37256
rect 33876 37247 33928 37256
rect 25136 37068 25188 37120
rect 26884 37179 26936 37188
rect 26884 37145 26893 37179
rect 26893 37145 26927 37179
rect 26927 37145 26936 37179
rect 26884 37136 26936 37145
rect 33876 37213 33885 37247
rect 33885 37213 33919 37247
rect 33919 37213 33928 37247
rect 33876 37204 33928 37213
rect 34796 37204 34848 37256
rect 36636 37204 36688 37256
rect 33600 37136 33652 37188
rect 34704 37136 34756 37188
rect 33140 37068 33192 37120
rect 33416 37068 33468 37120
rect 34152 37068 34204 37120
rect 47860 37136 47912 37188
rect 47676 37068 47728 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 1768 36864 1820 36916
rect 12900 36864 12952 36916
rect 13636 36907 13688 36916
rect 13636 36873 13645 36907
rect 13645 36873 13679 36907
rect 13679 36873 13688 36907
rect 13636 36864 13688 36873
rect 16120 36864 16172 36916
rect 18328 36796 18380 36848
rect 21732 36864 21784 36916
rect 23388 36864 23440 36916
rect 26884 36864 26936 36916
rect 31668 36864 31720 36916
rect 33692 36864 33744 36916
rect 33876 36864 33928 36916
rect 20076 36796 20128 36848
rect 17132 36728 17184 36780
rect 18420 36728 18472 36780
rect 19892 36728 19944 36780
rect 19984 36728 20036 36780
rect 14096 36660 14148 36712
rect 16028 36703 16080 36712
rect 16028 36669 16037 36703
rect 16037 36669 16071 36703
rect 16071 36669 16080 36703
rect 16028 36660 16080 36669
rect 16120 36703 16172 36712
rect 16120 36669 16129 36703
rect 16129 36669 16163 36703
rect 16163 36669 16172 36703
rect 16120 36660 16172 36669
rect 19432 36524 19484 36576
rect 19708 36567 19760 36576
rect 19708 36533 19717 36567
rect 19717 36533 19751 36567
rect 19751 36533 19760 36567
rect 20628 36771 20680 36780
rect 20628 36737 20642 36771
rect 20642 36737 20676 36771
rect 20676 36737 20680 36771
rect 20628 36728 20680 36737
rect 21732 36728 21784 36780
rect 22468 36728 22520 36780
rect 23572 36796 23624 36848
rect 26424 36796 26476 36848
rect 24584 36771 24636 36780
rect 24584 36737 24593 36771
rect 24593 36737 24627 36771
rect 24627 36737 24636 36771
rect 24584 36728 24636 36737
rect 25504 36728 25556 36780
rect 25780 36728 25832 36780
rect 22008 36660 22060 36712
rect 25872 36660 25924 36712
rect 27068 36728 27120 36780
rect 28632 36728 28684 36780
rect 32312 36728 32364 36780
rect 32956 36771 33008 36780
rect 32956 36737 32965 36771
rect 32965 36737 32999 36771
rect 32999 36737 33008 36771
rect 32956 36728 33008 36737
rect 33416 36771 33468 36780
rect 33416 36737 33425 36771
rect 33425 36737 33459 36771
rect 33459 36737 33468 36771
rect 33416 36728 33468 36737
rect 33600 36771 33652 36780
rect 33600 36737 33609 36771
rect 33609 36737 33643 36771
rect 33643 36737 33652 36771
rect 33600 36728 33652 36737
rect 33324 36660 33376 36712
rect 20536 36592 20588 36644
rect 19708 36524 19760 36533
rect 21272 36524 21324 36576
rect 28724 36524 28776 36576
rect 33048 36524 33100 36576
rect 46480 36524 46532 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 16028 36320 16080 36372
rect 20168 36363 20220 36372
rect 20168 36329 20177 36363
rect 20177 36329 20211 36363
rect 20211 36329 20220 36363
rect 20168 36320 20220 36329
rect 25780 36320 25832 36372
rect 16120 36184 16172 36236
rect 16948 36184 17000 36236
rect 18328 36184 18380 36236
rect 20628 36227 20680 36236
rect 20628 36193 20637 36227
rect 20637 36193 20671 36227
rect 20671 36193 20680 36227
rect 20628 36184 20680 36193
rect 11796 36116 11848 36168
rect 12348 36159 12400 36168
rect 12348 36125 12357 36159
rect 12357 36125 12391 36159
rect 12391 36125 12400 36159
rect 12348 36116 12400 36125
rect 15200 36159 15252 36168
rect 15200 36125 15209 36159
rect 15209 36125 15243 36159
rect 15243 36125 15252 36159
rect 15200 36116 15252 36125
rect 16304 36159 16356 36168
rect 16304 36125 16313 36159
rect 16313 36125 16347 36159
rect 16347 36125 16356 36159
rect 16304 36116 16356 36125
rect 12808 36048 12860 36100
rect 20168 36116 20220 36168
rect 20352 36159 20404 36168
rect 20352 36125 20361 36159
rect 20361 36125 20395 36159
rect 20395 36125 20404 36159
rect 20352 36116 20404 36125
rect 20536 36159 20588 36168
rect 20536 36125 20545 36159
rect 20545 36125 20579 36159
rect 20579 36125 20588 36159
rect 20536 36116 20588 36125
rect 22192 36159 22244 36168
rect 22192 36125 22201 36159
rect 22201 36125 22235 36159
rect 22235 36125 22244 36159
rect 22192 36116 22244 36125
rect 22652 36116 22704 36168
rect 24768 36252 24820 36304
rect 25872 36184 25924 36236
rect 28632 36320 28684 36372
rect 32680 36320 32732 36372
rect 33324 36320 33376 36372
rect 33140 36252 33192 36304
rect 34428 36252 34480 36304
rect 25044 36116 25096 36168
rect 19708 36048 19760 36100
rect 20076 36048 20128 36100
rect 22284 36048 22336 36100
rect 22836 36048 22888 36100
rect 13820 35980 13872 36032
rect 14832 36023 14884 36032
rect 14832 35989 14841 36023
rect 14841 35989 14875 36023
rect 14875 35989 14884 36023
rect 14832 35980 14884 35989
rect 15292 36023 15344 36032
rect 15292 35989 15301 36023
rect 15301 35989 15335 36023
rect 15335 35989 15344 36023
rect 15292 35980 15344 35989
rect 19340 35980 19392 36032
rect 22744 35980 22796 36032
rect 25228 36023 25280 36032
rect 25228 35989 25237 36023
rect 25237 35989 25271 36023
rect 25271 35989 25280 36023
rect 25228 35980 25280 35989
rect 25688 36159 25740 36168
rect 25688 36125 25697 36159
rect 25697 36125 25731 36159
rect 25731 36125 25740 36159
rect 25688 36116 25740 36125
rect 26332 36116 26384 36168
rect 26424 36159 26476 36168
rect 26424 36125 26433 36159
rect 26433 36125 26467 36159
rect 26467 36125 26476 36159
rect 26884 36159 26936 36168
rect 26424 36116 26476 36125
rect 26884 36125 26893 36159
rect 26893 36125 26927 36159
rect 26927 36125 26936 36159
rect 26884 36116 26936 36125
rect 32680 36184 32732 36236
rect 46480 36227 46532 36236
rect 46480 36193 46489 36227
rect 46489 36193 46523 36227
rect 46523 36193 46532 36227
rect 46480 36184 46532 36193
rect 48228 36227 48280 36236
rect 48228 36193 48237 36227
rect 48237 36193 48271 36227
rect 48271 36193 48280 36227
rect 48228 36184 48280 36193
rect 28264 36116 28316 36168
rect 26700 36048 26752 36100
rect 27620 36048 27672 36100
rect 30288 36116 30340 36168
rect 28448 35980 28500 36032
rect 33048 36159 33100 36168
rect 33048 36125 33057 36159
rect 33057 36125 33091 36159
rect 33091 36125 33100 36159
rect 33876 36159 33928 36168
rect 33048 36116 33100 36125
rect 33876 36125 33885 36159
rect 33885 36125 33919 36159
rect 33919 36125 33928 36159
rect 33876 36116 33928 36125
rect 33140 36091 33192 36100
rect 33140 36057 33149 36091
rect 33149 36057 33183 36091
rect 33183 36057 33192 36091
rect 33140 36048 33192 36057
rect 33232 36091 33284 36100
rect 33232 36057 33267 36091
rect 33267 36057 33284 36091
rect 33232 36048 33284 36057
rect 47860 36048 47912 36100
rect 33416 35980 33468 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 12808 35819 12860 35828
rect 12808 35785 12817 35819
rect 12817 35785 12851 35819
rect 12851 35785 12860 35819
rect 12808 35776 12860 35785
rect 13820 35819 13872 35828
rect 13820 35785 13829 35819
rect 13829 35785 13863 35819
rect 13863 35785 13872 35819
rect 13820 35776 13872 35785
rect 14832 35776 14884 35828
rect 16948 35819 17000 35828
rect 16948 35785 16957 35819
rect 16957 35785 16991 35819
rect 16991 35785 17000 35819
rect 16948 35776 17000 35785
rect 19984 35776 20036 35828
rect 22192 35776 22244 35828
rect 23296 35776 23348 35828
rect 25228 35776 25280 35828
rect 26884 35776 26936 35828
rect 30104 35776 30156 35828
rect 30932 35776 30984 35828
rect 33140 35776 33192 35828
rect 33416 35819 33468 35828
rect 33416 35785 33425 35819
rect 33425 35785 33459 35819
rect 33459 35785 33468 35819
rect 33416 35776 33468 35785
rect 47860 35819 47912 35828
rect 47860 35785 47869 35819
rect 47869 35785 47903 35819
rect 47903 35785 47912 35819
rect 47860 35776 47912 35785
rect 13636 35708 13688 35760
rect 15384 35708 15436 35760
rect 13728 35640 13780 35692
rect 17684 35683 17736 35692
rect 17684 35649 17693 35683
rect 17693 35649 17727 35683
rect 17727 35649 17736 35683
rect 17684 35640 17736 35649
rect 17868 35683 17920 35692
rect 17868 35649 17877 35683
rect 17877 35649 17911 35683
rect 17911 35649 17920 35683
rect 17868 35640 17920 35649
rect 19340 35708 19392 35760
rect 26332 35708 26384 35760
rect 14096 35615 14148 35624
rect 14096 35581 14105 35615
rect 14105 35581 14139 35615
rect 14139 35581 14148 35615
rect 14096 35572 14148 35581
rect 16304 35572 16356 35624
rect 19064 35683 19116 35692
rect 19064 35649 19073 35683
rect 19073 35649 19107 35683
rect 19107 35649 19116 35683
rect 19248 35683 19300 35692
rect 19064 35640 19116 35649
rect 19248 35649 19257 35683
rect 19257 35649 19291 35683
rect 19291 35649 19300 35683
rect 19248 35640 19300 35649
rect 19616 35640 19668 35692
rect 20076 35683 20128 35692
rect 20076 35649 20085 35683
rect 20085 35649 20119 35683
rect 20119 35649 20128 35683
rect 20076 35640 20128 35649
rect 22100 35640 22152 35692
rect 26424 35640 26476 35692
rect 27436 35640 27488 35692
rect 30288 35708 30340 35760
rect 30472 35751 30524 35760
rect 30472 35717 30481 35751
rect 30481 35717 30515 35751
rect 30515 35717 30524 35751
rect 30472 35708 30524 35717
rect 32956 35708 33008 35760
rect 29000 35640 29052 35692
rect 30104 35640 30156 35692
rect 31668 35640 31720 35692
rect 33324 35683 33376 35692
rect 33324 35649 33333 35683
rect 33333 35649 33367 35683
rect 33367 35649 33376 35683
rect 33324 35640 33376 35649
rect 33692 35640 33744 35692
rect 47400 35640 47452 35692
rect 18880 35572 18932 35624
rect 20168 35572 20220 35624
rect 22008 35615 22060 35624
rect 22008 35581 22017 35615
rect 22017 35581 22051 35615
rect 22051 35581 22060 35615
rect 22008 35572 22060 35581
rect 25412 35572 25464 35624
rect 32680 35572 32732 35624
rect 33876 35572 33928 35624
rect 19800 35504 19852 35556
rect 30472 35504 30524 35556
rect 31668 35504 31720 35556
rect 33232 35504 33284 35556
rect 15660 35436 15712 35488
rect 19524 35436 19576 35488
rect 20904 35436 20956 35488
rect 22652 35436 22704 35488
rect 24584 35436 24636 35488
rect 30196 35436 30248 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 15292 35232 15344 35284
rect 16948 35232 17000 35284
rect 19616 35275 19668 35284
rect 19616 35241 19625 35275
rect 19625 35241 19659 35275
rect 19659 35241 19668 35275
rect 19616 35232 19668 35241
rect 23388 35232 23440 35284
rect 15384 35164 15436 35216
rect 17684 35164 17736 35216
rect 19064 35164 19116 35216
rect 19524 35207 19576 35216
rect 19524 35173 19533 35207
rect 19533 35173 19567 35207
rect 19567 35173 19576 35207
rect 19524 35164 19576 35173
rect 19800 35164 19852 35216
rect 26332 35232 26384 35284
rect 27896 35164 27948 35216
rect 13820 35096 13872 35148
rect 15660 35139 15712 35148
rect 15660 35105 15669 35139
rect 15669 35105 15703 35139
rect 15703 35105 15712 35139
rect 15660 35096 15712 35105
rect 13636 35028 13688 35080
rect 13728 35071 13780 35080
rect 13728 35037 13737 35071
rect 13737 35037 13771 35071
rect 13771 35037 13780 35071
rect 14556 35071 14608 35080
rect 13728 35028 13780 35037
rect 14556 35037 14565 35071
rect 14565 35037 14599 35071
rect 14599 35037 14608 35071
rect 14556 35028 14608 35037
rect 14740 35071 14792 35080
rect 14740 35037 14749 35071
rect 14749 35037 14783 35071
rect 14783 35037 14792 35071
rect 14740 35028 14792 35037
rect 15844 35028 15896 35080
rect 21640 35139 21692 35148
rect 21640 35105 21649 35139
rect 21649 35105 21683 35139
rect 21683 35105 21692 35139
rect 21640 35096 21692 35105
rect 22376 35096 22428 35148
rect 27528 35096 27580 35148
rect 18880 35028 18932 35080
rect 19340 35028 19392 35080
rect 21732 35071 21784 35080
rect 21732 35037 21746 35071
rect 21746 35037 21780 35071
rect 21780 35037 21784 35071
rect 22284 35071 22336 35080
rect 21732 35028 21784 35037
rect 22284 35037 22293 35071
rect 22293 35037 22327 35071
rect 22327 35037 22336 35071
rect 22284 35028 22336 35037
rect 22652 35028 22704 35080
rect 27068 35028 27120 35080
rect 27160 35071 27212 35080
rect 27160 35037 27169 35071
rect 27169 35037 27203 35071
rect 27203 35037 27212 35071
rect 27160 35028 27212 35037
rect 28724 35071 28776 35080
rect 20076 34960 20128 35012
rect 15016 34892 15068 34944
rect 16672 34892 16724 34944
rect 17868 34892 17920 34944
rect 21456 34960 21508 35012
rect 21916 34960 21968 35012
rect 23112 34960 23164 35012
rect 23296 35003 23348 35012
rect 23296 34969 23305 35003
rect 23305 34969 23339 35003
rect 23339 34969 23348 35003
rect 23296 34960 23348 34969
rect 24400 34960 24452 35012
rect 26424 34960 26476 35012
rect 28724 35037 28733 35071
rect 28733 35037 28767 35071
rect 28767 35037 28776 35071
rect 28724 35028 28776 35037
rect 29092 35028 29144 35080
rect 30196 35028 30248 35080
rect 30748 35071 30800 35080
rect 30748 35037 30757 35071
rect 30757 35037 30791 35071
rect 30791 35037 30800 35071
rect 30748 35028 30800 35037
rect 31024 35071 31076 35080
rect 31024 35037 31033 35071
rect 31033 35037 31067 35071
rect 31067 35037 31076 35071
rect 31024 35028 31076 35037
rect 30932 35003 30984 35012
rect 30932 34969 30941 35003
rect 30941 34969 30975 35003
rect 30975 34969 30984 35003
rect 30932 34960 30984 34969
rect 22192 34892 22244 34944
rect 22468 34892 22520 34944
rect 23664 34935 23716 34944
rect 23664 34901 23673 34935
rect 23673 34901 23707 34935
rect 23707 34901 23716 34935
rect 23664 34892 23716 34901
rect 26976 34935 27028 34944
rect 26976 34901 26985 34935
rect 26985 34901 27019 34935
rect 27019 34901 27028 34935
rect 26976 34892 27028 34901
rect 29184 34892 29236 34944
rect 30564 34935 30616 34944
rect 30564 34901 30573 34935
rect 30573 34901 30607 34935
rect 30607 34901 30616 34935
rect 30564 34892 30616 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 15844 34731 15896 34740
rect 15844 34697 15853 34731
rect 15853 34697 15887 34731
rect 15887 34697 15896 34731
rect 15844 34688 15896 34697
rect 22284 34688 22336 34740
rect 1584 34595 1636 34604
rect 1584 34561 1593 34595
rect 1593 34561 1627 34595
rect 1627 34561 1636 34595
rect 1584 34552 1636 34561
rect 14556 34595 14608 34604
rect 14556 34561 14565 34595
rect 14565 34561 14599 34595
rect 14599 34561 14608 34595
rect 14556 34552 14608 34561
rect 14740 34595 14792 34604
rect 14740 34561 14749 34595
rect 14749 34561 14783 34595
rect 14783 34561 14792 34595
rect 14740 34552 14792 34561
rect 22652 34688 22704 34740
rect 23388 34731 23440 34740
rect 23388 34697 23397 34731
rect 23397 34697 23431 34731
rect 23431 34697 23440 34731
rect 23388 34688 23440 34697
rect 24400 34731 24452 34740
rect 24400 34697 24409 34731
rect 24409 34697 24443 34731
rect 24443 34697 24452 34731
rect 24400 34688 24452 34697
rect 25688 34688 25740 34740
rect 15200 34484 15252 34536
rect 18696 34484 18748 34536
rect 21456 34484 21508 34536
rect 22192 34484 22244 34536
rect 22560 34595 22612 34604
rect 22560 34561 22569 34595
rect 22569 34561 22603 34595
rect 22603 34561 22612 34595
rect 24584 34595 24636 34604
rect 22560 34552 22612 34561
rect 24584 34561 24593 34595
rect 24593 34561 24627 34595
rect 24627 34561 24636 34595
rect 24584 34552 24636 34561
rect 26976 34620 27028 34672
rect 28356 34688 28408 34740
rect 29000 34731 29052 34740
rect 29000 34697 29009 34731
rect 29009 34697 29043 34731
rect 29043 34697 29052 34731
rect 29000 34688 29052 34697
rect 30104 34620 30156 34672
rect 30564 34663 30616 34672
rect 30564 34629 30598 34663
rect 30598 34629 30616 34663
rect 30564 34620 30616 34629
rect 25136 34552 25188 34604
rect 25412 34552 25464 34604
rect 25964 34484 26016 34536
rect 26700 34552 26752 34604
rect 27068 34552 27120 34604
rect 26332 34527 26384 34536
rect 25872 34459 25924 34468
rect 25872 34425 25881 34459
rect 25881 34425 25915 34459
rect 25915 34425 25924 34459
rect 25872 34416 25924 34425
rect 26332 34493 26341 34527
rect 26341 34493 26375 34527
rect 26375 34493 26384 34527
rect 26332 34484 26384 34493
rect 28172 34552 28224 34604
rect 29184 34595 29236 34604
rect 29184 34561 29193 34595
rect 29193 34561 29227 34595
rect 29227 34561 29236 34595
rect 29184 34552 29236 34561
rect 30288 34595 30340 34604
rect 30288 34561 30297 34595
rect 30297 34561 30331 34595
rect 30331 34561 30340 34595
rect 30288 34552 30340 34561
rect 29368 34527 29420 34536
rect 29368 34493 29377 34527
rect 29377 34493 29411 34527
rect 29411 34493 29420 34527
rect 29368 34484 29420 34493
rect 30840 34552 30892 34604
rect 32220 34552 32272 34604
rect 1768 34391 1820 34400
rect 1768 34357 1777 34391
rect 1777 34357 1811 34391
rect 1811 34357 1820 34391
rect 1768 34348 1820 34357
rect 15016 34348 15068 34400
rect 22560 34348 22612 34400
rect 31392 34348 31444 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 1768 34144 1820 34196
rect 12992 34144 13044 34196
rect 13728 34144 13780 34196
rect 11796 34051 11848 34060
rect 11796 34017 11805 34051
rect 11805 34017 11839 34051
rect 11839 34017 11848 34051
rect 11796 34008 11848 34017
rect 22100 34144 22152 34196
rect 22652 34187 22704 34196
rect 22652 34153 22661 34187
rect 22661 34153 22695 34187
rect 22695 34153 22704 34187
rect 22652 34144 22704 34153
rect 27160 34144 27212 34196
rect 30748 34144 30800 34196
rect 31024 34144 31076 34196
rect 15016 33983 15068 33992
rect 15016 33949 15025 33983
rect 15025 33949 15059 33983
rect 15059 33949 15068 33983
rect 15200 33983 15252 33992
rect 15016 33940 15068 33949
rect 15200 33949 15209 33983
rect 15209 33949 15243 33983
rect 15243 33949 15252 33983
rect 15200 33940 15252 33949
rect 15384 33940 15436 33992
rect 17500 33940 17552 33992
rect 20168 33983 20220 33992
rect 20168 33949 20177 33983
rect 20177 33949 20211 33983
rect 20211 33949 20220 33983
rect 20168 33940 20220 33949
rect 20536 34008 20588 34060
rect 20812 34008 20864 34060
rect 21456 33940 21508 33992
rect 21640 33940 21692 33992
rect 22468 33940 22520 33992
rect 23664 34008 23716 34060
rect 22744 33983 22796 33992
rect 22744 33949 22753 33983
rect 22753 33949 22787 33983
rect 22787 33949 22796 33983
rect 22744 33940 22796 33949
rect 26884 33940 26936 33992
rect 12072 33915 12124 33924
rect 12072 33881 12106 33915
rect 12106 33881 12124 33915
rect 12072 33872 12124 33881
rect 16856 33872 16908 33924
rect 27068 33872 27120 33924
rect 28356 33940 28408 33992
rect 31392 34008 31444 34060
rect 30196 33983 30248 33992
rect 30196 33949 30205 33983
rect 30205 33949 30239 33983
rect 30239 33949 30248 33983
rect 30196 33940 30248 33949
rect 31300 33983 31352 33992
rect 30104 33915 30156 33924
rect 30104 33881 30113 33915
rect 30113 33881 30147 33915
rect 30147 33881 30156 33915
rect 30104 33872 30156 33881
rect 31300 33949 31309 33983
rect 31309 33949 31343 33983
rect 31343 33949 31352 33983
rect 31300 33940 31352 33949
rect 31760 33940 31812 33992
rect 31576 33872 31628 33924
rect 15752 33804 15804 33856
rect 17132 33847 17184 33856
rect 17132 33813 17141 33847
rect 17141 33813 17175 33847
rect 17175 33813 17184 33847
rect 17132 33804 17184 33813
rect 19984 33847 20036 33856
rect 19984 33813 19993 33847
rect 19993 33813 20027 33847
rect 20027 33813 20036 33847
rect 19984 33804 20036 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 12072 33600 12124 33652
rect 16856 33643 16908 33652
rect 11796 33532 11848 33584
rect 16856 33609 16865 33643
rect 16865 33609 16899 33643
rect 16899 33609 16908 33643
rect 16856 33600 16908 33609
rect 20904 33643 20956 33652
rect 20904 33609 20913 33643
rect 20913 33609 20947 33643
rect 20947 33609 20956 33643
rect 20904 33600 20956 33609
rect 12164 33507 12216 33516
rect 12164 33473 12173 33507
rect 12173 33473 12207 33507
rect 12207 33473 12216 33507
rect 12164 33464 12216 33473
rect 14740 33532 14792 33584
rect 14280 33464 14332 33516
rect 14924 33507 14976 33516
rect 14924 33473 14933 33507
rect 14933 33473 14967 33507
rect 14967 33473 14976 33507
rect 14924 33464 14976 33473
rect 17500 33532 17552 33584
rect 19432 33532 19484 33584
rect 17040 33507 17092 33516
rect 12440 33439 12492 33448
rect 12440 33405 12449 33439
rect 12449 33405 12483 33439
rect 12483 33405 12492 33439
rect 12440 33396 12492 33405
rect 12808 33396 12860 33448
rect 17040 33473 17049 33507
rect 17049 33473 17083 33507
rect 17083 33473 17092 33507
rect 17040 33464 17092 33473
rect 17224 33507 17276 33516
rect 17224 33473 17233 33507
rect 17233 33473 17267 33507
rect 17267 33473 17276 33507
rect 17224 33464 17276 33473
rect 18236 33507 18288 33516
rect 18236 33473 18245 33507
rect 18245 33473 18279 33507
rect 18279 33473 18288 33507
rect 18236 33464 18288 33473
rect 19984 33532 20036 33584
rect 31392 33507 31444 33516
rect 31392 33473 31401 33507
rect 31401 33473 31435 33507
rect 31435 33473 31444 33507
rect 31392 33464 31444 33473
rect 35900 33507 35952 33516
rect 35900 33473 35909 33507
rect 35909 33473 35943 33507
rect 35943 33473 35952 33507
rect 35900 33464 35952 33473
rect 17316 33439 17368 33448
rect 17316 33405 17325 33439
rect 17325 33405 17359 33439
rect 17359 33405 17368 33439
rect 17316 33396 17368 33405
rect 17960 33396 18012 33448
rect 19064 33396 19116 33448
rect 36636 33439 36688 33448
rect 36636 33405 36645 33439
rect 36645 33405 36679 33439
rect 36679 33405 36688 33439
rect 36636 33396 36688 33405
rect 15200 33328 15252 33380
rect 18604 33328 18656 33380
rect 31392 33328 31444 33380
rect 12532 33260 12584 33312
rect 13820 33260 13872 33312
rect 14464 33260 14516 33312
rect 18052 33303 18104 33312
rect 18052 33269 18061 33303
rect 18061 33269 18095 33303
rect 18095 33269 18104 33303
rect 18052 33260 18104 33269
rect 18328 33260 18380 33312
rect 21732 33260 21784 33312
rect 23204 33260 23256 33312
rect 31760 33260 31812 33312
rect 32220 33260 32272 33312
rect 47952 33303 48004 33312
rect 47952 33269 47961 33303
rect 47961 33269 47995 33303
rect 47995 33269 48004 33303
rect 47952 33260 48004 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 12164 33056 12216 33108
rect 14280 33099 14332 33108
rect 14280 33065 14289 33099
rect 14289 33065 14323 33099
rect 14323 33065 14332 33099
rect 14280 33056 14332 33065
rect 17040 33056 17092 33108
rect 20168 33056 20220 33108
rect 21916 33056 21968 33108
rect 22284 33056 22336 33108
rect 22836 33056 22888 33108
rect 2136 32852 2188 32904
rect 2504 32895 2556 32904
rect 2504 32861 2513 32895
rect 2513 32861 2547 32895
rect 2547 32861 2556 32895
rect 2504 32852 2556 32861
rect 5264 32852 5316 32904
rect 14924 32988 14976 33040
rect 22008 32988 22060 33040
rect 22100 32988 22152 33040
rect 26332 33056 26384 33108
rect 29368 33056 29420 33108
rect 31300 33056 31352 33108
rect 27068 32988 27120 33040
rect 31852 33031 31904 33040
rect 31852 32997 31861 33031
rect 31861 32997 31895 33031
rect 31895 32997 31904 33031
rect 31852 32988 31904 32997
rect 14372 32920 14424 32972
rect 15016 32920 15068 32972
rect 17500 32963 17552 32972
rect 17500 32929 17509 32963
rect 17509 32929 17543 32963
rect 17543 32929 17552 32963
rect 17500 32920 17552 32929
rect 12624 32852 12676 32904
rect 12992 32895 13044 32904
rect 12992 32861 13001 32895
rect 13001 32861 13035 32895
rect 13035 32861 13044 32895
rect 12992 32852 13044 32861
rect 14464 32895 14516 32904
rect 14464 32861 14473 32895
rect 14473 32861 14507 32895
rect 14507 32861 14516 32895
rect 14464 32852 14516 32861
rect 16856 32895 16908 32904
rect 12900 32784 12952 32836
rect 13820 32784 13872 32836
rect 16856 32861 16865 32895
rect 16865 32861 16899 32895
rect 16899 32861 16908 32895
rect 16856 32852 16908 32861
rect 17132 32852 17184 32904
rect 18052 32852 18104 32904
rect 18512 32852 18564 32904
rect 21548 32920 21600 32972
rect 24584 32963 24636 32972
rect 24584 32929 24593 32963
rect 24593 32929 24627 32963
rect 24627 32929 24636 32963
rect 24584 32920 24636 32929
rect 25596 32920 25648 32972
rect 30656 32920 30708 32972
rect 20996 32852 21048 32904
rect 21824 32895 21876 32904
rect 21824 32861 21833 32895
rect 21833 32861 21867 32895
rect 21867 32861 21876 32895
rect 21824 32852 21876 32861
rect 22284 32895 22336 32904
rect 22284 32861 22293 32895
rect 22293 32861 22327 32895
rect 22327 32861 22336 32895
rect 22284 32852 22336 32861
rect 23020 32852 23072 32904
rect 23204 32895 23256 32904
rect 23204 32861 23213 32895
rect 23213 32861 23247 32895
rect 23247 32861 23256 32895
rect 23204 32852 23256 32861
rect 2320 32716 2372 32768
rect 22376 32784 22428 32836
rect 23940 32784 23992 32836
rect 28540 32852 28592 32904
rect 31484 32920 31536 32972
rect 47952 32920 48004 32972
rect 31392 32895 31444 32904
rect 31392 32861 31401 32895
rect 31401 32861 31435 32895
rect 31435 32861 31444 32895
rect 31392 32852 31444 32861
rect 32220 32852 32272 32904
rect 31576 32784 31628 32836
rect 33508 32784 33560 32836
rect 47860 32784 47912 32836
rect 48320 32827 48372 32836
rect 48320 32793 48329 32827
rect 48329 32793 48363 32827
rect 48363 32793 48372 32827
rect 48320 32784 48372 32793
rect 18328 32716 18380 32768
rect 18880 32759 18932 32768
rect 18880 32725 18889 32759
rect 18889 32725 18923 32759
rect 18923 32725 18932 32759
rect 18880 32716 18932 32725
rect 21180 32716 21232 32768
rect 21732 32716 21784 32768
rect 22100 32716 22152 32768
rect 23388 32716 23440 32768
rect 29092 32716 29144 32768
rect 32128 32716 32180 32768
rect 47308 32716 47360 32768
rect 48136 32716 48188 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 12900 32512 12952 32564
rect 15200 32512 15252 32564
rect 17132 32512 17184 32564
rect 18236 32555 18288 32564
rect 18236 32521 18245 32555
rect 18245 32521 18279 32555
rect 18279 32521 18288 32555
rect 18236 32512 18288 32521
rect 23388 32555 23440 32564
rect 23388 32521 23397 32555
rect 23397 32521 23431 32555
rect 23431 32521 23440 32555
rect 23388 32512 23440 32521
rect 23940 32555 23992 32564
rect 23940 32521 23949 32555
rect 23949 32521 23983 32555
rect 23983 32521 23992 32555
rect 23940 32512 23992 32521
rect 24400 32512 24452 32564
rect 26424 32512 26476 32564
rect 2320 32487 2372 32496
rect 2320 32453 2329 32487
rect 2329 32453 2363 32487
rect 2363 32453 2372 32487
rect 2320 32444 2372 32453
rect 18604 32444 18656 32496
rect 26240 32444 26292 32496
rect 2136 32419 2188 32428
rect 2136 32385 2145 32419
rect 2145 32385 2179 32419
rect 2179 32385 2188 32419
rect 2136 32376 2188 32385
rect 14924 32376 14976 32428
rect 18512 32376 18564 32428
rect 18880 32419 18932 32428
rect 18880 32385 18889 32419
rect 18889 32385 18923 32419
rect 18923 32385 18932 32419
rect 18880 32376 18932 32385
rect 22008 32419 22060 32428
rect 22008 32385 22017 32419
rect 22017 32385 22051 32419
rect 22051 32385 22060 32419
rect 22008 32376 22060 32385
rect 22100 32376 22152 32428
rect 24952 32376 25004 32428
rect 25228 32376 25280 32428
rect 26332 32376 26384 32428
rect 2780 32351 2832 32360
rect 2780 32317 2789 32351
rect 2789 32317 2823 32351
rect 2823 32317 2832 32351
rect 2780 32308 2832 32317
rect 15844 32351 15896 32360
rect 15844 32317 15853 32351
rect 15853 32317 15887 32351
rect 15887 32317 15896 32351
rect 15844 32308 15896 32317
rect 16120 32308 16172 32360
rect 16856 32308 16908 32360
rect 17592 32308 17644 32360
rect 20076 32308 20128 32360
rect 24400 32351 24452 32360
rect 24400 32317 24409 32351
rect 24409 32317 24443 32351
rect 24443 32317 24452 32351
rect 24400 32308 24452 32317
rect 24584 32308 24636 32360
rect 30288 32444 30340 32496
rect 27252 32376 27304 32428
rect 29000 32419 29052 32428
rect 29000 32385 29009 32419
rect 29009 32385 29043 32419
rect 29043 32385 29052 32419
rect 29000 32376 29052 32385
rect 29092 32376 29144 32428
rect 31116 32419 31168 32428
rect 31116 32385 31125 32419
rect 31125 32385 31159 32419
rect 31159 32385 31168 32419
rect 31116 32376 31168 32385
rect 32680 32512 32732 32564
rect 47860 32555 47912 32564
rect 47860 32521 47869 32555
rect 47869 32521 47903 32555
rect 47903 32521 47912 32555
rect 47860 32512 47912 32521
rect 31668 32444 31720 32496
rect 31576 32419 31628 32428
rect 36636 32444 36688 32496
rect 31576 32385 31590 32419
rect 31590 32385 31624 32419
rect 31624 32385 31628 32419
rect 31576 32376 31628 32385
rect 48136 32376 48188 32428
rect 15384 32215 15436 32224
rect 15384 32181 15393 32215
rect 15393 32181 15427 32215
rect 15427 32181 15436 32215
rect 15384 32172 15436 32181
rect 24308 32215 24360 32224
rect 24308 32181 24317 32215
rect 24317 32181 24351 32215
rect 24351 32181 24360 32215
rect 24308 32172 24360 32181
rect 27436 32172 27488 32224
rect 30380 32215 30432 32224
rect 30380 32181 30389 32215
rect 30389 32181 30423 32215
rect 30423 32181 30432 32215
rect 30380 32172 30432 32181
rect 32680 32172 32732 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 21916 32011 21968 32020
rect 21916 31977 21925 32011
rect 21925 31977 21959 32011
rect 21959 31977 21968 32011
rect 21916 31968 21968 31977
rect 23940 32011 23992 32020
rect 23940 31977 23949 32011
rect 23949 31977 23983 32011
rect 23983 31977 23992 32011
rect 23940 31968 23992 31977
rect 24308 31968 24360 32020
rect 24952 31968 25004 32020
rect 25320 31968 25372 32020
rect 25964 32011 26016 32020
rect 25964 31977 25973 32011
rect 25973 31977 26007 32011
rect 26007 31977 26016 32011
rect 25964 31968 26016 31977
rect 1584 31875 1636 31884
rect 1584 31841 1593 31875
rect 1593 31841 1627 31875
rect 1627 31841 1636 31875
rect 1584 31832 1636 31841
rect 6644 31764 6696 31816
rect 13820 31764 13872 31816
rect 17132 31832 17184 31884
rect 19432 31832 19484 31884
rect 16488 31807 16540 31816
rect 16488 31773 16497 31807
rect 16497 31773 16531 31807
rect 16531 31773 16540 31807
rect 16488 31764 16540 31773
rect 21824 31764 21876 31816
rect 24584 31875 24636 31884
rect 20996 31696 21048 31748
rect 22376 31696 22428 31748
rect 23388 31764 23440 31816
rect 23756 31807 23808 31816
rect 23756 31773 23765 31807
rect 23765 31773 23799 31807
rect 23799 31773 23808 31807
rect 23756 31764 23808 31773
rect 24584 31841 24593 31875
rect 24593 31841 24627 31875
rect 24627 31841 24636 31875
rect 24584 31832 24636 31841
rect 27804 31968 27856 32020
rect 28540 32011 28592 32020
rect 28540 31977 28549 32011
rect 28549 31977 28583 32011
rect 28583 31977 28592 32011
rect 28540 31968 28592 31977
rect 31116 31968 31168 32020
rect 32220 31968 32272 32020
rect 30472 31900 30524 31952
rect 27068 31832 27120 31884
rect 32128 31875 32180 31884
rect 26884 31764 26936 31816
rect 32128 31841 32137 31875
rect 32137 31841 32171 31875
rect 32171 31841 32180 31875
rect 32128 31832 32180 31841
rect 27436 31807 27488 31816
rect 27436 31773 27445 31807
rect 27445 31773 27479 31807
rect 27479 31773 27488 31807
rect 27436 31764 27488 31773
rect 28724 31807 28776 31816
rect 28724 31773 28733 31807
rect 28733 31773 28767 31807
rect 28767 31773 28776 31807
rect 28724 31764 28776 31773
rect 29092 31764 29144 31816
rect 30380 31764 30432 31816
rect 31852 31807 31904 31816
rect 31852 31773 31861 31807
rect 31861 31773 31895 31807
rect 31895 31773 31904 31807
rect 31852 31764 31904 31773
rect 32772 31807 32824 31816
rect 32772 31773 32781 31807
rect 32781 31773 32815 31807
rect 32815 31773 32824 31807
rect 32772 31764 32824 31773
rect 32588 31739 32640 31748
rect 12440 31671 12492 31680
rect 12440 31637 12449 31671
rect 12449 31637 12483 31671
rect 12483 31637 12492 31671
rect 12440 31628 12492 31637
rect 16764 31628 16816 31680
rect 22284 31628 22336 31680
rect 32588 31705 32597 31739
rect 32597 31705 32631 31739
rect 32631 31705 32640 31739
rect 32588 31696 32640 31705
rect 25228 31628 25280 31680
rect 26792 31671 26844 31680
rect 26792 31637 26801 31671
rect 26801 31637 26835 31671
rect 26835 31637 26844 31671
rect 26792 31628 26844 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 13820 31467 13872 31476
rect 13820 31433 13829 31467
rect 13829 31433 13863 31467
rect 13863 31433 13872 31467
rect 13820 31424 13872 31433
rect 15384 31424 15436 31476
rect 20996 31467 21048 31476
rect 20996 31433 21005 31467
rect 21005 31433 21039 31467
rect 21039 31433 21048 31467
rect 20996 31424 21048 31433
rect 22100 31467 22152 31476
rect 22100 31433 22109 31467
rect 22109 31433 22143 31467
rect 22143 31433 22152 31467
rect 22100 31424 22152 31433
rect 23756 31424 23808 31476
rect 27252 31424 27304 31476
rect 31392 31424 31444 31476
rect 12440 31356 12492 31408
rect 12624 31356 12676 31408
rect 17316 31356 17368 31408
rect 6000 31288 6052 31340
rect 8392 31331 8444 31340
rect 8392 31297 8401 31331
rect 8401 31297 8435 31331
rect 8435 31297 8444 31331
rect 8392 31288 8444 31297
rect 11796 31288 11848 31340
rect 16856 31331 16908 31340
rect 16856 31297 16865 31331
rect 16865 31297 16899 31331
rect 16899 31297 16908 31331
rect 16856 31288 16908 31297
rect 17040 31331 17092 31340
rect 17040 31297 17049 31331
rect 17049 31297 17083 31331
rect 17083 31297 17092 31331
rect 17040 31288 17092 31297
rect 17592 31331 17644 31340
rect 17592 31297 17601 31331
rect 17601 31297 17635 31331
rect 17635 31297 17644 31331
rect 17592 31288 17644 31297
rect 21180 31331 21232 31340
rect 14096 31220 14148 31272
rect 14464 31263 14516 31272
rect 14464 31229 14473 31263
rect 14473 31229 14507 31263
rect 14507 31229 14516 31263
rect 14464 31220 14516 31229
rect 15568 31263 15620 31272
rect 15568 31229 15577 31263
rect 15577 31229 15611 31263
rect 15611 31229 15620 31263
rect 15568 31220 15620 31229
rect 15844 31263 15896 31272
rect 15844 31229 15853 31263
rect 15853 31229 15887 31263
rect 15887 31229 15896 31263
rect 15844 31220 15896 31229
rect 16580 31220 16632 31272
rect 21180 31297 21189 31331
rect 21189 31297 21223 31331
rect 21223 31297 21232 31331
rect 21180 31288 21232 31297
rect 22284 31331 22336 31340
rect 22284 31297 22293 31331
rect 22293 31297 22327 31331
rect 22327 31297 22336 31331
rect 22284 31288 22336 31297
rect 24860 31331 24912 31340
rect 24860 31297 24869 31331
rect 24869 31297 24903 31331
rect 24903 31297 24912 31331
rect 24860 31288 24912 31297
rect 25320 31331 25372 31340
rect 21548 31220 21600 31272
rect 22468 31220 22520 31272
rect 23204 31220 23256 31272
rect 25320 31297 25329 31331
rect 25329 31297 25363 31331
rect 25363 31297 25372 31331
rect 25320 31288 25372 31297
rect 26792 31288 26844 31340
rect 29000 31288 29052 31340
rect 30196 31331 30248 31340
rect 30196 31297 30230 31331
rect 30230 31297 30248 31331
rect 30196 31288 30248 31297
rect 32128 31288 32180 31340
rect 25228 31220 25280 31272
rect 27804 31220 27856 31272
rect 32680 31220 32732 31272
rect 32772 31220 32824 31272
rect 13636 31152 13688 31204
rect 4712 31084 4764 31136
rect 5356 31084 5408 31136
rect 8208 31127 8260 31136
rect 8208 31093 8217 31127
rect 8217 31093 8251 31127
rect 8251 31093 8260 31127
rect 8208 31084 8260 31093
rect 13544 31084 13596 31136
rect 16488 31084 16540 31136
rect 22376 31152 22428 31204
rect 20444 31084 20496 31136
rect 23940 31084 23992 31136
rect 24768 31084 24820 31136
rect 27528 31127 27580 31136
rect 27528 31093 27537 31127
rect 27537 31093 27571 31127
rect 27571 31093 27580 31127
rect 27528 31084 27580 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 5356 30923 5408 30932
rect 5356 30889 5365 30923
rect 5365 30889 5399 30923
rect 5399 30889 5408 30923
rect 5356 30880 5408 30889
rect 6000 30923 6052 30932
rect 6000 30889 6009 30923
rect 6009 30889 6043 30923
rect 6043 30889 6052 30923
rect 6000 30880 6052 30889
rect 12532 30923 12584 30932
rect 6920 30744 6972 30796
rect 12532 30889 12541 30923
rect 12541 30889 12575 30923
rect 12575 30889 12584 30923
rect 12532 30880 12584 30889
rect 15568 30880 15620 30932
rect 17960 30880 18012 30932
rect 19248 30880 19300 30932
rect 32588 30880 32640 30932
rect 9128 30787 9180 30796
rect 9128 30753 9137 30787
rect 9137 30753 9171 30787
rect 9171 30753 9180 30787
rect 9128 30744 9180 30753
rect 5172 30676 5224 30728
rect 6184 30719 6236 30728
rect 6184 30685 6193 30719
rect 6193 30685 6227 30719
rect 6227 30685 6236 30719
rect 6184 30676 6236 30685
rect 8208 30676 8260 30728
rect 15936 30812 15988 30864
rect 16304 30855 16356 30864
rect 16304 30821 16313 30855
rect 16313 30821 16347 30855
rect 16347 30821 16356 30855
rect 16304 30812 16356 30821
rect 16580 30812 16632 30864
rect 16764 30812 16816 30864
rect 17592 30812 17644 30864
rect 1860 30608 1912 30660
rect 12440 30676 12492 30728
rect 12624 30719 12676 30728
rect 12624 30685 12633 30719
rect 12633 30685 12667 30719
rect 12667 30685 12676 30719
rect 12624 30676 12676 30685
rect 13544 30719 13596 30728
rect 13544 30685 13553 30719
rect 13553 30685 13587 30719
rect 13587 30685 13596 30719
rect 13544 30676 13596 30685
rect 13728 30719 13780 30728
rect 13728 30685 13737 30719
rect 13737 30685 13771 30719
rect 13771 30685 13780 30719
rect 13728 30676 13780 30685
rect 9496 30608 9548 30660
rect 5540 30583 5592 30592
rect 5540 30549 5549 30583
rect 5549 30549 5583 30583
rect 5583 30549 5592 30583
rect 5540 30540 5592 30549
rect 7840 30540 7892 30592
rect 9128 30540 9180 30592
rect 13636 30608 13688 30660
rect 15476 30676 15528 30728
rect 16488 30676 16540 30728
rect 19432 30787 19484 30796
rect 19432 30753 19441 30787
rect 19441 30753 19475 30787
rect 19475 30753 19484 30787
rect 19432 30744 19484 30753
rect 28080 30744 28132 30796
rect 16948 30719 17000 30728
rect 16948 30685 16957 30719
rect 16957 30685 16991 30719
rect 16991 30685 17000 30719
rect 16948 30676 17000 30685
rect 17684 30676 17736 30728
rect 30564 30719 30616 30728
rect 17868 30608 17920 30660
rect 19340 30608 19392 30660
rect 30564 30685 30573 30719
rect 30573 30685 30607 30719
rect 30607 30685 30616 30719
rect 30564 30676 30616 30685
rect 30748 30676 30800 30728
rect 31392 30676 31444 30728
rect 32128 30719 32180 30728
rect 32128 30685 32137 30719
rect 32137 30685 32171 30719
rect 32171 30685 32180 30719
rect 32128 30676 32180 30685
rect 32680 30676 32732 30728
rect 30104 30608 30156 30660
rect 10508 30583 10560 30592
rect 10508 30549 10517 30583
rect 10517 30549 10551 30583
rect 10551 30549 10560 30583
rect 10508 30540 10560 30549
rect 12256 30540 12308 30592
rect 15200 30540 15252 30592
rect 16304 30540 16356 30592
rect 18052 30583 18104 30592
rect 18052 30549 18061 30583
rect 18061 30549 18095 30583
rect 18095 30549 18104 30583
rect 18052 30540 18104 30549
rect 18604 30540 18656 30592
rect 18788 30540 18840 30592
rect 28816 30583 28868 30592
rect 28816 30549 28825 30583
rect 28825 30549 28859 30583
rect 28859 30549 28868 30583
rect 28816 30540 28868 30549
rect 30380 30583 30432 30592
rect 30380 30549 30389 30583
rect 30389 30549 30423 30583
rect 30423 30549 30432 30583
rect 30380 30540 30432 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 5540 30336 5592 30388
rect 6184 30336 6236 30388
rect 6644 30311 6696 30320
rect 6644 30277 6653 30311
rect 6653 30277 6687 30311
rect 6687 30277 6696 30311
rect 8392 30336 8444 30388
rect 9496 30379 9548 30388
rect 9496 30345 9505 30379
rect 9505 30345 9539 30379
rect 9539 30345 9548 30379
rect 9496 30336 9548 30345
rect 16948 30336 17000 30388
rect 17868 30336 17920 30388
rect 19248 30336 19300 30388
rect 23296 30336 23348 30388
rect 23756 30336 23808 30388
rect 30196 30379 30248 30388
rect 30196 30345 30205 30379
rect 30205 30345 30239 30379
rect 30239 30345 30248 30379
rect 30196 30336 30248 30345
rect 6644 30268 6696 30277
rect 11888 30268 11940 30320
rect 17040 30311 17092 30320
rect 17040 30277 17049 30311
rect 17049 30277 17083 30311
rect 17083 30277 17092 30311
rect 17040 30268 17092 30277
rect 17132 30268 17184 30320
rect 18052 30268 18104 30320
rect 18512 30268 18564 30320
rect 5172 30200 5224 30252
rect 7380 30200 7432 30252
rect 7840 30200 7892 30252
rect 7748 30175 7800 30184
rect 4896 30039 4948 30048
rect 4896 30005 4905 30039
rect 4905 30005 4939 30039
rect 4939 30005 4948 30039
rect 4896 29996 4948 30005
rect 7748 30141 7757 30175
rect 7757 30141 7791 30175
rect 7791 30141 7800 30175
rect 8668 30200 8720 30252
rect 12256 30243 12308 30252
rect 12256 30209 12290 30243
rect 12290 30209 12308 30243
rect 12256 30200 12308 30209
rect 15200 30243 15252 30252
rect 15200 30209 15209 30243
rect 15209 30209 15243 30243
rect 15243 30209 15252 30243
rect 15200 30200 15252 30209
rect 15476 30243 15528 30252
rect 15476 30209 15485 30243
rect 15485 30209 15519 30243
rect 15519 30209 15528 30243
rect 15476 30200 15528 30209
rect 16856 30243 16908 30252
rect 16856 30209 16865 30243
rect 16865 30209 16899 30243
rect 16899 30209 16908 30243
rect 16856 30200 16908 30209
rect 17684 30243 17736 30252
rect 17684 30209 17693 30243
rect 17693 30209 17727 30243
rect 17727 30209 17736 30243
rect 17684 30200 17736 30209
rect 17868 30243 17920 30252
rect 17868 30209 17877 30243
rect 17877 30209 17911 30243
rect 17911 30209 17920 30243
rect 17868 30200 17920 30209
rect 18604 30243 18656 30252
rect 18604 30209 18613 30243
rect 18613 30209 18647 30243
rect 18647 30209 18656 30243
rect 18604 30200 18656 30209
rect 18788 30243 18840 30252
rect 18788 30209 18795 30243
rect 18795 30209 18840 30243
rect 18788 30200 18840 30209
rect 11980 30175 12032 30184
rect 7748 30132 7800 30141
rect 11980 30141 11989 30175
rect 11989 30141 12023 30175
rect 12023 30141 12032 30175
rect 11980 30132 12032 30141
rect 19432 30268 19484 30320
rect 22376 30311 22428 30320
rect 22376 30277 22385 30311
rect 22385 30277 22419 30311
rect 22419 30277 22428 30311
rect 22376 30268 22428 30277
rect 23020 30268 23072 30320
rect 19064 30243 19116 30252
rect 19064 30209 19078 30243
rect 19078 30209 19112 30243
rect 19112 30209 19116 30243
rect 19064 30200 19116 30209
rect 20628 30200 20680 30252
rect 20260 30132 20312 30184
rect 22468 30243 22520 30252
rect 22468 30209 22477 30243
rect 22477 30209 22511 30243
rect 22511 30209 22520 30243
rect 22468 30200 22520 30209
rect 23572 30268 23624 30320
rect 7472 30064 7524 30116
rect 8392 29996 8444 30048
rect 10508 29996 10560 30048
rect 13084 29996 13136 30048
rect 13728 29996 13780 30048
rect 16764 30064 16816 30116
rect 17684 30064 17736 30116
rect 19340 30064 19392 30116
rect 19524 30064 19576 30116
rect 22560 30064 22612 30116
rect 22652 30064 22704 30116
rect 25136 30268 25188 30320
rect 26608 30268 26660 30320
rect 27896 30311 27948 30320
rect 27896 30277 27905 30311
rect 27905 30277 27939 30311
rect 27939 30277 27948 30311
rect 27896 30268 27948 30277
rect 41328 30268 41380 30320
rect 47676 30268 47728 30320
rect 25688 30200 25740 30252
rect 26240 30200 26292 30252
rect 26516 30243 26568 30252
rect 26516 30209 26525 30243
rect 26525 30209 26559 30243
rect 26559 30209 26568 30243
rect 26516 30200 26568 30209
rect 28080 30243 28132 30252
rect 28080 30209 28089 30243
rect 28089 30209 28123 30243
rect 28123 30209 28132 30243
rect 28080 30200 28132 30209
rect 28816 30200 28868 30252
rect 30380 30243 30432 30252
rect 30380 30209 30389 30243
rect 30389 30209 30423 30243
rect 30423 30209 30432 30243
rect 30380 30200 30432 30209
rect 30840 30200 30892 30252
rect 30472 30132 30524 30184
rect 32864 30200 32916 30252
rect 47308 30200 47360 30252
rect 31852 30132 31904 30184
rect 15752 30039 15804 30048
rect 15752 30005 15761 30039
rect 15761 30005 15795 30039
rect 15795 30005 15804 30039
rect 15752 29996 15804 30005
rect 15936 29996 15988 30048
rect 21640 29996 21692 30048
rect 22376 29996 22428 30048
rect 22468 29996 22520 30048
rect 23296 30039 23348 30048
rect 23296 30005 23305 30039
rect 23305 30005 23339 30039
rect 23339 30005 23348 30039
rect 23296 29996 23348 30005
rect 26332 29996 26384 30048
rect 29276 29996 29328 30048
rect 31024 29996 31076 30048
rect 46480 29996 46532 30048
rect 47860 30039 47912 30048
rect 47860 30005 47869 30039
rect 47869 30005 47903 30039
rect 47903 30005 47912 30039
rect 47860 29996 47912 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 12440 29835 12492 29844
rect 12440 29801 12449 29835
rect 12449 29801 12483 29835
rect 12483 29801 12492 29835
rect 15752 29835 15804 29844
rect 12440 29792 12492 29801
rect 15752 29801 15761 29835
rect 15761 29801 15795 29835
rect 15795 29801 15804 29835
rect 15752 29792 15804 29801
rect 20628 29835 20680 29844
rect 20628 29801 20637 29835
rect 20637 29801 20671 29835
rect 20671 29801 20680 29835
rect 20628 29792 20680 29801
rect 22192 29792 22244 29844
rect 22376 29792 22428 29844
rect 23480 29792 23532 29844
rect 30104 29835 30156 29844
rect 6920 29699 6972 29708
rect 6920 29665 6929 29699
rect 6929 29665 6963 29699
rect 6963 29665 6972 29699
rect 6920 29656 6972 29665
rect 19524 29656 19576 29708
rect 22468 29724 22520 29776
rect 23296 29724 23348 29776
rect 30104 29801 30113 29835
rect 30113 29801 30147 29835
rect 30147 29801 30156 29835
rect 30104 29792 30156 29801
rect 31668 29724 31720 29776
rect 4896 29588 4948 29640
rect 12716 29588 12768 29640
rect 12900 29631 12952 29640
rect 12900 29597 12909 29631
rect 12909 29597 12943 29631
rect 12943 29597 12952 29631
rect 12900 29588 12952 29597
rect 13084 29631 13136 29640
rect 13084 29597 13093 29631
rect 13093 29597 13127 29631
rect 13127 29597 13136 29631
rect 13084 29588 13136 29597
rect 15936 29631 15988 29640
rect 15936 29597 15945 29631
rect 15945 29597 15979 29631
rect 15979 29597 15988 29631
rect 15936 29588 15988 29597
rect 16028 29588 16080 29640
rect 20720 29631 20772 29640
rect 4712 29520 4764 29572
rect 6920 29520 6972 29572
rect 7288 29520 7340 29572
rect 20720 29597 20729 29631
rect 20729 29597 20763 29631
rect 20763 29597 20772 29631
rect 20720 29588 20772 29597
rect 21272 29588 21324 29640
rect 21640 29699 21692 29708
rect 21640 29665 21649 29699
rect 21649 29665 21683 29699
rect 21683 29665 21692 29699
rect 21640 29656 21692 29665
rect 23664 29656 23716 29708
rect 24584 29656 24636 29708
rect 46480 29699 46532 29708
rect 5724 29495 5776 29504
rect 5724 29461 5733 29495
rect 5733 29461 5767 29495
rect 5767 29461 5776 29495
rect 5724 29452 5776 29461
rect 8300 29495 8352 29504
rect 8300 29461 8309 29495
rect 8309 29461 8343 29495
rect 8343 29461 8352 29495
rect 8300 29452 8352 29461
rect 16672 29452 16724 29504
rect 20720 29452 20772 29504
rect 21364 29452 21416 29504
rect 22836 29588 22888 29640
rect 23756 29588 23808 29640
rect 46480 29665 46489 29699
rect 46489 29665 46523 29699
rect 46523 29665 46532 29699
rect 46480 29656 46532 29665
rect 47860 29656 47912 29708
rect 23020 29520 23072 29572
rect 23388 29520 23440 29572
rect 24676 29520 24728 29572
rect 28540 29588 28592 29640
rect 23204 29452 23256 29504
rect 23664 29452 23716 29504
rect 24952 29495 25004 29504
rect 24952 29461 24961 29495
rect 24961 29461 24995 29495
rect 24995 29461 25004 29495
rect 24952 29452 25004 29461
rect 26148 29520 26200 29572
rect 27620 29563 27672 29572
rect 27620 29529 27654 29563
rect 27654 29529 27672 29563
rect 27620 29520 27672 29529
rect 26516 29452 26568 29504
rect 27988 29452 28040 29504
rect 48320 29563 48372 29572
rect 48320 29529 48329 29563
rect 48329 29529 48363 29563
rect 48363 29529 48372 29563
rect 48320 29520 48372 29529
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 7288 29291 7340 29300
rect 7288 29257 7297 29291
rect 7297 29257 7331 29291
rect 7331 29257 7340 29291
rect 7288 29248 7340 29257
rect 7840 29248 7892 29300
rect 8668 29291 8720 29300
rect 8668 29257 8677 29291
rect 8677 29257 8711 29291
rect 8711 29257 8720 29291
rect 8668 29248 8720 29257
rect 16580 29248 16632 29300
rect 19064 29248 19116 29300
rect 22836 29248 22888 29300
rect 16672 29180 16724 29232
rect 20720 29180 20772 29232
rect 5172 29155 5224 29164
rect 5172 29121 5181 29155
rect 5181 29121 5215 29155
rect 5215 29121 5224 29155
rect 5172 29112 5224 29121
rect 7472 29155 7524 29164
rect 7472 29121 7481 29155
rect 7481 29121 7515 29155
rect 7515 29121 7524 29155
rect 7472 29112 7524 29121
rect 7840 29112 7892 29164
rect 15384 29112 15436 29164
rect 15936 29155 15988 29164
rect 15936 29121 15945 29155
rect 15945 29121 15979 29155
rect 15979 29121 15988 29155
rect 15936 29112 15988 29121
rect 16028 29112 16080 29164
rect 18512 29112 18564 29164
rect 22376 29155 22428 29164
rect 22376 29121 22385 29155
rect 22385 29121 22419 29155
rect 22419 29121 22428 29155
rect 22376 29112 22428 29121
rect 22652 29155 22704 29164
rect 22652 29121 22661 29155
rect 22661 29121 22695 29155
rect 22695 29121 22704 29155
rect 22652 29112 22704 29121
rect 23204 29155 23256 29164
rect 23204 29121 23213 29155
rect 23213 29121 23247 29155
rect 23247 29121 23256 29155
rect 23204 29112 23256 29121
rect 23388 29155 23440 29164
rect 23388 29121 23395 29155
rect 23395 29121 23440 29155
rect 23388 29112 23440 29121
rect 23480 29155 23532 29164
rect 23480 29121 23489 29155
rect 23489 29121 23523 29155
rect 23523 29121 23532 29155
rect 23480 29112 23532 29121
rect 23756 29112 23808 29164
rect 24400 29180 24452 29232
rect 24676 29248 24728 29300
rect 26148 29291 26200 29300
rect 26148 29257 26157 29291
rect 26157 29257 26191 29291
rect 26191 29257 26200 29291
rect 26148 29248 26200 29257
rect 27988 29291 28040 29300
rect 27988 29257 27997 29291
rect 27997 29257 28031 29291
rect 28031 29257 28040 29291
rect 27988 29248 28040 29257
rect 29276 29291 29328 29300
rect 29276 29257 29285 29291
rect 29285 29257 29319 29291
rect 29319 29257 29328 29291
rect 29276 29248 29328 29257
rect 25044 29180 25096 29232
rect 8392 29044 8444 29096
rect 9220 29044 9272 29096
rect 16948 29044 17000 29096
rect 26332 29155 26384 29164
rect 26332 29121 26341 29155
rect 26341 29121 26375 29155
rect 26375 29121 26384 29155
rect 26332 29112 26384 29121
rect 27528 29112 27580 29164
rect 27896 29112 27948 29164
rect 29184 29155 29236 29164
rect 29184 29121 29193 29155
rect 29193 29121 29227 29155
rect 29227 29121 29236 29155
rect 29184 29112 29236 29121
rect 30840 29155 30892 29164
rect 30840 29121 30849 29155
rect 30849 29121 30883 29155
rect 30883 29121 30892 29155
rect 30840 29112 30892 29121
rect 5724 28976 5776 29028
rect 21272 29019 21324 29028
rect 21272 28985 21281 29019
rect 21281 28985 21315 29019
rect 21315 28985 21324 29019
rect 21272 28976 21324 28985
rect 22100 28976 22152 29028
rect 23664 28976 23716 29028
rect 5632 28951 5684 28960
rect 5632 28917 5641 28951
rect 5641 28917 5675 28951
rect 5675 28917 5684 28951
rect 5632 28908 5684 28917
rect 8300 28951 8352 28960
rect 8300 28917 8309 28951
rect 8309 28917 8343 28951
rect 8343 28917 8352 28951
rect 8300 28908 8352 28917
rect 16948 28908 17000 28960
rect 17224 28951 17276 28960
rect 17224 28917 17233 28951
rect 17233 28917 17267 28951
rect 17267 28917 17276 28951
rect 17224 28908 17276 28917
rect 22376 28908 22428 28960
rect 25412 28908 25464 28960
rect 28172 29087 28224 29096
rect 28172 29053 28181 29087
rect 28181 29053 28215 29087
rect 28215 29053 28224 29087
rect 28172 29044 28224 29053
rect 30656 29044 30708 29096
rect 33416 29112 33468 29164
rect 38016 29112 38068 29164
rect 47676 29112 47728 29164
rect 31024 29019 31076 29028
rect 26700 28908 26752 28960
rect 31024 28985 31033 29019
rect 31033 28985 31067 29019
rect 31067 28985 31076 29019
rect 31024 28976 31076 28985
rect 31852 28976 31904 29028
rect 38476 28976 38528 29028
rect 27712 28908 27764 28960
rect 30656 28951 30708 28960
rect 30656 28917 30665 28951
rect 30665 28917 30699 28951
rect 30699 28917 30708 28951
rect 30656 28908 30708 28917
rect 47216 28951 47268 28960
rect 47216 28917 47225 28951
rect 47225 28917 47259 28951
rect 47259 28917 47268 28951
rect 47216 28908 47268 28917
rect 47860 28951 47912 28960
rect 47860 28917 47869 28951
rect 47869 28917 47903 28951
rect 47903 28917 47912 28951
rect 47860 28908 47912 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 9220 28747 9272 28756
rect 9220 28713 9229 28747
rect 9229 28713 9263 28747
rect 9263 28713 9272 28747
rect 9220 28704 9272 28713
rect 13820 28704 13872 28756
rect 14464 28704 14516 28756
rect 23572 28747 23624 28756
rect 14556 28568 14608 28620
rect 23572 28713 23581 28747
rect 23581 28713 23615 28747
rect 23615 28713 23624 28747
rect 23572 28704 23624 28713
rect 27620 28704 27672 28756
rect 28080 28704 28132 28756
rect 32128 28747 32180 28756
rect 32128 28713 32137 28747
rect 32137 28713 32171 28747
rect 32171 28713 32180 28747
rect 32128 28704 32180 28713
rect 5632 28500 5684 28552
rect 9404 28500 9456 28552
rect 13452 28543 13504 28552
rect 13452 28509 13461 28543
rect 13461 28509 13495 28543
rect 13495 28509 13504 28543
rect 13452 28500 13504 28509
rect 13636 28543 13688 28552
rect 13636 28509 13645 28543
rect 13645 28509 13679 28543
rect 13679 28509 13688 28543
rect 13636 28500 13688 28509
rect 14832 28432 14884 28484
rect 15752 28500 15804 28552
rect 15844 28500 15896 28552
rect 16580 28500 16632 28552
rect 16948 28500 17000 28552
rect 17408 28500 17460 28552
rect 22652 28568 22704 28620
rect 22100 28543 22152 28552
rect 22100 28509 22109 28543
rect 22109 28509 22143 28543
rect 22143 28509 22152 28543
rect 22100 28500 22152 28509
rect 22284 28500 22336 28552
rect 24952 28568 25004 28620
rect 27160 28568 27212 28620
rect 47216 28568 47268 28620
rect 48228 28611 48280 28620
rect 48228 28577 48237 28611
rect 48237 28577 48271 28611
rect 48271 28577 48280 28611
rect 48228 28568 48280 28577
rect 23664 28543 23716 28552
rect 23664 28509 23673 28543
rect 23673 28509 23707 28543
rect 23707 28509 23716 28543
rect 23664 28500 23716 28509
rect 27712 28543 27764 28552
rect 27712 28509 27721 28543
rect 27721 28509 27755 28543
rect 27755 28509 27764 28543
rect 27712 28500 27764 28509
rect 27988 28500 28040 28552
rect 28540 28543 28592 28552
rect 28540 28509 28549 28543
rect 28549 28509 28583 28543
rect 28583 28509 28592 28543
rect 28540 28500 28592 28509
rect 30656 28500 30708 28552
rect 35900 28500 35952 28552
rect 18788 28432 18840 28484
rect 4988 28407 5040 28416
rect 4988 28373 4997 28407
rect 4997 28373 5031 28407
rect 5031 28373 5040 28407
rect 4988 28364 5040 28373
rect 13544 28407 13596 28416
rect 13544 28373 13553 28407
rect 13553 28373 13587 28407
rect 13587 28373 13596 28407
rect 13544 28364 13596 28373
rect 15200 28407 15252 28416
rect 15200 28373 15209 28407
rect 15209 28373 15243 28407
rect 15243 28373 15252 28407
rect 15200 28364 15252 28373
rect 16212 28407 16264 28416
rect 16212 28373 16221 28407
rect 16221 28373 16255 28407
rect 16255 28373 16264 28407
rect 16212 28364 16264 28373
rect 16672 28364 16724 28416
rect 17500 28364 17552 28416
rect 18420 28364 18472 28416
rect 20168 28364 20220 28416
rect 20812 28407 20864 28416
rect 20812 28373 20821 28407
rect 20821 28373 20855 28407
rect 20855 28373 20864 28407
rect 20812 28364 20864 28373
rect 20904 28407 20956 28416
rect 20904 28373 20913 28407
rect 20913 28373 20947 28407
rect 20947 28373 20956 28407
rect 22192 28407 22244 28416
rect 38108 28432 38160 28484
rect 47860 28432 47912 28484
rect 20904 28364 20956 28373
rect 22192 28373 22207 28407
rect 22207 28373 22241 28407
rect 22241 28373 22244 28407
rect 22192 28364 22244 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 4712 28160 4764 28212
rect 13452 28160 13504 28212
rect 16028 28160 16080 28212
rect 4988 28092 5040 28144
rect 6920 28092 6972 28144
rect 14556 28135 14608 28144
rect 14556 28101 14565 28135
rect 14565 28101 14599 28135
rect 14599 28101 14608 28135
rect 14556 28092 14608 28101
rect 15476 28092 15528 28144
rect 9404 28024 9456 28076
rect 12808 28024 12860 28076
rect 12992 28024 13044 28076
rect 14372 28024 14424 28076
rect 8852 27999 8904 28008
rect 8852 27965 8861 27999
rect 8861 27965 8895 27999
rect 8895 27965 8904 27999
rect 8852 27956 8904 27965
rect 13820 27956 13872 28008
rect 14832 28067 14884 28076
rect 14832 28033 14841 28067
rect 14841 28033 14875 28067
rect 14875 28033 14884 28067
rect 17960 28092 18012 28144
rect 14832 28024 14884 28033
rect 9588 27888 9640 27940
rect 15844 27956 15896 28008
rect 15752 27888 15804 27940
rect 4988 27820 5040 27872
rect 8024 27863 8076 27872
rect 8024 27829 8033 27863
rect 8033 27829 8067 27863
rect 8067 27829 8076 27863
rect 8024 27820 8076 27829
rect 12716 27820 12768 27872
rect 14556 27863 14608 27872
rect 14556 27829 14565 27863
rect 14565 27829 14599 27863
rect 14599 27829 14608 27863
rect 14556 27820 14608 27829
rect 15568 27820 15620 27872
rect 17224 28024 17276 28076
rect 18788 28160 18840 28212
rect 20812 28203 20864 28212
rect 20812 28169 20821 28203
rect 20821 28169 20855 28203
rect 20855 28169 20864 28203
rect 20812 28160 20864 28169
rect 20904 28160 20956 28212
rect 30840 28160 30892 28212
rect 18512 28135 18564 28144
rect 18512 28101 18521 28135
rect 18521 28101 18555 28135
rect 18555 28101 18564 28135
rect 18512 28092 18564 28101
rect 18420 28067 18472 28076
rect 18420 28033 18427 28067
rect 18427 28033 18472 28067
rect 18420 28024 18472 28033
rect 19064 28024 19116 28076
rect 19984 28024 20036 28076
rect 17408 27956 17460 28008
rect 19432 27999 19484 28008
rect 19432 27965 19441 27999
rect 19441 27965 19475 27999
rect 19475 27965 19484 27999
rect 19432 27956 19484 27965
rect 21364 28135 21416 28144
rect 21364 28101 21373 28135
rect 21373 28101 21407 28135
rect 21407 28101 21416 28135
rect 21364 28092 21416 28101
rect 30748 28092 30800 28144
rect 21456 28067 21508 28076
rect 21456 28033 21465 28067
rect 21465 28033 21499 28067
rect 21499 28033 21508 28067
rect 21456 28024 21508 28033
rect 22192 28024 22244 28076
rect 22376 28067 22428 28076
rect 22376 28033 22385 28067
rect 22385 28033 22419 28067
rect 22419 28033 22428 28067
rect 22652 28067 22704 28076
rect 22376 28024 22428 28033
rect 22652 28033 22661 28067
rect 22661 28033 22695 28067
rect 22695 28033 22704 28067
rect 22652 28024 22704 28033
rect 24584 28067 24636 28076
rect 24584 28033 24593 28067
rect 24593 28033 24627 28067
rect 24627 28033 24636 28067
rect 24584 28024 24636 28033
rect 21364 27956 21416 28008
rect 22560 27999 22612 28008
rect 22560 27965 22569 27999
rect 22569 27965 22603 27999
rect 22603 27965 22612 27999
rect 26700 28024 26752 28076
rect 30472 28024 30524 28076
rect 32128 28024 32180 28076
rect 47492 28024 47544 28076
rect 47768 28067 47820 28076
rect 47768 28033 47777 28067
rect 47777 28033 47811 28067
rect 47811 28033 47820 28067
rect 47768 28024 47820 28033
rect 22560 27956 22612 27965
rect 25412 27956 25464 28008
rect 16212 27820 16264 27872
rect 24768 27863 24820 27872
rect 24768 27829 24777 27863
rect 24777 27829 24811 27863
rect 24811 27829 24820 27863
rect 24768 27820 24820 27829
rect 24860 27820 24912 27872
rect 47216 27863 47268 27872
rect 47216 27829 47225 27863
rect 47225 27829 47259 27863
rect 47259 27829 47268 27863
rect 47216 27820 47268 27829
rect 47860 27863 47912 27872
rect 47860 27829 47869 27863
rect 47869 27829 47903 27863
rect 47903 27829 47912 27863
rect 47860 27820 47912 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 4988 27616 5040 27668
rect 5724 27659 5776 27668
rect 5724 27625 5733 27659
rect 5733 27625 5767 27659
rect 5767 27625 5776 27659
rect 5724 27616 5776 27625
rect 8392 27659 8444 27668
rect 8392 27625 8401 27659
rect 8401 27625 8435 27659
rect 8435 27625 8444 27659
rect 8392 27616 8444 27625
rect 19984 27659 20036 27668
rect 14372 27591 14424 27600
rect 14372 27557 14381 27591
rect 14381 27557 14415 27591
rect 14415 27557 14424 27591
rect 14372 27548 14424 27557
rect 15384 27591 15436 27600
rect 15384 27557 15393 27591
rect 15393 27557 15427 27591
rect 15427 27557 15436 27591
rect 15384 27548 15436 27557
rect 5172 27412 5224 27464
rect 11980 27480 12032 27532
rect 16120 27548 16172 27600
rect 16580 27548 16632 27600
rect 16856 27480 16908 27532
rect 19984 27625 19993 27659
rect 19993 27625 20027 27659
rect 20027 27625 20036 27659
rect 19984 27616 20036 27625
rect 21272 27548 21324 27600
rect 26608 27591 26660 27600
rect 26608 27557 26617 27591
rect 26617 27557 26651 27591
rect 26651 27557 26660 27591
rect 26608 27548 26660 27557
rect 29368 27548 29420 27600
rect 14556 27455 14608 27464
rect 7012 27344 7064 27396
rect 14556 27421 14565 27455
rect 14565 27421 14599 27455
rect 14599 27421 14608 27455
rect 14556 27412 14608 27421
rect 12532 27344 12584 27396
rect 15292 27412 15344 27464
rect 15568 27455 15620 27464
rect 15568 27421 15577 27455
rect 15577 27421 15611 27455
rect 15611 27421 15620 27455
rect 15568 27412 15620 27421
rect 15660 27455 15712 27464
rect 15660 27421 15669 27455
rect 15669 27421 15703 27455
rect 15703 27421 15712 27455
rect 15660 27412 15712 27421
rect 16580 27455 16632 27464
rect 15200 27344 15252 27396
rect 16580 27421 16589 27455
rect 16589 27421 16623 27455
rect 16623 27421 16632 27455
rect 16580 27412 16632 27421
rect 17500 27412 17552 27464
rect 22560 27480 22612 27532
rect 47216 27480 47268 27532
rect 48228 27523 48280 27532
rect 48228 27489 48237 27523
rect 48237 27489 48271 27523
rect 48271 27489 48280 27523
rect 48228 27480 48280 27489
rect 20168 27455 20220 27464
rect 5908 27319 5960 27328
rect 5908 27285 5917 27319
rect 5917 27285 5951 27319
rect 5951 27285 5960 27319
rect 5908 27276 5960 27285
rect 6368 27319 6420 27328
rect 6368 27285 6377 27319
rect 6377 27285 6411 27319
rect 6411 27285 6420 27319
rect 6368 27276 6420 27285
rect 7564 27276 7616 27328
rect 13452 27319 13504 27328
rect 13452 27285 13461 27319
rect 13461 27285 13495 27319
rect 13495 27285 13504 27319
rect 13452 27276 13504 27285
rect 13544 27276 13596 27328
rect 15476 27276 15528 27328
rect 17224 27344 17276 27396
rect 15752 27276 15804 27328
rect 20168 27421 20177 27455
rect 20177 27421 20211 27455
rect 20211 27421 20220 27455
rect 20168 27412 20220 27421
rect 20812 27412 20864 27464
rect 21088 27455 21140 27464
rect 21088 27421 21097 27455
rect 21097 27421 21131 27455
rect 21131 27421 21140 27455
rect 21088 27412 21140 27421
rect 21456 27412 21508 27464
rect 26424 27455 26476 27464
rect 24860 27387 24912 27396
rect 24860 27353 24894 27387
rect 24894 27353 24912 27387
rect 24860 27344 24912 27353
rect 26424 27421 26433 27455
rect 26433 27421 26467 27455
rect 26467 27421 26476 27455
rect 26424 27412 26476 27421
rect 28540 27412 28592 27464
rect 29276 27412 29328 27464
rect 31208 27455 31260 27464
rect 31208 27421 31217 27455
rect 31217 27421 31251 27455
rect 31251 27421 31260 27455
rect 31208 27412 31260 27421
rect 32772 27412 32824 27464
rect 33600 27455 33652 27464
rect 33600 27421 33609 27455
rect 33609 27421 33643 27455
rect 33643 27421 33652 27455
rect 33600 27412 33652 27421
rect 34888 27455 34940 27464
rect 34888 27421 34897 27455
rect 34897 27421 34931 27455
rect 34931 27421 34940 27455
rect 34888 27412 34940 27421
rect 35072 27455 35124 27464
rect 35072 27421 35081 27455
rect 35081 27421 35115 27455
rect 35115 27421 35124 27455
rect 35072 27412 35124 27421
rect 35716 27455 35768 27464
rect 35716 27421 35725 27455
rect 35725 27421 35759 27455
rect 35759 27421 35768 27455
rect 35716 27412 35768 27421
rect 36176 27412 36228 27464
rect 38108 27455 38160 27464
rect 38108 27421 38117 27455
rect 38117 27421 38151 27455
rect 38151 27421 38160 27455
rect 38108 27412 38160 27421
rect 26240 27344 26292 27396
rect 27160 27344 27212 27396
rect 31300 27344 31352 27396
rect 36452 27344 36504 27396
rect 38568 27344 38620 27396
rect 47860 27344 47912 27396
rect 25044 27276 25096 27328
rect 28724 27319 28776 27328
rect 28724 27285 28733 27319
rect 28733 27285 28767 27319
rect 28767 27285 28776 27319
rect 28724 27276 28776 27285
rect 32128 27276 32180 27328
rect 33508 27276 33560 27328
rect 35808 27319 35860 27328
rect 35808 27285 35817 27319
rect 35817 27285 35851 27319
rect 35851 27285 35860 27319
rect 35808 27276 35860 27285
rect 39488 27319 39540 27328
rect 39488 27285 39497 27319
rect 39497 27285 39531 27319
rect 39531 27285 39540 27319
rect 39488 27276 39540 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 5724 27115 5776 27124
rect 5724 27081 5733 27115
rect 5733 27081 5767 27115
rect 5767 27081 5776 27115
rect 5724 27072 5776 27081
rect 9404 27115 9456 27124
rect 6368 27004 6420 27056
rect 9404 27081 9413 27115
rect 9413 27081 9447 27115
rect 9447 27081 9456 27115
rect 9404 27072 9456 27081
rect 12532 27115 12584 27124
rect 12532 27081 12541 27115
rect 12541 27081 12575 27115
rect 12575 27081 12584 27115
rect 12532 27072 12584 27081
rect 14648 27072 14700 27124
rect 15660 27072 15712 27124
rect 16856 27072 16908 27124
rect 18604 27072 18656 27124
rect 24584 27072 24636 27124
rect 28632 27072 28684 27124
rect 32128 27072 32180 27124
rect 34888 27072 34940 27124
rect 5172 26936 5224 26988
rect 5908 26936 5960 26988
rect 7564 26979 7616 26988
rect 7564 26945 7573 26979
rect 7573 26945 7607 26979
rect 7607 26945 7616 26979
rect 7564 26936 7616 26945
rect 12716 26979 12768 26988
rect 12716 26945 12725 26979
rect 12725 26945 12759 26979
rect 12759 26945 12768 26979
rect 12716 26936 12768 26945
rect 13544 26979 13596 26988
rect 13544 26945 13553 26979
rect 13553 26945 13587 26979
rect 13587 26945 13596 26979
rect 13544 26936 13596 26945
rect 16580 26936 16632 26988
rect 17224 26979 17276 26988
rect 17224 26945 17233 26979
rect 17233 26945 17267 26979
rect 17267 26945 17276 26979
rect 17224 26936 17276 26945
rect 20536 26979 20588 26988
rect 20536 26945 20545 26979
rect 20545 26945 20579 26979
rect 20579 26945 20588 26979
rect 20536 26936 20588 26945
rect 20720 26979 20772 26988
rect 20720 26945 20729 26979
rect 20729 26945 20763 26979
rect 20763 26945 20772 26979
rect 20720 26936 20772 26945
rect 22468 26979 22520 26988
rect 22468 26945 22477 26979
rect 22477 26945 22511 26979
rect 22511 26945 22520 26979
rect 22468 26936 22520 26945
rect 7104 26868 7156 26920
rect 8024 26911 8076 26920
rect 8024 26877 8033 26911
rect 8033 26877 8067 26911
rect 8067 26877 8076 26911
rect 8024 26868 8076 26877
rect 14188 26911 14240 26920
rect 14188 26877 14197 26911
rect 14197 26877 14231 26911
rect 14231 26877 14240 26911
rect 14188 26868 14240 26877
rect 15568 26868 15620 26920
rect 22560 26868 22612 26920
rect 24676 26936 24728 26988
rect 25228 27004 25280 27056
rect 26700 27004 26752 27056
rect 28724 27004 28776 27056
rect 29460 27004 29512 27056
rect 35716 27072 35768 27124
rect 38568 27115 38620 27124
rect 38568 27081 38577 27115
rect 38577 27081 38611 27115
rect 38611 27081 38620 27115
rect 38568 27072 38620 27081
rect 25044 26979 25096 26988
rect 25044 26945 25053 26979
rect 25053 26945 25087 26979
rect 25087 26945 25096 26979
rect 25044 26936 25096 26945
rect 25872 26979 25924 26988
rect 25872 26945 25881 26979
rect 25881 26945 25915 26979
rect 25915 26945 25924 26979
rect 25872 26936 25924 26945
rect 27160 26979 27212 26988
rect 24952 26868 25004 26920
rect 25596 26868 25648 26920
rect 27160 26945 27169 26979
rect 27169 26945 27203 26979
rect 27203 26945 27212 26979
rect 27160 26936 27212 26945
rect 27252 26936 27304 26988
rect 31208 26936 31260 26988
rect 31576 26979 31628 26988
rect 31576 26945 31585 26979
rect 31585 26945 31619 26979
rect 31619 26945 31628 26979
rect 31576 26936 31628 26945
rect 31760 26979 31812 26988
rect 31760 26945 31769 26979
rect 31769 26945 31803 26979
rect 31803 26945 31812 26979
rect 33508 26979 33560 26988
rect 31760 26936 31812 26945
rect 33508 26945 33542 26979
rect 33542 26945 33560 26979
rect 33508 26936 33560 26945
rect 32404 26868 32456 26920
rect 32772 26868 32824 26920
rect 23664 26800 23716 26852
rect 34612 26936 34664 26988
rect 35072 26979 35124 26988
rect 35072 26945 35081 26979
rect 35081 26945 35115 26979
rect 35115 26945 35124 26979
rect 35072 26936 35124 26945
rect 37648 26979 37700 26988
rect 37648 26945 37657 26979
rect 37657 26945 37691 26979
rect 37691 26945 37700 26979
rect 37648 26936 37700 26945
rect 38384 27004 38436 27056
rect 38016 26936 38068 26988
rect 38936 26936 38988 26988
rect 39488 26936 39540 26988
rect 6552 26775 6604 26784
rect 6552 26741 6561 26775
rect 6561 26741 6595 26775
rect 6595 26741 6604 26775
rect 6552 26732 6604 26741
rect 20352 26775 20404 26784
rect 20352 26741 20361 26775
rect 20361 26741 20395 26775
rect 20395 26741 20404 26775
rect 20352 26732 20404 26741
rect 22284 26775 22336 26784
rect 22284 26741 22293 26775
rect 22293 26741 22327 26775
rect 22327 26741 22336 26775
rect 22284 26732 22336 26741
rect 24584 26732 24636 26784
rect 24768 26732 24820 26784
rect 25136 26732 25188 26784
rect 25780 26732 25832 26784
rect 28908 26732 28960 26784
rect 29184 26732 29236 26784
rect 31484 26732 31536 26784
rect 34612 26775 34664 26784
rect 34612 26741 34621 26775
rect 34621 26741 34655 26775
rect 34655 26741 34664 26775
rect 34612 26732 34664 26741
rect 36176 26732 36228 26784
rect 38844 26732 38896 26784
rect 46480 26732 46532 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 8392 26528 8444 26580
rect 14188 26528 14240 26580
rect 17224 26528 17276 26580
rect 6920 26460 6972 26512
rect 18052 26460 18104 26512
rect 5264 26367 5316 26376
rect 5264 26333 5273 26367
rect 5273 26333 5307 26367
rect 5307 26333 5316 26367
rect 5264 26324 5316 26333
rect 6552 26324 6604 26376
rect 7104 26367 7156 26376
rect 7104 26333 7113 26367
rect 7113 26333 7147 26367
rect 7147 26333 7156 26367
rect 7104 26324 7156 26333
rect 13452 26367 13504 26376
rect 13452 26333 13461 26367
rect 13461 26333 13495 26367
rect 13495 26333 13504 26367
rect 13452 26324 13504 26333
rect 13636 26367 13688 26376
rect 13636 26333 13645 26367
rect 13645 26333 13679 26367
rect 13679 26333 13688 26367
rect 13636 26324 13688 26333
rect 7748 26256 7800 26308
rect 17408 26324 17460 26376
rect 18604 26367 18656 26376
rect 18604 26333 18613 26367
rect 18613 26333 18647 26367
rect 18647 26333 18656 26367
rect 18604 26324 18656 26333
rect 20720 26528 20772 26580
rect 21088 26571 21140 26580
rect 21088 26537 21097 26571
rect 21097 26537 21131 26571
rect 21131 26537 21140 26571
rect 21088 26528 21140 26537
rect 22652 26528 22704 26580
rect 23112 26528 23164 26580
rect 25136 26528 25188 26580
rect 25504 26528 25556 26580
rect 30380 26528 30432 26580
rect 25688 26503 25740 26512
rect 25688 26469 25697 26503
rect 25697 26469 25731 26503
rect 25731 26469 25740 26503
rect 25688 26460 25740 26469
rect 26332 26460 26384 26512
rect 28540 26503 28592 26512
rect 19432 26392 19484 26444
rect 20352 26324 20404 26376
rect 26240 26392 26292 26444
rect 28540 26469 28549 26503
rect 28549 26469 28583 26503
rect 28583 26469 28592 26503
rect 28540 26460 28592 26469
rect 31944 26460 31996 26512
rect 32772 26435 32824 26444
rect 24676 26367 24728 26376
rect 14832 26188 14884 26240
rect 17868 26256 17920 26308
rect 18512 26256 18564 26308
rect 20628 26256 20680 26308
rect 24676 26333 24685 26367
rect 24685 26333 24719 26367
rect 24719 26333 24728 26367
rect 24676 26324 24728 26333
rect 25596 26324 25648 26376
rect 25688 26324 25740 26376
rect 32772 26401 32781 26435
rect 32781 26401 32815 26435
rect 32815 26401 32824 26435
rect 32772 26392 32824 26401
rect 22284 26299 22336 26308
rect 22284 26265 22318 26299
rect 22318 26265 22336 26299
rect 22284 26256 22336 26265
rect 19984 26188 20036 26240
rect 25136 26256 25188 26308
rect 25044 26188 25096 26240
rect 27068 26256 27120 26308
rect 28632 26324 28684 26376
rect 28724 26367 28776 26376
rect 28724 26333 28733 26367
rect 28733 26333 28767 26367
rect 28767 26333 28776 26367
rect 28724 26324 28776 26333
rect 28908 26324 28960 26376
rect 29184 26367 29236 26376
rect 29184 26333 29193 26367
rect 29193 26333 29227 26367
rect 29227 26333 29236 26367
rect 29184 26324 29236 26333
rect 30748 26324 30800 26376
rect 31944 26367 31996 26376
rect 31944 26333 31953 26367
rect 31953 26333 31987 26367
rect 31987 26333 31996 26367
rect 31944 26324 31996 26333
rect 35900 26460 35952 26512
rect 38844 26460 38896 26512
rect 35716 26392 35768 26444
rect 46480 26435 46532 26444
rect 35808 26324 35860 26376
rect 36084 26324 36136 26376
rect 36544 26367 36596 26376
rect 36544 26333 36553 26367
rect 36553 26333 36587 26367
rect 36587 26333 36596 26367
rect 36544 26324 36596 26333
rect 37648 26324 37700 26376
rect 38292 26324 38344 26376
rect 38384 26367 38436 26376
rect 38384 26333 38393 26367
rect 38393 26333 38427 26367
rect 38427 26333 38436 26367
rect 38384 26324 38436 26333
rect 38568 26367 38620 26376
rect 38568 26333 38577 26367
rect 38577 26333 38611 26367
rect 38611 26333 38620 26367
rect 46480 26401 46489 26435
rect 46489 26401 46523 26435
rect 46523 26401 46532 26435
rect 46480 26392 46532 26401
rect 48228 26435 48280 26444
rect 48228 26401 48237 26435
rect 48237 26401 48271 26435
rect 48271 26401 48280 26435
rect 48228 26392 48280 26401
rect 38568 26324 38620 26333
rect 40684 26324 40736 26376
rect 29736 26299 29788 26308
rect 29736 26265 29745 26299
rect 29745 26265 29779 26299
rect 29779 26265 29788 26299
rect 29736 26256 29788 26265
rect 33784 26256 33836 26308
rect 35992 26256 36044 26308
rect 47860 26256 47912 26308
rect 27344 26188 27396 26240
rect 35440 26231 35492 26240
rect 35440 26197 35449 26231
rect 35449 26197 35483 26231
rect 35483 26197 35492 26231
rect 35440 26188 35492 26197
rect 39028 26231 39080 26240
rect 39028 26197 39037 26231
rect 39037 26197 39071 26231
rect 39071 26197 39080 26231
rect 39028 26188 39080 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 7748 26027 7800 26036
rect 7748 25993 7757 26027
rect 7757 25993 7791 26027
rect 7791 25993 7800 26027
rect 7748 25984 7800 25993
rect 17868 26027 17920 26036
rect 17868 25993 17877 26027
rect 17877 25993 17911 26027
rect 17911 25993 17920 26027
rect 17868 25984 17920 25993
rect 20536 26027 20588 26036
rect 20536 25993 20545 26027
rect 20545 25993 20579 26027
rect 20579 25993 20588 26027
rect 20536 25984 20588 25993
rect 22468 26027 22520 26036
rect 22468 25993 22477 26027
rect 22477 25993 22511 26027
rect 22511 25993 22520 26027
rect 22468 25984 22520 25993
rect 12900 25916 12952 25968
rect 25688 25984 25740 26036
rect 26424 25984 26476 26036
rect 27252 25984 27304 26036
rect 31300 26027 31352 26036
rect 31300 25993 31309 26027
rect 31309 25993 31343 26027
rect 31343 25993 31352 26027
rect 31300 25984 31352 25993
rect 33600 25984 33652 26036
rect 35440 25984 35492 26036
rect 40684 26027 40736 26036
rect 40684 25993 40693 26027
rect 40693 25993 40727 26027
rect 40727 25993 40736 26027
rect 40684 25984 40736 25993
rect 47860 26027 47912 26036
rect 47860 25993 47869 26027
rect 47869 25993 47903 26027
rect 47903 25993 47912 26027
rect 47860 25984 47912 25993
rect 2228 25891 2280 25900
rect 2228 25857 2237 25891
rect 2237 25857 2271 25891
rect 2271 25857 2280 25891
rect 2228 25848 2280 25857
rect 7012 25848 7064 25900
rect 12808 25848 12860 25900
rect 13636 25848 13688 25900
rect 16580 25848 16632 25900
rect 17040 25848 17092 25900
rect 18052 25891 18104 25900
rect 18052 25857 18061 25891
rect 18061 25857 18095 25891
rect 18095 25857 18104 25891
rect 18052 25848 18104 25857
rect 1768 25644 1820 25696
rect 6920 25687 6972 25696
rect 6920 25653 6929 25687
rect 6929 25653 6963 25687
rect 6963 25653 6972 25687
rect 6920 25644 6972 25653
rect 12532 25687 12584 25696
rect 12532 25653 12541 25687
rect 12541 25653 12575 25687
rect 12575 25653 12584 25687
rect 12532 25644 12584 25653
rect 16856 25644 16908 25696
rect 17040 25644 17092 25696
rect 18236 25687 18288 25696
rect 18236 25653 18245 25687
rect 18245 25653 18279 25687
rect 18279 25653 18288 25687
rect 18236 25644 18288 25653
rect 21088 25848 21140 25900
rect 21916 25848 21968 25900
rect 23756 25916 23808 25968
rect 24676 25916 24728 25968
rect 25872 25959 25924 25968
rect 25872 25925 25881 25959
rect 25881 25925 25915 25959
rect 25915 25925 25924 25959
rect 25872 25916 25924 25925
rect 32496 25916 32548 25968
rect 36084 25916 36136 25968
rect 36176 25959 36228 25968
rect 36176 25925 36201 25959
rect 36201 25925 36228 25959
rect 36176 25916 36228 25925
rect 39028 25916 39080 25968
rect 23112 25891 23164 25900
rect 23112 25857 23121 25891
rect 23121 25857 23155 25891
rect 23155 25857 23164 25891
rect 23112 25848 23164 25857
rect 25688 25891 25740 25900
rect 25688 25857 25697 25891
rect 25697 25857 25731 25891
rect 25731 25857 25740 25891
rect 25688 25848 25740 25857
rect 27344 25891 27396 25900
rect 27344 25857 27353 25891
rect 27353 25857 27387 25891
rect 27387 25857 27396 25891
rect 27344 25848 27396 25857
rect 23664 25780 23716 25832
rect 27896 25848 27948 25900
rect 28356 25848 28408 25900
rect 31484 25891 31536 25900
rect 27988 25780 28040 25832
rect 29276 25780 29328 25832
rect 31484 25857 31493 25891
rect 31493 25857 31527 25891
rect 31527 25857 31536 25891
rect 31484 25848 31536 25857
rect 32128 25848 32180 25900
rect 32220 25848 32272 25900
rect 34612 25848 34664 25900
rect 38292 25891 38344 25900
rect 25044 25712 25096 25764
rect 30196 25712 30248 25764
rect 34244 25780 34296 25832
rect 35440 25780 35492 25832
rect 22468 25644 22520 25696
rect 27528 25687 27580 25696
rect 27528 25653 27537 25687
rect 27537 25653 27571 25687
rect 27571 25653 27580 25687
rect 27528 25644 27580 25653
rect 30472 25644 30524 25696
rect 33508 25712 33560 25764
rect 32404 25644 32456 25696
rect 38292 25857 38301 25891
rect 38301 25857 38335 25891
rect 38335 25857 38344 25891
rect 38292 25848 38344 25857
rect 38384 25848 38436 25900
rect 38568 25891 38620 25900
rect 38568 25857 38577 25891
rect 38577 25857 38611 25891
rect 38611 25857 38620 25891
rect 38568 25848 38620 25857
rect 38752 25891 38804 25900
rect 38752 25857 38761 25891
rect 38761 25857 38795 25891
rect 38795 25857 38804 25891
rect 38752 25848 38804 25857
rect 47768 25891 47820 25900
rect 47768 25857 47777 25891
rect 47777 25857 47811 25891
rect 47811 25857 47820 25891
rect 47768 25848 47820 25857
rect 37280 25780 37332 25832
rect 38108 25780 38160 25832
rect 36544 25712 36596 25764
rect 36728 25712 36780 25764
rect 36912 25644 36964 25696
rect 38200 25644 38252 25696
rect 46480 25644 46532 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 13636 25440 13688 25492
rect 16580 25440 16632 25492
rect 17316 25440 17368 25492
rect 18788 25483 18840 25492
rect 18788 25449 18797 25483
rect 18797 25449 18831 25483
rect 18831 25449 18840 25483
rect 18788 25440 18840 25449
rect 20812 25440 20864 25492
rect 21916 25440 21968 25492
rect 24952 25440 25004 25492
rect 32496 25483 32548 25492
rect 32496 25449 32505 25483
rect 32505 25449 32539 25483
rect 32539 25449 32548 25483
rect 32496 25440 32548 25449
rect 18236 25372 18288 25424
rect 27528 25372 27580 25424
rect 31024 25372 31076 25424
rect 1768 25347 1820 25356
rect 1768 25313 1777 25347
rect 1777 25313 1811 25347
rect 1811 25313 1820 25347
rect 1768 25304 1820 25313
rect 2780 25347 2832 25356
rect 2780 25313 2789 25347
rect 2789 25313 2823 25347
rect 2823 25313 2832 25347
rect 2780 25304 2832 25313
rect 11980 25304 12032 25356
rect 1584 25279 1636 25288
rect 1584 25245 1593 25279
rect 1593 25245 1627 25279
rect 1627 25245 1636 25279
rect 1584 25236 1636 25245
rect 19340 25304 19392 25356
rect 23664 25347 23716 25356
rect 13820 25236 13872 25288
rect 14832 25279 14884 25288
rect 14832 25245 14841 25279
rect 14841 25245 14875 25279
rect 14875 25245 14884 25279
rect 14832 25236 14884 25245
rect 16856 25279 16908 25288
rect 16856 25245 16865 25279
rect 16865 25245 16899 25279
rect 16899 25245 16908 25279
rect 16856 25236 16908 25245
rect 17040 25279 17092 25288
rect 17040 25245 17049 25279
rect 17049 25245 17083 25279
rect 17083 25245 17092 25279
rect 17040 25236 17092 25245
rect 17592 25236 17644 25288
rect 12348 25211 12400 25220
rect 12348 25177 12382 25211
rect 12382 25177 12400 25211
rect 12348 25168 12400 25177
rect 19248 25236 19300 25288
rect 19984 25236 20036 25288
rect 23664 25313 23673 25347
rect 23673 25313 23707 25347
rect 23707 25313 23716 25347
rect 23664 25304 23716 25313
rect 21364 25236 21416 25288
rect 20812 25168 20864 25220
rect 22376 25236 22428 25288
rect 29368 25304 29420 25356
rect 25688 25236 25740 25288
rect 27712 25279 27764 25288
rect 27712 25245 27721 25279
rect 27721 25245 27755 25279
rect 27755 25245 27764 25279
rect 27712 25236 27764 25245
rect 28356 25236 28408 25288
rect 30104 25279 30156 25288
rect 30104 25245 30113 25279
rect 30113 25245 30147 25279
rect 30147 25245 30156 25279
rect 30104 25236 30156 25245
rect 30196 25236 30248 25288
rect 30840 25236 30892 25288
rect 33784 25236 33836 25288
rect 36176 25304 36228 25356
rect 36452 25347 36504 25356
rect 36452 25313 36461 25347
rect 36461 25313 36495 25347
rect 36495 25313 36504 25347
rect 36452 25304 36504 25313
rect 46480 25347 46532 25356
rect 46480 25313 46489 25347
rect 46489 25313 46523 25347
rect 46523 25313 46532 25347
rect 46480 25304 46532 25313
rect 48228 25347 48280 25356
rect 48228 25313 48237 25347
rect 48237 25313 48271 25347
rect 48271 25313 48280 25347
rect 48228 25304 48280 25313
rect 36360 25279 36412 25288
rect 18420 25143 18472 25152
rect 18420 25109 18429 25143
rect 18429 25109 18463 25143
rect 18463 25109 18472 25143
rect 18420 25100 18472 25109
rect 18788 25100 18840 25152
rect 23664 25168 23716 25220
rect 24584 25168 24636 25220
rect 31392 25211 31444 25220
rect 31392 25177 31426 25211
rect 31426 25177 31444 25211
rect 36360 25245 36369 25279
rect 36369 25245 36403 25279
rect 36403 25245 36412 25279
rect 36360 25236 36412 25245
rect 36912 25279 36964 25288
rect 36912 25245 36921 25279
rect 36921 25245 36955 25279
rect 36955 25245 36964 25279
rect 36912 25236 36964 25245
rect 37280 25236 37332 25288
rect 31392 25168 31444 25177
rect 36452 25168 36504 25220
rect 21640 25143 21692 25152
rect 21640 25109 21649 25143
rect 21649 25109 21683 25143
rect 21683 25109 21692 25143
rect 21640 25100 21692 25109
rect 27896 25143 27948 25152
rect 27896 25109 27905 25143
rect 27905 25109 27939 25143
rect 27939 25109 27948 25143
rect 27896 25100 27948 25109
rect 28724 25100 28776 25152
rect 29920 25143 29972 25152
rect 29920 25109 29929 25143
rect 29929 25109 29963 25143
rect 29963 25109 29972 25143
rect 29920 25100 29972 25109
rect 34152 25100 34204 25152
rect 38016 25168 38068 25220
rect 47124 25168 47176 25220
rect 38476 25100 38528 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 12348 24939 12400 24948
rect 12348 24905 12357 24939
rect 12357 24905 12391 24939
rect 12391 24905 12400 24939
rect 12348 24896 12400 24905
rect 17592 24896 17644 24948
rect 18420 24871 18472 24880
rect 1584 24760 1636 24812
rect 12532 24803 12584 24812
rect 12532 24769 12541 24803
rect 12541 24769 12575 24803
rect 12575 24769 12584 24803
rect 12532 24760 12584 24769
rect 13820 24803 13872 24812
rect 13820 24769 13829 24803
rect 13829 24769 13863 24803
rect 13863 24769 13872 24803
rect 13820 24760 13872 24769
rect 14372 24760 14424 24812
rect 15844 24803 15896 24812
rect 15844 24769 15853 24803
rect 15853 24769 15887 24803
rect 15887 24769 15896 24803
rect 15844 24760 15896 24769
rect 18420 24837 18454 24871
rect 18454 24837 18472 24871
rect 18420 24828 18472 24837
rect 19340 24896 19392 24948
rect 21640 24896 21692 24948
rect 12808 24735 12860 24744
rect 12808 24701 12817 24735
rect 12817 24701 12851 24735
rect 12851 24701 12860 24735
rect 12808 24692 12860 24701
rect 19984 24760 20036 24812
rect 20260 24760 20312 24812
rect 22100 24760 22152 24812
rect 22376 24803 22428 24812
rect 18144 24735 18196 24744
rect 18144 24701 18153 24735
rect 18153 24701 18187 24735
rect 18187 24701 18196 24735
rect 18144 24692 18196 24701
rect 15292 24624 15344 24676
rect 17040 24624 17092 24676
rect 22376 24769 22385 24803
rect 22385 24769 22419 24803
rect 22419 24769 22428 24803
rect 22376 24760 22428 24769
rect 23112 24803 23164 24812
rect 23112 24769 23121 24803
rect 23121 24769 23155 24803
rect 23155 24769 23164 24803
rect 23112 24760 23164 24769
rect 23204 24760 23256 24812
rect 23756 24803 23808 24812
rect 23756 24769 23765 24803
rect 23765 24769 23799 24803
rect 23799 24769 23808 24803
rect 23756 24760 23808 24769
rect 22468 24735 22520 24744
rect 22468 24701 22477 24735
rect 22477 24701 22511 24735
rect 22511 24701 22520 24735
rect 24216 24760 24268 24812
rect 25688 24760 25740 24812
rect 25872 24760 25924 24812
rect 24400 24735 24452 24744
rect 22468 24692 22520 24701
rect 24400 24701 24409 24735
rect 24409 24701 24443 24735
rect 24443 24701 24452 24735
rect 24400 24692 24452 24701
rect 15660 24599 15712 24608
rect 15660 24565 15669 24599
rect 15669 24565 15703 24599
rect 15703 24565 15712 24599
rect 15660 24556 15712 24565
rect 22008 24599 22060 24608
rect 22008 24565 22017 24599
rect 22017 24565 22051 24599
rect 22051 24565 22060 24599
rect 22008 24556 22060 24565
rect 23388 24556 23440 24608
rect 24768 24624 24820 24676
rect 24676 24599 24728 24608
rect 24676 24565 24685 24599
rect 24685 24565 24719 24599
rect 24719 24565 24728 24599
rect 24676 24556 24728 24565
rect 29644 24896 29696 24948
rect 29920 24828 29972 24880
rect 27528 24760 27580 24812
rect 27620 24803 27672 24812
rect 27620 24769 27629 24803
rect 27629 24769 27663 24803
rect 27663 24769 27672 24803
rect 27620 24760 27672 24769
rect 30656 24760 30708 24812
rect 29460 24735 29512 24744
rect 29460 24701 29469 24735
rect 29469 24701 29503 24735
rect 29503 24701 29512 24735
rect 29460 24692 29512 24701
rect 31392 24896 31444 24948
rect 32496 24896 32548 24948
rect 38016 24939 38068 24948
rect 38016 24905 38025 24939
rect 38025 24905 38059 24939
rect 38059 24905 38068 24939
rect 38016 24896 38068 24905
rect 32772 24803 32824 24812
rect 31668 24735 31720 24744
rect 31668 24701 31677 24735
rect 31677 24701 31711 24735
rect 31711 24701 31720 24735
rect 31668 24692 31720 24701
rect 31760 24735 31812 24744
rect 31760 24701 31769 24735
rect 31769 24701 31803 24735
rect 31803 24701 31812 24735
rect 32772 24769 32781 24803
rect 32781 24769 32815 24803
rect 32815 24769 32824 24803
rect 32772 24760 32824 24769
rect 33140 24760 33192 24812
rect 36360 24828 36412 24880
rect 37372 24828 37424 24880
rect 47400 24828 47452 24880
rect 47768 24828 47820 24880
rect 33876 24803 33928 24812
rect 33876 24769 33885 24803
rect 33885 24769 33919 24803
rect 33919 24769 33928 24803
rect 33876 24760 33928 24769
rect 34060 24803 34112 24812
rect 34060 24769 34069 24803
rect 34069 24769 34103 24803
rect 34103 24769 34112 24803
rect 34060 24760 34112 24769
rect 35716 24760 35768 24812
rect 35992 24803 36044 24812
rect 35992 24769 36001 24803
rect 36001 24769 36035 24803
rect 36035 24769 36044 24803
rect 35992 24760 36044 24769
rect 36452 24760 36504 24812
rect 36728 24803 36780 24812
rect 36728 24769 36737 24803
rect 36737 24769 36771 24803
rect 36771 24769 36780 24803
rect 36728 24760 36780 24769
rect 38200 24803 38252 24812
rect 31760 24692 31812 24701
rect 33968 24692 34020 24744
rect 36084 24692 36136 24744
rect 38200 24769 38209 24803
rect 38209 24769 38243 24803
rect 38243 24769 38252 24803
rect 38200 24760 38252 24769
rect 47032 24803 47084 24812
rect 47032 24769 47041 24803
rect 47041 24769 47075 24803
rect 47075 24769 47084 24803
rect 47032 24760 47084 24769
rect 47124 24803 47176 24812
rect 47124 24769 47133 24803
rect 47133 24769 47167 24803
rect 47167 24769 47176 24803
rect 47124 24760 47176 24769
rect 48228 24760 48280 24812
rect 38476 24735 38528 24744
rect 38476 24701 38485 24735
rect 38485 24701 38519 24735
rect 38519 24701 38528 24735
rect 38476 24692 38528 24701
rect 26240 24556 26292 24608
rect 27160 24599 27212 24608
rect 27160 24565 27169 24599
rect 27169 24565 27203 24599
rect 27203 24565 27212 24599
rect 27160 24556 27212 24565
rect 29644 24556 29696 24608
rect 29736 24556 29788 24608
rect 46848 24624 46900 24676
rect 30840 24599 30892 24608
rect 30840 24565 30849 24599
rect 30849 24565 30883 24599
rect 30883 24565 30892 24599
rect 30840 24556 30892 24565
rect 32772 24556 32824 24608
rect 36360 24556 36412 24608
rect 38384 24599 38436 24608
rect 38384 24565 38393 24599
rect 38393 24565 38427 24599
rect 38427 24565 38436 24599
rect 38384 24556 38436 24565
rect 38844 24556 38896 24608
rect 46940 24556 46992 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 14372 24395 14424 24404
rect 14372 24361 14381 24395
rect 14381 24361 14415 24395
rect 14415 24361 14424 24395
rect 14372 24352 14424 24361
rect 15844 24352 15896 24404
rect 23020 24352 23072 24404
rect 23204 24395 23256 24404
rect 23204 24361 23213 24395
rect 23213 24361 23247 24395
rect 23247 24361 23256 24395
rect 23204 24352 23256 24361
rect 23664 24395 23716 24404
rect 23664 24361 23673 24395
rect 23673 24361 23707 24395
rect 23707 24361 23716 24395
rect 23664 24352 23716 24361
rect 17316 24284 17368 24336
rect 23388 24284 23440 24336
rect 15660 24216 15712 24268
rect 22100 24216 22152 24268
rect 24492 24216 24544 24268
rect 12808 24080 12860 24132
rect 17500 24148 17552 24200
rect 19248 24148 19300 24200
rect 20628 24191 20680 24200
rect 20628 24157 20637 24191
rect 20637 24157 20671 24191
rect 20671 24157 20680 24191
rect 20628 24148 20680 24157
rect 22008 24148 22060 24200
rect 23112 24191 23164 24200
rect 23112 24157 23121 24191
rect 23121 24157 23155 24191
rect 23155 24157 23164 24191
rect 23112 24148 23164 24157
rect 23388 24191 23440 24200
rect 23388 24157 23397 24191
rect 23397 24157 23431 24191
rect 23431 24157 23440 24191
rect 23388 24148 23440 24157
rect 30104 24352 30156 24404
rect 25596 24284 25648 24336
rect 42892 24352 42944 24404
rect 26240 24216 26292 24268
rect 27160 24148 27212 24200
rect 17408 24080 17460 24132
rect 18512 24123 18564 24132
rect 18512 24089 18521 24123
rect 18521 24089 18555 24123
rect 18555 24089 18564 24123
rect 18512 24080 18564 24089
rect 20260 24080 20312 24132
rect 23480 24080 23532 24132
rect 24768 24080 24820 24132
rect 25780 24123 25832 24132
rect 16948 24055 17000 24064
rect 16948 24021 16957 24055
rect 16957 24021 16991 24055
rect 16991 24021 17000 24055
rect 16948 24012 17000 24021
rect 21364 24012 21416 24064
rect 24400 24012 24452 24064
rect 25780 24089 25789 24123
rect 25789 24089 25823 24123
rect 25823 24089 25832 24123
rect 25780 24080 25832 24089
rect 25872 24080 25924 24132
rect 34060 24284 34112 24336
rect 39764 24284 39816 24336
rect 31576 24216 31628 24268
rect 35992 24216 36044 24268
rect 30288 24191 30340 24200
rect 30288 24157 30297 24191
rect 30297 24157 30331 24191
rect 30331 24157 30340 24191
rect 30288 24148 30340 24157
rect 30748 24080 30800 24132
rect 28172 24012 28224 24064
rect 29828 24012 29880 24064
rect 33784 24148 33836 24200
rect 33876 24148 33928 24200
rect 34060 24148 34112 24200
rect 36360 24191 36412 24200
rect 36360 24157 36369 24191
rect 36369 24157 36403 24191
rect 36403 24157 36412 24191
rect 36360 24148 36412 24157
rect 37280 24216 37332 24268
rect 39396 24148 39448 24200
rect 32588 24123 32640 24132
rect 32588 24089 32622 24123
rect 32622 24089 32640 24123
rect 32588 24080 32640 24089
rect 36452 24012 36504 24064
rect 40868 24012 40920 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 17500 23851 17552 23860
rect 17500 23817 17509 23851
rect 17509 23817 17543 23851
rect 17543 23817 17552 23851
rect 17500 23808 17552 23817
rect 25044 23851 25096 23860
rect 25044 23817 25053 23851
rect 25053 23817 25087 23851
rect 25087 23817 25096 23851
rect 25044 23808 25096 23817
rect 25688 23851 25740 23860
rect 25688 23817 25697 23851
rect 25697 23817 25731 23851
rect 25731 23817 25740 23851
rect 25688 23808 25740 23817
rect 27528 23851 27580 23860
rect 27528 23817 27537 23851
rect 27537 23817 27571 23851
rect 27571 23817 27580 23851
rect 27528 23808 27580 23817
rect 11888 23783 11940 23792
rect 11888 23749 11897 23783
rect 11897 23749 11931 23783
rect 11931 23749 11940 23783
rect 11888 23740 11940 23749
rect 16856 23740 16908 23792
rect 18512 23740 18564 23792
rect 19432 23740 19484 23792
rect 20168 23740 20220 23792
rect 24400 23740 24452 23792
rect 17960 23715 18012 23724
rect 17960 23681 17969 23715
rect 17969 23681 18003 23715
rect 18003 23681 18012 23715
rect 17960 23672 18012 23681
rect 18880 23672 18932 23724
rect 21916 23672 21968 23724
rect 24216 23672 24268 23724
rect 25596 23715 25648 23724
rect 25596 23681 25605 23715
rect 25605 23681 25639 23715
rect 25639 23681 25648 23715
rect 25596 23672 25648 23681
rect 25780 23715 25832 23724
rect 25780 23681 25789 23715
rect 25789 23681 25823 23715
rect 25823 23681 25832 23715
rect 25780 23672 25832 23681
rect 29920 23740 29972 23792
rect 30748 23808 30800 23860
rect 32404 23808 32456 23860
rect 32588 23851 32640 23860
rect 32588 23817 32597 23851
rect 32597 23817 32631 23851
rect 32631 23817 32640 23851
rect 32588 23808 32640 23817
rect 39396 23851 39448 23860
rect 39396 23817 39405 23851
rect 39405 23817 39439 23851
rect 39439 23817 39448 23851
rect 39396 23808 39448 23817
rect 39764 23851 39816 23860
rect 39764 23817 39773 23851
rect 39773 23817 39807 23851
rect 39807 23817 39816 23851
rect 39764 23808 39816 23817
rect 46940 23740 46992 23792
rect 28172 23715 28224 23724
rect 18052 23536 18104 23588
rect 4068 23468 4120 23520
rect 11060 23468 11112 23520
rect 13360 23468 13412 23520
rect 21456 23468 21508 23520
rect 22284 23468 22336 23520
rect 26700 23604 26752 23656
rect 28172 23681 28181 23715
rect 28181 23681 28215 23715
rect 28215 23681 28224 23715
rect 28172 23672 28224 23681
rect 29552 23715 29604 23724
rect 29552 23681 29561 23715
rect 29561 23681 29595 23715
rect 29595 23681 29604 23715
rect 29552 23672 29604 23681
rect 29644 23672 29696 23724
rect 32772 23715 32824 23724
rect 32772 23681 32781 23715
rect 32781 23681 32815 23715
rect 32815 23681 32824 23715
rect 32772 23672 32824 23681
rect 33784 23715 33836 23724
rect 33784 23681 33793 23715
rect 33793 23681 33827 23715
rect 33827 23681 33836 23715
rect 33784 23672 33836 23681
rect 33876 23672 33928 23724
rect 36452 23715 36504 23724
rect 36452 23681 36461 23715
rect 36461 23681 36495 23715
rect 36495 23681 36504 23715
rect 36452 23672 36504 23681
rect 37372 23672 37424 23724
rect 40868 23672 40920 23724
rect 46296 23715 46348 23724
rect 46296 23681 46305 23715
rect 46305 23681 46339 23715
rect 46339 23681 46348 23715
rect 46296 23672 46348 23681
rect 29828 23647 29880 23656
rect 23020 23536 23072 23588
rect 27896 23536 27948 23588
rect 29828 23613 29837 23647
rect 29837 23613 29871 23647
rect 29871 23613 29880 23647
rect 29828 23604 29880 23613
rect 31852 23604 31904 23656
rect 39948 23647 40000 23656
rect 39948 23613 39957 23647
rect 39957 23613 39991 23647
rect 39991 23613 40000 23647
rect 40684 23647 40736 23656
rect 39948 23604 40000 23613
rect 40684 23613 40693 23647
rect 40693 23613 40727 23647
rect 40727 23613 40736 23647
rect 40684 23604 40736 23613
rect 30104 23536 30156 23588
rect 31668 23536 31720 23588
rect 33140 23536 33192 23588
rect 23388 23468 23440 23520
rect 24768 23468 24820 23520
rect 25780 23468 25832 23520
rect 28264 23468 28316 23520
rect 29460 23468 29512 23520
rect 31484 23468 31536 23520
rect 34060 23468 34112 23520
rect 35348 23468 35400 23520
rect 36544 23511 36596 23520
rect 36544 23477 36553 23511
rect 36553 23477 36587 23511
rect 36587 23477 36596 23511
rect 36544 23468 36596 23477
rect 46388 23511 46440 23520
rect 46388 23477 46397 23511
rect 46397 23477 46431 23511
rect 46431 23477 46440 23511
rect 46388 23468 46440 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 12992 23264 13044 23316
rect 18052 23307 18104 23316
rect 11060 23171 11112 23180
rect 11060 23137 11069 23171
rect 11069 23137 11103 23171
rect 11103 23137 11112 23171
rect 11060 23128 11112 23137
rect 13912 23128 13964 23180
rect 18052 23273 18061 23307
rect 18061 23273 18095 23307
rect 18095 23273 18104 23307
rect 18052 23264 18104 23273
rect 23480 23264 23532 23316
rect 24584 23264 24636 23316
rect 29552 23264 29604 23316
rect 40684 23264 40736 23316
rect 10140 23103 10192 23112
rect 10140 23069 10149 23103
rect 10149 23069 10183 23103
rect 10183 23069 10192 23103
rect 10140 23060 10192 23069
rect 14556 23103 14608 23112
rect 14556 23069 14565 23103
rect 14565 23069 14599 23103
rect 14599 23069 14608 23103
rect 14556 23060 14608 23069
rect 18144 23060 18196 23112
rect 18420 23128 18472 23180
rect 19432 23171 19484 23180
rect 19432 23137 19441 23171
rect 19441 23137 19475 23171
rect 19475 23137 19484 23171
rect 19432 23128 19484 23137
rect 18512 23103 18564 23112
rect 18512 23069 18521 23103
rect 18521 23069 18555 23103
rect 18555 23069 18564 23103
rect 18512 23060 18564 23069
rect 18880 23060 18932 23112
rect 21456 23103 21508 23112
rect 21456 23069 21465 23103
rect 21465 23069 21499 23103
rect 21499 23069 21508 23103
rect 21456 23060 21508 23069
rect 24676 23103 24728 23112
rect 24676 23069 24685 23103
rect 24685 23069 24719 23103
rect 24719 23069 24728 23103
rect 24676 23060 24728 23069
rect 26240 23060 26292 23112
rect 27712 23060 27764 23112
rect 29920 23103 29972 23112
rect 29920 23069 29929 23103
rect 29929 23069 29963 23103
rect 29963 23069 29972 23103
rect 29920 23060 29972 23069
rect 30104 23060 30156 23112
rect 10508 22992 10560 23044
rect 16948 22992 17000 23044
rect 17316 22924 17368 22976
rect 20536 22924 20588 22976
rect 22652 22992 22704 23044
rect 23388 22992 23440 23044
rect 30564 23060 30616 23112
rect 40040 23128 40092 23180
rect 47584 23171 47636 23180
rect 47584 23137 47593 23171
rect 47593 23137 47627 23171
rect 47627 23137 47636 23171
rect 47584 23128 47636 23137
rect 33968 23060 34020 23112
rect 34060 23060 34112 23112
rect 35348 23060 35400 23112
rect 36268 23060 36320 23112
rect 36544 23103 36596 23112
rect 36544 23069 36553 23103
rect 36553 23069 36587 23103
rect 36587 23069 36596 23103
rect 36544 23060 36596 23069
rect 39120 23103 39172 23112
rect 39120 23069 39129 23103
rect 39129 23069 39163 23103
rect 39163 23069 39172 23103
rect 39120 23060 39172 23069
rect 31484 22992 31536 23044
rect 36452 22992 36504 23044
rect 39396 23103 39448 23112
rect 39396 23069 39405 23103
rect 39405 23069 39439 23103
rect 39439 23069 39448 23103
rect 39396 23060 39448 23069
rect 40316 23060 40368 23112
rect 22928 22967 22980 22976
rect 22928 22933 22937 22967
rect 22937 22933 22971 22967
rect 22971 22933 22980 22967
rect 22928 22924 22980 22933
rect 27712 22924 27764 22976
rect 31852 22924 31904 22976
rect 33692 22967 33744 22976
rect 33692 22933 33701 22967
rect 33701 22933 33735 22967
rect 33735 22933 33744 22967
rect 33692 22924 33744 22933
rect 35808 22924 35860 22976
rect 39580 22992 39632 23044
rect 40592 23060 40644 23112
rect 45928 23103 45980 23112
rect 45928 23069 45937 23103
rect 45937 23069 45971 23103
rect 45971 23069 45980 23103
rect 45928 23060 45980 23069
rect 46112 23035 46164 23044
rect 46112 23001 46121 23035
rect 46121 23001 46155 23035
rect 46155 23001 46164 23035
rect 46112 22992 46164 23001
rect 37372 22924 37424 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 10508 22763 10560 22772
rect 10508 22729 10517 22763
rect 10517 22729 10551 22763
rect 10551 22729 10560 22763
rect 10508 22720 10560 22729
rect 18972 22720 19024 22772
rect 20168 22763 20220 22772
rect 20168 22729 20177 22763
rect 20177 22729 20211 22763
rect 20211 22729 20220 22763
rect 20168 22720 20220 22729
rect 20536 22763 20588 22772
rect 20536 22729 20545 22763
rect 20545 22729 20579 22763
rect 20579 22729 20588 22763
rect 20536 22720 20588 22729
rect 27712 22720 27764 22772
rect 10416 22627 10468 22636
rect 10416 22593 10425 22627
rect 10425 22593 10459 22627
rect 10459 22593 10468 22627
rect 10416 22584 10468 22593
rect 12164 22516 12216 22568
rect 12532 22627 12584 22636
rect 12532 22593 12566 22627
rect 12566 22593 12584 22627
rect 14556 22652 14608 22704
rect 16856 22695 16908 22704
rect 16856 22661 16865 22695
rect 16865 22661 16899 22695
rect 16899 22661 16908 22695
rect 16856 22652 16908 22661
rect 12532 22584 12584 22593
rect 14280 22584 14332 22636
rect 18788 22584 18840 22636
rect 22928 22652 22980 22704
rect 31760 22720 31812 22772
rect 33876 22720 33928 22772
rect 23480 22627 23532 22636
rect 23480 22593 23489 22627
rect 23489 22593 23523 22627
rect 23523 22593 23532 22627
rect 23480 22584 23532 22593
rect 18420 22559 18472 22568
rect 18420 22525 18429 22559
rect 18429 22525 18463 22559
rect 18463 22525 18472 22559
rect 18420 22516 18472 22525
rect 19340 22516 19392 22568
rect 21732 22516 21784 22568
rect 22652 22516 22704 22568
rect 23204 22516 23256 22568
rect 29000 22584 29052 22636
rect 29368 22652 29420 22704
rect 30840 22652 30892 22704
rect 29460 22627 29512 22636
rect 29460 22593 29494 22627
rect 29494 22593 29512 22627
rect 29460 22584 29512 22593
rect 33508 22652 33560 22704
rect 38752 22720 38804 22772
rect 39672 22720 39724 22772
rect 40040 22720 40092 22772
rect 40868 22720 40920 22772
rect 46112 22763 46164 22772
rect 46112 22729 46121 22763
rect 46121 22729 46155 22763
rect 46155 22729 46164 22763
rect 46112 22720 46164 22729
rect 31852 22516 31904 22568
rect 33692 22584 33744 22636
rect 35348 22652 35400 22704
rect 35808 22627 35860 22636
rect 35808 22593 35817 22627
rect 35817 22593 35851 22627
rect 35851 22593 35860 22627
rect 35808 22584 35860 22593
rect 35900 22584 35952 22636
rect 39120 22652 39172 22704
rect 38476 22627 38528 22636
rect 38476 22593 38485 22627
rect 38485 22593 38519 22627
rect 38519 22593 38528 22627
rect 38476 22584 38528 22593
rect 38936 22584 38988 22636
rect 39304 22627 39356 22636
rect 39304 22593 39313 22627
rect 39313 22593 39347 22627
rect 39347 22593 39356 22627
rect 39304 22584 39356 22593
rect 39580 22627 39632 22636
rect 39580 22593 39589 22627
rect 39589 22593 39623 22627
rect 39623 22593 39632 22627
rect 39580 22584 39632 22593
rect 40040 22584 40092 22636
rect 33140 22516 33192 22568
rect 36084 22559 36136 22568
rect 36084 22525 36093 22559
rect 36093 22525 36127 22559
rect 36127 22525 36136 22559
rect 36084 22516 36136 22525
rect 36176 22559 36228 22568
rect 36176 22525 36185 22559
rect 36185 22525 36219 22559
rect 36219 22525 36228 22559
rect 36176 22516 36228 22525
rect 39212 22516 39264 22568
rect 40592 22584 40644 22636
rect 43076 22627 43128 22636
rect 43076 22593 43085 22627
rect 43085 22593 43119 22627
rect 43119 22593 43128 22627
rect 43076 22584 43128 22593
rect 43812 22584 43864 22636
rect 46296 22584 46348 22636
rect 46848 22584 46900 22636
rect 42892 22559 42944 22568
rect 42892 22525 42901 22559
rect 42901 22525 42935 22559
rect 42935 22525 42944 22559
rect 42892 22516 42944 22525
rect 13176 22380 13228 22432
rect 15568 22423 15620 22432
rect 15568 22389 15577 22423
rect 15577 22389 15611 22423
rect 15611 22389 15620 22423
rect 15568 22380 15620 22389
rect 18052 22380 18104 22432
rect 21732 22380 21784 22432
rect 24216 22448 24268 22500
rect 32864 22448 32916 22500
rect 40224 22448 40276 22500
rect 23664 22380 23716 22432
rect 24400 22380 24452 22432
rect 30564 22423 30616 22432
rect 30564 22389 30573 22423
rect 30573 22389 30607 22423
rect 30607 22389 30616 22423
rect 30564 22380 30616 22389
rect 31392 22380 31444 22432
rect 32680 22423 32732 22432
rect 32680 22389 32689 22423
rect 32689 22389 32723 22423
rect 32723 22389 32732 22423
rect 32680 22380 32732 22389
rect 36544 22423 36596 22432
rect 36544 22389 36553 22423
rect 36553 22389 36587 22423
rect 36587 22389 36596 22423
rect 36544 22380 36596 22389
rect 40040 22380 40092 22432
rect 41512 22423 41564 22432
rect 41512 22389 41521 22423
rect 41521 22389 41555 22423
rect 41555 22389 41564 22423
rect 41512 22380 41564 22389
rect 43628 22380 43680 22432
rect 44364 22380 44416 22432
rect 45468 22380 45520 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 12532 22176 12584 22228
rect 14280 22219 14332 22228
rect 14280 22185 14289 22219
rect 14289 22185 14323 22219
rect 14323 22185 14332 22219
rect 14280 22176 14332 22185
rect 18512 22176 18564 22228
rect 29828 22176 29880 22228
rect 33968 22176 34020 22228
rect 39304 22176 39356 22228
rect 39396 22176 39448 22228
rect 40132 22176 40184 22228
rect 40500 22176 40552 22228
rect 4620 22108 4672 22160
rect 5264 22108 5316 22160
rect 11520 22108 11572 22160
rect 14924 22108 14976 22160
rect 23112 22108 23164 22160
rect 23572 22108 23624 22160
rect 33140 22151 33192 22160
rect 33140 22117 33149 22151
rect 33149 22117 33183 22151
rect 33183 22117 33192 22151
rect 33140 22108 33192 22117
rect 37188 22108 37240 22160
rect 42892 22108 42944 22160
rect 44088 22108 44140 22160
rect 13268 22083 13320 22092
rect 13268 22049 13277 22083
rect 13277 22049 13311 22083
rect 13311 22049 13320 22083
rect 13268 22040 13320 22049
rect 15568 22040 15620 22092
rect 15844 22083 15896 22092
rect 15844 22049 15853 22083
rect 15853 22049 15887 22083
rect 15887 22049 15896 22083
rect 15844 22040 15896 22049
rect 21732 22083 21784 22092
rect 2044 21972 2096 22024
rect 12808 21972 12860 22024
rect 13176 22015 13228 22024
rect 13176 21981 13185 22015
rect 13185 21981 13219 22015
rect 13219 21981 13228 22015
rect 13176 21972 13228 21981
rect 13912 21972 13964 22024
rect 17316 21972 17368 22024
rect 18144 21972 18196 22024
rect 21732 22049 21741 22083
rect 21741 22049 21775 22083
rect 21775 22049 21784 22083
rect 21732 22040 21784 22049
rect 22928 22040 22980 22092
rect 23112 22015 23164 22024
rect 23112 21981 23121 22015
rect 23121 21981 23155 22015
rect 23155 21981 23164 22015
rect 23112 21972 23164 21981
rect 23204 21972 23256 22024
rect 24492 21972 24544 22024
rect 25044 22015 25096 22024
rect 17776 21904 17828 21956
rect 20260 21947 20312 21956
rect 20260 21913 20269 21947
rect 20269 21913 20303 21947
rect 20303 21913 20312 21947
rect 25044 21981 25053 22015
rect 25053 21981 25087 22015
rect 25087 21981 25096 22015
rect 25044 21972 25096 21981
rect 26700 21972 26752 22024
rect 30472 22040 30524 22092
rect 20260 21904 20312 21913
rect 25596 21904 25648 21956
rect 25872 21947 25924 21956
rect 15936 21836 15988 21888
rect 18788 21879 18840 21888
rect 18788 21845 18797 21879
rect 18797 21845 18831 21879
rect 18831 21845 18840 21879
rect 18788 21836 18840 21845
rect 21456 21836 21508 21888
rect 21640 21879 21692 21888
rect 21640 21845 21649 21879
rect 21649 21845 21683 21879
rect 21683 21845 21692 21879
rect 22376 21879 22428 21888
rect 21640 21836 21692 21845
rect 22376 21845 22385 21879
rect 22385 21845 22419 21879
rect 22419 21845 22428 21879
rect 22376 21836 22428 21845
rect 23480 21879 23532 21888
rect 23480 21845 23489 21879
rect 23489 21845 23523 21879
rect 23523 21845 23532 21879
rect 23480 21836 23532 21845
rect 24584 21879 24636 21888
rect 24584 21845 24593 21879
rect 24593 21845 24627 21879
rect 24627 21845 24636 21879
rect 24584 21836 24636 21845
rect 25872 21913 25881 21947
rect 25881 21913 25915 21947
rect 25915 21913 25924 21947
rect 25872 21904 25924 21913
rect 26240 21904 26292 21956
rect 27620 21972 27672 22024
rect 30656 21972 30708 22024
rect 31208 21972 31260 22024
rect 34244 22040 34296 22092
rect 35900 22040 35952 22092
rect 40132 22040 40184 22092
rect 40960 22040 41012 22092
rect 41512 22040 41564 22092
rect 27160 21904 27212 21956
rect 30288 21904 30340 21956
rect 31576 21904 31628 21956
rect 33416 21972 33468 22024
rect 33876 22015 33928 22024
rect 33876 21981 33885 22015
rect 33885 21981 33919 22015
rect 33919 21981 33928 22015
rect 33876 21972 33928 21981
rect 34060 21972 34112 22024
rect 35072 21972 35124 22024
rect 37280 21972 37332 22024
rect 38476 22015 38528 22024
rect 38476 21981 38485 22015
rect 38485 21981 38519 22015
rect 38519 21981 38528 22015
rect 38476 21972 38528 21981
rect 39212 22015 39264 22024
rect 39212 21981 39221 22015
rect 39221 21981 39255 22015
rect 39255 21981 39264 22015
rect 39212 21972 39264 21981
rect 36544 21904 36596 21956
rect 39764 21972 39816 22024
rect 41052 21972 41104 22024
rect 46572 22108 46624 22160
rect 45928 22040 45980 22092
rect 46388 22083 46440 22092
rect 46388 22049 46397 22083
rect 46397 22049 46431 22083
rect 46431 22049 46440 22083
rect 46388 22040 46440 22049
rect 46664 22083 46716 22092
rect 46664 22049 46673 22083
rect 46673 22049 46707 22083
rect 46707 22049 46716 22083
rect 46664 22040 46716 22049
rect 40040 21947 40092 21956
rect 40040 21913 40049 21947
rect 40049 21913 40083 21947
rect 40083 21913 40092 21947
rect 40040 21904 40092 21913
rect 40224 21947 40276 21956
rect 40224 21913 40249 21947
rect 40249 21913 40276 21947
rect 40224 21904 40276 21913
rect 40868 21904 40920 21956
rect 45468 21972 45520 22024
rect 26148 21836 26200 21888
rect 27344 21836 27396 21888
rect 31116 21836 31168 21888
rect 31852 21836 31904 21888
rect 36084 21836 36136 21888
rect 36728 21836 36780 21888
rect 39488 21836 39540 21888
rect 43996 21879 44048 21888
rect 43996 21845 44005 21879
rect 44005 21845 44039 21879
rect 44039 21845 44048 21879
rect 43996 21836 44048 21845
rect 44088 21879 44140 21888
rect 44088 21845 44097 21879
rect 44097 21845 44131 21879
rect 44131 21845 44140 21879
rect 45192 21879 45244 21888
rect 44088 21836 44140 21845
rect 45192 21845 45201 21879
rect 45201 21845 45235 21879
rect 45235 21845 45244 21879
rect 45192 21836 45244 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 13268 21675 13320 21684
rect 13268 21641 13277 21675
rect 13277 21641 13311 21675
rect 13311 21641 13320 21675
rect 13268 21632 13320 21641
rect 13912 21675 13964 21684
rect 13912 21641 13921 21675
rect 13921 21641 13955 21675
rect 13955 21641 13964 21675
rect 13912 21632 13964 21641
rect 17776 21675 17828 21684
rect 17776 21641 17785 21675
rect 17785 21641 17819 21675
rect 17819 21641 17828 21675
rect 17776 21632 17828 21641
rect 21456 21675 21508 21684
rect 13176 21564 13228 21616
rect 21456 21641 21465 21675
rect 21465 21641 21499 21675
rect 21499 21641 21508 21675
rect 21456 21632 21508 21641
rect 21640 21632 21692 21684
rect 2044 21539 2096 21548
rect 2044 21505 2053 21539
rect 2053 21505 2087 21539
rect 2087 21505 2096 21539
rect 2044 21496 2096 21505
rect 9588 21539 9640 21548
rect 9588 21505 9597 21539
rect 9597 21505 9631 21539
rect 9631 21505 9640 21539
rect 9588 21496 9640 21505
rect 10416 21539 10468 21548
rect 10416 21505 10425 21539
rect 10425 21505 10459 21539
rect 10459 21505 10468 21539
rect 10416 21496 10468 21505
rect 12440 21496 12492 21548
rect 2320 21428 2372 21480
rect 2780 21471 2832 21480
rect 2780 21437 2789 21471
rect 2789 21437 2823 21471
rect 2823 21437 2832 21471
rect 2780 21428 2832 21437
rect 10324 21428 10376 21480
rect 10048 21360 10100 21412
rect 10232 21292 10284 21344
rect 13360 21428 13412 21480
rect 15844 21428 15896 21480
rect 16028 21471 16080 21480
rect 16028 21437 16037 21471
rect 16037 21437 16071 21471
rect 16071 21437 16080 21471
rect 16028 21428 16080 21437
rect 18052 21496 18104 21548
rect 20628 21564 20680 21616
rect 24584 21564 24636 21616
rect 25872 21632 25924 21684
rect 31208 21632 31260 21684
rect 31576 21675 31628 21684
rect 31576 21641 31585 21675
rect 31585 21641 31619 21675
rect 31619 21641 31628 21675
rect 31576 21632 31628 21641
rect 35624 21632 35676 21684
rect 40868 21675 40920 21684
rect 22376 21496 22428 21548
rect 23664 21496 23716 21548
rect 23848 21539 23900 21548
rect 23848 21505 23857 21539
rect 23857 21505 23891 21539
rect 23891 21505 23900 21539
rect 23848 21496 23900 21505
rect 25872 21539 25924 21548
rect 25872 21505 25881 21539
rect 25881 21505 25915 21539
rect 25915 21505 25924 21539
rect 25872 21496 25924 21505
rect 26240 21539 26292 21548
rect 26240 21505 26249 21539
rect 26249 21505 26283 21539
rect 26283 21505 26292 21539
rect 26240 21496 26292 21505
rect 30656 21564 30708 21616
rect 27252 21496 27304 21548
rect 28172 21496 28224 21548
rect 28724 21496 28776 21548
rect 29000 21539 29052 21548
rect 29000 21505 29016 21539
rect 29016 21505 29050 21539
rect 29050 21505 29052 21539
rect 29276 21539 29328 21548
rect 29000 21496 29052 21505
rect 29276 21505 29299 21539
rect 29299 21505 29328 21539
rect 29276 21496 29328 21505
rect 31024 21539 31076 21548
rect 18788 21428 18840 21480
rect 25228 21428 25280 21480
rect 12164 21292 12216 21344
rect 13820 21292 13872 21344
rect 23112 21292 23164 21344
rect 29000 21360 29052 21412
rect 31024 21505 31033 21539
rect 31033 21505 31067 21539
rect 31067 21505 31076 21539
rect 31024 21496 31076 21505
rect 31116 21539 31168 21548
rect 31116 21505 31125 21539
rect 31125 21505 31159 21539
rect 31159 21505 31168 21539
rect 31392 21539 31444 21548
rect 31116 21496 31168 21505
rect 31392 21505 31401 21539
rect 31401 21505 31435 21539
rect 31435 21505 31444 21539
rect 31392 21496 31444 21505
rect 32956 21539 33008 21548
rect 32956 21505 32965 21539
rect 32965 21505 32999 21539
rect 32999 21505 33008 21539
rect 32956 21496 33008 21505
rect 33140 21539 33192 21548
rect 33140 21505 33149 21539
rect 33149 21505 33183 21539
rect 33183 21505 33192 21539
rect 33140 21496 33192 21505
rect 33232 21539 33284 21548
rect 33232 21505 33241 21539
rect 33241 21505 33275 21539
rect 33275 21505 33284 21539
rect 33784 21564 33836 21616
rect 33968 21607 34020 21616
rect 33968 21573 34002 21607
rect 34002 21573 34020 21607
rect 33968 21564 34020 21573
rect 39856 21607 39908 21616
rect 39856 21573 39865 21607
rect 39865 21573 39899 21607
rect 39899 21573 39908 21607
rect 39856 21564 39908 21573
rect 40868 21641 40877 21675
rect 40877 21641 40911 21675
rect 40911 21641 40920 21675
rect 40868 21632 40920 21641
rect 43076 21632 43128 21684
rect 43812 21632 43864 21684
rect 45928 21632 45980 21684
rect 33232 21496 33284 21505
rect 31208 21471 31260 21480
rect 31208 21437 31217 21471
rect 31217 21437 31251 21471
rect 31251 21437 31260 21471
rect 36176 21496 36228 21548
rect 37188 21496 37240 21548
rect 39488 21496 39540 21548
rect 39764 21539 39816 21546
rect 39764 21505 39771 21539
rect 39771 21505 39816 21539
rect 39764 21494 39816 21505
rect 31208 21428 31260 21437
rect 35072 21403 35124 21412
rect 35072 21369 35081 21403
rect 35081 21369 35115 21403
rect 35115 21369 35124 21403
rect 40592 21496 40644 21548
rect 40776 21539 40828 21548
rect 40776 21505 40785 21539
rect 40785 21505 40819 21539
rect 40819 21505 40828 21539
rect 40776 21496 40828 21505
rect 43076 21496 43128 21548
rect 35072 21360 35124 21369
rect 40592 21360 40644 21412
rect 42800 21428 42852 21480
rect 40960 21360 41012 21412
rect 43352 21496 43404 21548
rect 43628 21496 43680 21548
rect 44364 21539 44416 21548
rect 44364 21505 44373 21539
rect 44373 21505 44407 21539
rect 44407 21505 44416 21539
rect 44364 21496 44416 21505
rect 45192 21564 45244 21616
rect 47032 21539 47084 21548
rect 47032 21505 47041 21539
rect 47041 21505 47075 21539
rect 47075 21505 47084 21539
rect 47032 21496 47084 21505
rect 43444 21360 43496 21412
rect 28540 21335 28592 21344
rect 28540 21301 28549 21335
rect 28549 21301 28583 21335
rect 28583 21301 28592 21335
rect 28540 21292 28592 21301
rect 28908 21292 28960 21344
rect 32956 21292 33008 21344
rect 36268 21292 36320 21344
rect 38108 21292 38160 21344
rect 38568 21292 38620 21344
rect 38936 21292 38988 21344
rect 40316 21292 40368 21344
rect 46664 21292 46716 21344
rect 47952 21335 48004 21344
rect 47952 21301 47961 21335
rect 47961 21301 47995 21335
rect 47995 21301 48004 21335
rect 47952 21292 48004 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 2320 21131 2372 21140
rect 2320 21097 2329 21131
rect 2329 21097 2363 21131
rect 2363 21097 2372 21131
rect 2320 21088 2372 21097
rect 12808 21131 12860 21140
rect 12808 21097 12817 21131
rect 12817 21097 12851 21131
rect 12851 21097 12860 21131
rect 12808 21088 12860 21097
rect 16028 21088 16080 21140
rect 25044 21088 25096 21140
rect 27160 21131 27212 21140
rect 27160 21097 27169 21131
rect 27169 21097 27203 21131
rect 27203 21097 27212 21131
rect 27160 21088 27212 21097
rect 29276 21088 29328 21140
rect 33232 21088 33284 21140
rect 2320 20884 2372 20936
rect 4160 20884 4212 20936
rect 3516 20816 3568 20868
rect 10232 20995 10284 21004
rect 10232 20961 10241 20995
rect 10241 20961 10275 20995
rect 10275 20961 10284 20995
rect 10232 20952 10284 20961
rect 23480 21020 23532 21072
rect 13268 20995 13320 21004
rect 13268 20961 13277 20995
rect 13277 20961 13311 20995
rect 13311 20961 13320 20995
rect 13268 20952 13320 20961
rect 13360 20995 13412 21004
rect 13360 20961 13369 20995
rect 13369 20961 13403 20995
rect 13403 20961 13412 20995
rect 23848 20995 23900 21004
rect 13360 20952 13412 20961
rect 23848 20961 23857 20995
rect 23857 20961 23891 20995
rect 23891 20961 23900 20995
rect 23848 20952 23900 20961
rect 10048 20927 10100 20936
rect 10048 20893 10057 20927
rect 10057 20893 10091 20927
rect 10091 20893 10100 20927
rect 10048 20884 10100 20893
rect 12164 20884 12216 20936
rect 19984 20927 20036 20936
rect 19984 20893 19993 20927
rect 19993 20893 20027 20927
rect 20027 20893 20036 20927
rect 19984 20884 20036 20893
rect 23388 20884 23440 20936
rect 24400 20884 24452 20936
rect 28356 21020 28408 21072
rect 31024 21020 31076 21072
rect 34244 21020 34296 21072
rect 25872 20884 25924 20936
rect 15200 20816 15252 20868
rect 22100 20816 22152 20868
rect 30380 20952 30432 21004
rect 31392 20952 31444 21004
rect 41052 21088 41104 21140
rect 42892 21088 42944 21140
rect 43444 21131 43496 21140
rect 43444 21097 43453 21131
rect 43453 21097 43487 21131
rect 43487 21097 43496 21131
rect 43444 21088 43496 21097
rect 43996 21088 44048 21140
rect 48044 21088 48096 21140
rect 26148 20927 26200 20936
rect 26148 20893 26157 20927
rect 26157 20893 26191 20927
rect 26191 20893 26200 20927
rect 28172 20927 28224 20936
rect 26148 20884 26200 20893
rect 28172 20893 28181 20927
rect 28181 20893 28215 20927
rect 28215 20893 28224 20927
rect 28172 20884 28224 20893
rect 28356 20927 28408 20936
rect 28356 20893 28365 20927
rect 28365 20893 28399 20927
rect 28399 20893 28408 20927
rect 28356 20884 28408 20893
rect 13176 20791 13228 20800
rect 13176 20757 13185 20791
rect 13185 20757 13219 20791
rect 13219 20757 13228 20791
rect 13176 20748 13228 20757
rect 19432 20748 19484 20800
rect 23204 20748 23256 20800
rect 28632 20884 28684 20936
rect 28724 20927 28776 20936
rect 28724 20893 28733 20927
rect 28733 20893 28767 20927
rect 28767 20893 28776 20927
rect 28724 20884 28776 20893
rect 32680 20927 32732 20936
rect 32680 20893 32689 20927
rect 32689 20893 32723 20927
rect 32723 20893 32732 20927
rect 32680 20884 32732 20893
rect 32864 20927 32916 20936
rect 32864 20893 32873 20927
rect 32873 20893 32907 20927
rect 32907 20893 32916 20927
rect 32864 20884 32916 20893
rect 33692 20927 33744 20936
rect 33692 20893 33701 20927
rect 33701 20893 33735 20927
rect 33735 20893 33744 20927
rect 33692 20884 33744 20893
rect 34152 20884 34204 20936
rect 38108 20927 38160 20936
rect 31944 20816 31996 20868
rect 33876 20859 33928 20868
rect 33876 20825 33885 20859
rect 33885 20825 33919 20859
rect 33919 20825 33928 20859
rect 33876 20816 33928 20825
rect 38108 20893 38117 20927
rect 38117 20893 38151 20927
rect 38151 20893 38160 20927
rect 38108 20884 38160 20893
rect 42708 20952 42760 21004
rect 40040 20927 40092 20936
rect 40040 20893 40049 20927
rect 40049 20893 40083 20927
rect 40083 20893 40092 20927
rect 40040 20884 40092 20893
rect 40316 20927 40368 20936
rect 40316 20893 40350 20927
rect 40350 20893 40368 20927
rect 40316 20884 40368 20893
rect 42800 20927 42852 20936
rect 38752 20816 38804 20868
rect 26700 20748 26752 20800
rect 28448 20748 28500 20800
rect 28632 20748 28684 20800
rect 31208 20748 31260 20800
rect 37924 20748 37976 20800
rect 38292 20748 38344 20800
rect 42800 20893 42809 20927
rect 42809 20893 42843 20927
rect 42843 20893 42852 20927
rect 42800 20884 42852 20893
rect 42984 20884 43036 20936
rect 43076 20816 43128 20868
rect 45468 20952 45520 21004
rect 47952 21020 48004 21072
rect 46664 20995 46716 21004
rect 46664 20961 46673 20995
rect 46673 20961 46707 20995
rect 46707 20961 46716 20995
rect 46664 20952 46716 20961
rect 48228 20995 48280 21004
rect 48228 20961 48237 20995
rect 48237 20961 48271 20995
rect 48271 20961 48280 20995
rect 48228 20952 48280 20961
rect 45928 20884 45980 20936
rect 43352 20748 43404 20800
rect 44272 20748 44324 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 5080 20544 5132 20596
rect 9588 20544 9640 20596
rect 12440 20587 12492 20596
rect 12440 20553 12449 20587
rect 12449 20553 12483 20587
rect 12483 20553 12492 20587
rect 12440 20544 12492 20553
rect 17868 20544 17920 20596
rect 17960 20544 18012 20596
rect 22100 20544 22152 20596
rect 23388 20544 23440 20596
rect 13176 20476 13228 20528
rect 4160 20451 4212 20460
rect 4160 20417 4169 20451
rect 4169 20417 4203 20451
rect 4203 20417 4212 20451
rect 4160 20408 4212 20417
rect 12532 20408 12584 20460
rect 13820 20408 13872 20460
rect 19064 20408 19116 20460
rect 19432 20476 19484 20528
rect 24400 20519 24452 20528
rect 24400 20485 24409 20519
rect 24409 20485 24443 20519
rect 24443 20485 24452 20519
rect 24400 20476 24452 20485
rect 27252 20544 27304 20596
rect 29184 20587 29236 20596
rect 29184 20553 29193 20587
rect 29193 20553 29227 20587
rect 29227 20553 29236 20587
rect 29184 20544 29236 20553
rect 23388 20451 23440 20460
rect 4896 20340 4948 20392
rect 10140 20383 10192 20392
rect 2964 20272 3016 20324
rect 10140 20349 10149 20383
rect 10149 20349 10183 20383
rect 10183 20349 10192 20383
rect 10140 20340 10192 20349
rect 10324 20340 10376 20392
rect 15292 20340 15344 20392
rect 15844 20340 15896 20392
rect 18144 20340 18196 20392
rect 23388 20417 23397 20451
rect 23397 20417 23431 20451
rect 23431 20417 23440 20451
rect 23388 20408 23440 20417
rect 23480 20408 23532 20460
rect 27344 20451 27396 20460
rect 27344 20417 27353 20451
rect 27353 20417 27387 20451
rect 27387 20417 27396 20451
rect 27344 20408 27396 20417
rect 28540 20476 28592 20528
rect 28448 20408 28500 20460
rect 28908 20408 28960 20460
rect 33140 20544 33192 20596
rect 35624 20544 35676 20596
rect 41880 20544 41932 20596
rect 31024 20451 31076 20460
rect 23756 20383 23808 20392
rect 23756 20349 23765 20383
rect 23765 20349 23799 20383
rect 23799 20349 23808 20383
rect 23756 20340 23808 20349
rect 31024 20417 31033 20451
rect 31033 20417 31067 20451
rect 31067 20417 31076 20451
rect 31024 20408 31076 20417
rect 31208 20451 31260 20460
rect 31208 20417 31217 20451
rect 31217 20417 31251 20451
rect 31251 20417 31260 20451
rect 31208 20408 31260 20417
rect 31668 20408 31720 20460
rect 33692 20451 33744 20460
rect 33692 20417 33701 20451
rect 33701 20417 33735 20451
rect 33735 20417 33744 20451
rect 33692 20408 33744 20417
rect 33876 20451 33928 20460
rect 33876 20417 33885 20451
rect 33885 20417 33919 20451
rect 33919 20417 33928 20451
rect 33876 20408 33928 20417
rect 34520 20451 34572 20460
rect 31300 20383 31352 20392
rect 31300 20349 31309 20383
rect 31309 20349 31343 20383
rect 31343 20349 31352 20383
rect 31300 20340 31352 20349
rect 34520 20417 34529 20451
rect 34529 20417 34563 20451
rect 34563 20417 34572 20451
rect 34520 20408 34572 20417
rect 40040 20476 40092 20528
rect 40408 20476 40460 20528
rect 40500 20476 40552 20528
rect 42708 20476 42760 20528
rect 37740 20451 37792 20460
rect 37740 20417 37774 20451
rect 37774 20417 37792 20451
rect 40316 20451 40368 20460
rect 37740 20408 37792 20417
rect 40316 20417 40325 20451
rect 40325 20417 40359 20451
rect 40359 20417 40368 20451
rect 40316 20408 40368 20417
rect 40592 20408 40644 20460
rect 46572 20408 46624 20460
rect 46848 20408 46900 20460
rect 34796 20340 34848 20392
rect 39856 20340 39908 20392
rect 40868 20383 40920 20392
rect 40868 20349 40877 20383
rect 40877 20349 40911 20383
rect 40911 20349 40920 20383
rect 40868 20340 40920 20349
rect 15384 20204 15436 20256
rect 18236 20247 18288 20256
rect 18236 20213 18245 20247
rect 18245 20213 18279 20247
rect 18279 20213 18288 20247
rect 18236 20204 18288 20213
rect 20628 20272 20680 20324
rect 35624 20272 35676 20324
rect 23572 20204 23624 20256
rect 24860 20204 24912 20256
rect 26240 20204 26292 20256
rect 29000 20204 29052 20256
rect 29368 20204 29420 20256
rect 30932 20204 30984 20256
rect 33876 20204 33928 20256
rect 38200 20204 38252 20256
rect 46664 20204 46716 20256
rect 47952 20247 48004 20256
rect 47952 20213 47961 20247
rect 47961 20213 47995 20247
rect 47995 20213 48004 20247
rect 47952 20204 48004 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 4896 20043 4948 20052
rect 4896 20009 4905 20043
rect 4905 20009 4939 20043
rect 4939 20009 4948 20043
rect 4896 20000 4948 20009
rect 15200 20043 15252 20052
rect 15200 20009 15209 20043
rect 15209 20009 15243 20043
rect 15243 20009 15252 20043
rect 15200 20000 15252 20009
rect 17868 20000 17920 20052
rect 20536 20000 20588 20052
rect 23572 20000 23624 20052
rect 28172 20000 28224 20052
rect 29000 20000 29052 20052
rect 30104 20000 30156 20052
rect 32680 20000 32732 20052
rect 33692 20000 33744 20052
rect 34152 20043 34204 20052
rect 34152 20009 34161 20043
rect 34161 20009 34195 20043
rect 34195 20009 34204 20043
rect 34152 20000 34204 20009
rect 34244 20000 34296 20052
rect 35440 20000 35492 20052
rect 37740 20043 37792 20052
rect 23388 19932 23440 19984
rect 33968 19932 34020 19984
rect 37740 20009 37749 20043
rect 37749 20009 37783 20043
rect 37783 20009 37792 20043
rect 37740 20000 37792 20009
rect 40224 20000 40276 20052
rect 40684 20000 40736 20052
rect 39948 19932 40000 19984
rect 4804 19839 4856 19848
rect 4804 19805 4813 19839
rect 4813 19805 4847 19839
rect 4847 19805 4856 19839
rect 4804 19796 4856 19805
rect 5540 19796 5592 19848
rect 204 19728 256 19780
rect 18144 19864 18196 19916
rect 19340 19864 19392 19916
rect 30656 19907 30708 19916
rect 9588 19839 9640 19848
rect 9588 19805 9597 19839
rect 9597 19805 9631 19839
rect 9631 19805 9640 19839
rect 9588 19796 9640 19805
rect 10232 19839 10284 19848
rect 10232 19805 10241 19839
rect 10241 19805 10275 19839
rect 10275 19805 10284 19839
rect 10232 19796 10284 19805
rect 15384 19839 15436 19848
rect 15384 19805 15393 19839
rect 15393 19805 15427 19839
rect 15427 19805 15436 19839
rect 15384 19796 15436 19805
rect 15936 19796 15988 19848
rect 17960 19839 18012 19848
rect 17960 19805 17969 19839
rect 17969 19805 18003 19839
rect 18003 19805 18012 19839
rect 17960 19796 18012 19805
rect 20628 19839 20680 19848
rect 20628 19805 20637 19839
rect 20637 19805 20671 19839
rect 20671 19805 20680 19839
rect 20628 19796 20680 19805
rect 22376 19839 22428 19848
rect 22376 19805 22385 19839
rect 22385 19805 22419 19839
rect 22419 19805 22428 19839
rect 22376 19796 22428 19805
rect 22652 19839 22704 19848
rect 22652 19805 22661 19839
rect 22661 19805 22695 19839
rect 22695 19805 22704 19839
rect 22652 19796 22704 19805
rect 23480 19796 23532 19848
rect 30656 19873 30665 19907
rect 30665 19873 30699 19907
rect 30699 19873 30708 19907
rect 30656 19864 30708 19873
rect 27988 19796 28040 19848
rect 28448 19839 28500 19848
rect 28448 19805 28457 19839
rect 28457 19805 28491 19839
rect 28491 19805 28500 19839
rect 28448 19796 28500 19805
rect 28724 19839 28776 19848
rect 28724 19805 28733 19839
rect 28733 19805 28767 19839
rect 28767 19805 28776 19839
rect 28724 19796 28776 19805
rect 30932 19839 30984 19848
rect 30932 19805 30966 19839
rect 30966 19805 30984 19839
rect 30932 19796 30984 19805
rect 25136 19728 25188 19780
rect 32956 19864 33008 19916
rect 35440 19864 35492 19916
rect 38200 19907 38252 19916
rect 38200 19873 38209 19907
rect 38209 19873 38243 19907
rect 38243 19873 38252 19907
rect 38200 19864 38252 19873
rect 32496 19839 32548 19848
rect 32496 19805 32505 19839
rect 32505 19805 32539 19839
rect 32539 19805 32548 19839
rect 32496 19796 32548 19805
rect 32864 19796 32916 19848
rect 34520 19796 34572 19848
rect 15476 19660 15528 19712
rect 20076 19660 20128 19712
rect 22192 19703 22244 19712
rect 22192 19669 22201 19703
rect 22201 19669 22235 19703
rect 22235 19669 22244 19703
rect 22192 19660 22244 19669
rect 29460 19660 29512 19712
rect 32036 19703 32088 19712
rect 32036 19669 32045 19703
rect 32045 19669 32079 19703
rect 32079 19669 32088 19703
rect 32864 19703 32916 19712
rect 32036 19660 32088 19669
rect 32864 19669 32873 19703
rect 32873 19669 32907 19703
rect 32907 19669 32916 19703
rect 32864 19660 32916 19669
rect 37280 19796 37332 19848
rect 37924 19839 37976 19848
rect 37924 19805 37933 19839
rect 37933 19805 37967 19839
rect 37967 19805 37976 19839
rect 37924 19796 37976 19805
rect 40408 19864 40460 19916
rect 44456 19864 44508 19916
rect 47952 19932 48004 19984
rect 46664 19907 46716 19916
rect 46664 19873 46673 19907
rect 46673 19873 46707 19907
rect 46707 19873 46716 19907
rect 46664 19864 46716 19873
rect 48228 19907 48280 19916
rect 48228 19873 48237 19907
rect 48237 19873 48271 19907
rect 48271 19873 48280 19907
rect 48228 19864 48280 19873
rect 42156 19839 42208 19848
rect 35624 19728 35676 19780
rect 35992 19728 36044 19780
rect 42156 19805 42165 19839
rect 42165 19805 42199 19839
rect 42199 19805 42208 19839
rect 42156 19796 42208 19805
rect 44272 19796 44324 19848
rect 44548 19796 44600 19848
rect 34244 19660 34296 19712
rect 35348 19660 35400 19712
rect 35716 19660 35768 19712
rect 38384 19728 38436 19780
rect 39028 19728 39080 19780
rect 43444 19728 43496 19780
rect 37464 19660 37516 19712
rect 41880 19660 41932 19712
rect 43352 19660 43404 19712
rect 44180 19660 44232 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 12532 19456 12584 19508
rect 19064 19499 19116 19508
rect 19064 19465 19073 19499
rect 19073 19465 19107 19499
rect 19107 19465 19116 19499
rect 19064 19456 19116 19465
rect 19984 19456 20036 19508
rect 26424 19456 26476 19508
rect 28724 19456 28776 19508
rect 29460 19499 29512 19508
rect 29460 19465 29469 19499
rect 29469 19465 29503 19499
rect 29503 19465 29512 19499
rect 29460 19456 29512 19465
rect 31024 19499 31076 19508
rect 31024 19465 31033 19499
rect 31033 19465 31067 19499
rect 31067 19465 31076 19499
rect 31024 19456 31076 19465
rect 32680 19456 32732 19508
rect 35716 19456 35768 19508
rect 35992 19456 36044 19508
rect 9956 19363 10008 19372
rect 9956 19329 9965 19363
rect 9965 19329 9999 19363
rect 9999 19329 10008 19363
rect 9956 19320 10008 19329
rect 11520 19320 11572 19372
rect 11796 19320 11848 19372
rect 13912 19363 13964 19372
rect 13912 19329 13921 19363
rect 13921 19329 13955 19363
rect 13955 19329 13964 19363
rect 13912 19320 13964 19329
rect 14924 19363 14976 19372
rect 14924 19329 14933 19363
rect 14933 19329 14967 19363
rect 14967 19329 14976 19363
rect 14924 19320 14976 19329
rect 10048 19295 10100 19304
rect 10048 19261 10057 19295
rect 10057 19261 10091 19295
rect 10091 19261 10100 19295
rect 10048 19252 10100 19261
rect 10232 19252 10284 19304
rect 14096 19252 14148 19304
rect 15016 19252 15068 19304
rect 15200 19116 15252 19168
rect 18880 19431 18932 19440
rect 18880 19397 18889 19431
rect 18889 19397 18923 19431
rect 18923 19397 18932 19431
rect 18880 19388 18932 19397
rect 20260 19388 20312 19440
rect 24768 19388 24820 19440
rect 17868 19363 17920 19372
rect 17868 19329 17877 19363
rect 17877 19329 17911 19363
rect 17911 19329 17920 19363
rect 17868 19320 17920 19329
rect 22928 19363 22980 19372
rect 22928 19329 22937 19363
rect 22937 19329 22971 19363
rect 22971 19329 22980 19363
rect 22928 19320 22980 19329
rect 23112 19320 23164 19372
rect 19340 19252 19392 19304
rect 22652 19252 22704 19304
rect 24860 19320 24912 19372
rect 30288 19388 30340 19440
rect 32864 19388 32916 19440
rect 26792 19320 26844 19372
rect 27344 19363 27396 19372
rect 20076 19227 20128 19236
rect 20076 19193 20085 19227
rect 20085 19193 20119 19227
rect 20119 19193 20128 19227
rect 20076 19184 20128 19193
rect 22468 19116 22520 19168
rect 23756 19116 23808 19168
rect 24676 19159 24728 19168
rect 24676 19125 24685 19159
rect 24685 19125 24719 19159
rect 24719 19125 24728 19159
rect 24676 19116 24728 19125
rect 26332 19184 26384 19236
rect 27344 19329 27353 19363
rect 27353 19329 27387 19363
rect 27387 19329 27396 19363
rect 27344 19320 27396 19329
rect 28264 19320 28316 19372
rect 28724 19363 28776 19372
rect 28080 19295 28132 19304
rect 28080 19261 28089 19295
rect 28089 19261 28123 19295
rect 28123 19261 28132 19295
rect 28080 19252 28132 19261
rect 28724 19329 28733 19363
rect 28733 19329 28767 19363
rect 28767 19329 28776 19363
rect 28724 19320 28776 19329
rect 29368 19363 29420 19372
rect 28632 19252 28684 19304
rect 29368 19329 29377 19363
rect 29377 19329 29411 19363
rect 29411 19329 29420 19363
rect 29368 19320 29420 19329
rect 29920 19320 29972 19372
rect 31024 19320 31076 19372
rect 31484 19363 31536 19372
rect 31484 19329 31493 19363
rect 31493 19329 31527 19363
rect 31527 19329 31536 19363
rect 31484 19320 31536 19329
rect 32036 19320 32088 19372
rect 33692 19320 33744 19372
rect 33968 19320 34020 19372
rect 35348 19363 35400 19372
rect 35348 19329 35357 19363
rect 35357 19329 35391 19363
rect 35391 19329 35400 19363
rect 35348 19320 35400 19329
rect 27712 19184 27764 19236
rect 28724 19184 28776 19236
rect 31576 19252 31628 19304
rect 35256 19252 35308 19304
rect 35532 19388 35584 19440
rect 35808 19388 35860 19440
rect 40132 19499 40184 19508
rect 40132 19465 40141 19499
rect 40141 19465 40175 19499
rect 40175 19465 40184 19499
rect 40132 19456 40184 19465
rect 43536 19499 43588 19508
rect 43536 19465 43545 19499
rect 43545 19465 43579 19499
rect 43579 19465 43588 19499
rect 43536 19456 43588 19465
rect 37464 19431 37516 19440
rect 37464 19397 37473 19431
rect 37473 19397 37507 19431
rect 37507 19397 37516 19431
rect 37464 19388 37516 19397
rect 38200 19388 38252 19440
rect 43444 19388 43496 19440
rect 43812 19456 43864 19508
rect 39948 19363 40000 19372
rect 39948 19329 39957 19363
rect 39957 19329 39991 19363
rect 39991 19329 40000 19363
rect 39948 19320 40000 19329
rect 41880 19363 41932 19372
rect 41880 19329 41889 19363
rect 41889 19329 41923 19363
rect 41923 19329 41932 19363
rect 41880 19320 41932 19329
rect 42800 19320 42852 19372
rect 43352 19363 43404 19372
rect 43352 19329 43361 19363
rect 43361 19329 43395 19363
rect 43395 19329 43404 19363
rect 43352 19320 43404 19329
rect 44272 19388 44324 19440
rect 44456 19363 44508 19372
rect 44456 19329 44465 19363
rect 44465 19329 44499 19363
rect 44499 19329 44508 19363
rect 44456 19320 44508 19329
rect 47308 19320 47360 19372
rect 35900 19252 35952 19304
rect 39488 19252 39540 19304
rect 40316 19252 40368 19304
rect 33600 19184 33652 19236
rect 27068 19116 27120 19168
rect 27528 19116 27580 19168
rect 29000 19116 29052 19168
rect 34152 19159 34204 19168
rect 34152 19125 34161 19159
rect 34161 19125 34195 19159
rect 34195 19125 34204 19159
rect 34152 19116 34204 19125
rect 34428 19159 34480 19168
rect 34428 19125 34437 19159
rect 34437 19125 34471 19159
rect 34471 19125 34480 19159
rect 34428 19116 34480 19125
rect 36636 19116 36688 19168
rect 43076 19116 43128 19168
rect 44272 19159 44324 19168
rect 44272 19125 44281 19159
rect 44281 19125 44315 19159
rect 44315 19125 44324 19159
rect 44272 19116 44324 19125
rect 47124 19159 47176 19168
rect 47124 19125 47133 19159
rect 47133 19125 47167 19159
rect 47167 19125 47176 19159
rect 47124 19116 47176 19125
rect 47952 19159 48004 19168
rect 47952 19125 47961 19159
rect 47961 19125 47995 19159
rect 47995 19125 48004 19159
rect 47952 19116 48004 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 11796 18912 11848 18964
rect 22928 18912 22980 18964
rect 26792 18955 26844 18964
rect 13912 18844 13964 18896
rect 24676 18844 24728 18896
rect 25964 18844 26016 18896
rect 12716 18819 12768 18828
rect 12716 18785 12725 18819
rect 12725 18785 12759 18819
rect 12759 18785 12768 18819
rect 12716 18776 12768 18785
rect 2044 18708 2096 18760
rect 12256 18708 12308 18760
rect 12532 18708 12584 18760
rect 13912 18708 13964 18760
rect 15476 18708 15528 18760
rect 16764 18708 16816 18760
rect 18144 18708 18196 18760
rect 24768 18751 24820 18760
rect 24768 18717 24777 18751
rect 24777 18717 24811 18751
rect 24811 18717 24820 18751
rect 24768 18708 24820 18717
rect 26424 18844 26476 18896
rect 26332 18819 26384 18828
rect 26332 18785 26341 18819
rect 26341 18785 26375 18819
rect 26375 18785 26384 18819
rect 26332 18776 26384 18785
rect 26240 18751 26292 18760
rect 9956 18640 10008 18692
rect 16396 18640 16448 18692
rect 18236 18640 18288 18692
rect 22192 18640 22244 18692
rect 22744 18640 22796 18692
rect 16028 18572 16080 18624
rect 17868 18572 17920 18624
rect 24584 18615 24636 18624
rect 24584 18581 24593 18615
rect 24593 18581 24627 18615
rect 24627 18581 24636 18615
rect 24584 18572 24636 18581
rect 26240 18717 26249 18751
rect 26249 18717 26283 18751
rect 26283 18717 26292 18751
rect 26240 18708 26292 18717
rect 26792 18921 26801 18955
rect 26801 18921 26835 18955
rect 26835 18921 26844 18955
rect 26792 18912 26844 18921
rect 27528 18912 27580 18964
rect 29000 18912 29052 18964
rect 31484 18912 31536 18964
rect 31576 18912 31628 18964
rect 34152 18912 34204 18964
rect 35440 18912 35492 18964
rect 35532 18912 35584 18964
rect 36268 18912 36320 18964
rect 38292 18912 38344 18964
rect 39028 18955 39080 18964
rect 39028 18921 39037 18955
rect 39037 18921 39071 18955
rect 39071 18921 39080 18955
rect 39028 18912 39080 18921
rect 42156 18912 42208 18964
rect 27068 18844 27120 18896
rect 31300 18844 31352 18896
rect 34520 18844 34572 18896
rect 35900 18844 35952 18896
rect 37188 18844 37240 18896
rect 40868 18844 40920 18896
rect 28540 18776 28592 18828
rect 27528 18751 27580 18760
rect 27528 18717 27537 18751
rect 27537 18717 27571 18751
rect 27571 18717 27580 18751
rect 27528 18708 27580 18717
rect 27252 18640 27304 18692
rect 30380 18708 30432 18760
rect 30840 18776 30892 18828
rect 31208 18776 31260 18828
rect 33140 18776 33192 18828
rect 33784 18776 33836 18828
rect 34428 18776 34480 18828
rect 34796 18776 34848 18828
rect 28540 18640 28592 18692
rect 30564 18751 30616 18760
rect 30564 18717 30573 18751
rect 30573 18717 30607 18751
rect 30607 18717 30616 18751
rect 33876 18751 33928 18760
rect 30564 18708 30616 18717
rect 31116 18683 31168 18692
rect 31116 18649 31125 18683
rect 31125 18649 31159 18683
rect 31159 18649 31168 18683
rect 31116 18640 31168 18649
rect 26608 18572 26660 18624
rect 27436 18572 27488 18624
rect 29184 18572 29236 18624
rect 30104 18615 30156 18624
rect 30104 18581 30113 18615
rect 30113 18581 30147 18615
rect 30147 18581 30156 18615
rect 30104 18572 30156 18581
rect 33876 18717 33885 18751
rect 33885 18717 33919 18751
rect 33919 18717 33928 18751
rect 33876 18708 33928 18717
rect 35624 18776 35676 18828
rect 33692 18683 33744 18692
rect 33692 18649 33701 18683
rect 33701 18649 33735 18683
rect 33735 18649 33744 18683
rect 33692 18640 33744 18649
rect 34888 18640 34940 18692
rect 35808 18708 35860 18760
rect 44456 18844 44508 18896
rect 38476 18708 38528 18760
rect 39120 18751 39172 18760
rect 39120 18717 39129 18751
rect 39129 18717 39163 18751
rect 39163 18717 39172 18751
rect 39120 18708 39172 18717
rect 40132 18708 40184 18760
rect 40776 18751 40828 18760
rect 40776 18717 40785 18751
rect 40785 18717 40819 18751
rect 40819 18717 40828 18751
rect 40776 18708 40828 18717
rect 42800 18751 42852 18760
rect 42800 18717 42809 18751
rect 42809 18717 42843 18751
rect 42843 18717 42852 18751
rect 42800 18708 42852 18717
rect 42892 18751 42944 18760
rect 42892 18717 42901 18751
rect 42901 18717 42935 18751
rect 42935 18717 42944 18751
rect 42892 18708 42944 18717
rect 43076 18751 43128 18760
rect 43076 18717 43085 18751
rect 43085 18717 43119 18751
rect 43119 18717 43128 18751
rect 44180 18776 44232 18828
rect 47952 18844 48004 18896
rect 43076 18708 43128 18717
rect 44272 18751 44324 18760
rect 44272 18717 44281 18751
rect 44281 18717 44315 18751
rect 44315 18717 44324 18751
rect 44272 18708 44324 18717
rect 47124 18776 47176 18828
rect 48228 18819 48280 18828
rect 48228 18785 48237 18819
rect 48237 18785 48271 18819
rect 48271 18785 48280 18819
rect 48228 18776 48280 18785
rect 36636 18640 36688 18692
rect 43352 18640 43404 18692
rect 43536 18640 43588 18692
rect 44180 18640 44232 18692
rect 33968 18615 34020 18624
rect 33968 18581 33977 18615
rect 33977 18581 34011 18615
rect 34011 18581 34020 18615
rect 33968 18572 34020 18581
rect 35900 18615 35952 18624
rect 35900 18581 35909 18615
rect 35909 18581 35943 18615
rect 35943 18581 35952 18615
rect 35900 18572 35952 18581
rect 38660 18615 38712 18624
rect 38660 18581 38669 18615
rect 38669 18581 38703 18615
rect 38703 18581 38712 18615
rect 38660 18572 38712 18581
rect 44640 18615 44692 18624
rect 44640 18581 44649 18615
rect 44649 18581 44683 18615
rect 44683 18581 44692 18615
rect 44640 18572 44692 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 12256 18411 12308 18420
rect 12256 18377 12265 18411
rect 12265 18377 12299 18411
rect 12299 18377 12308 18411
rect 12256 18368 12308 18377
rect 16396 18368 16448 18420
rect 2044 18275 2096 18284
rect 2044 18241 2053 18275
rect 2053 18241 2087 18275
rect 2087 18241 2096 18275
rect 2044 18232 2096 18241
rect 17868 18300 17920 18352
rect 22376 18368 22428 18420
rect 33600 18368 33652 18420
rect 36636 18411 36688 18420
rect 36636 18377 36645 18411
rect 36645 18377 36679 18411
rect 36679 18377 36688 18411
rect 36636 18368 36688 18377
rect 38476 18411 38528 18420
rect 38476 18377 38485 18411
rect 38485 18377 38519 18411
rect 38519 18377 38528 18411
rect 38476 18368 38528 18377
rect 24584 18300 24636 18352
rect 27252 18300 27304 18352
rect 27528 18300 27580 18352
rect 19064 18275 19116 18284
rect 19064 18241 19073 18275
rect 19073 18241 19107 18275
rect 19107 18241 19116 18275
rect 19064 18232 19116 18241
rect 22284 18232 22336 18284
rect 2228 18207 2280 18216
rect 2228 18173 2237 18207
rect 2237 18173 2271 18207
rect 2271 18173 2280 18207
rect 2228 18164 2280 18173
rect 2780 18207 2832 18216
rect 2780 18173 2789 18207
rect 2789 18173 2823 18207
rect 2823 18173 2832 18207
rect 2780 18164 2832 18173
rect 12716 18207 12768 18216
rect 12716 18173 12725 18207
rect 12725 18173 12759 18207
rect 12759 18173 12768 18207
rect 12716 18164 12768 18173
rect 13360 18164 13412 18216
rect 16028 18207 16080 18216
rect 16028 18173 16037 18207
rect 16037 18173 16071 18207
rect 16071 18173 16080 18207
rect 16028 18164 16080 18173
rect 12624 18096 12676 18148
rect 15200 18028 15252 18080
rect 15844 18096 15896 18148
rect 19340 18164 19392 18216
rect 22376 18164 22428 18216
rect 22928 18275 22980 18284
rect 22928 18241 22937 18275
rect 22937 18241 22971 18275
rect 22971 18241 22980 18275
rect 22928 18232 22980 18241
rect 26332 18232 26384 18284
rect 26608 18275 26660 18284
rect 26608 18241 26617 18275
rect 26617 18241 26651 18275
rect 26651 18241 26660 18275
rect 26608 18232 26660 18241
rect 27344 18232 27396 18284
rect 27712 18275 27764 18284
rect 27712 18241 27721 18275
rect 27721 18241 27755 18275
rect 27755 18241 27764 18275
rect 27712 18232 27764 18241
rect 30104 18300 30156 18352
rect 33876 18300 33928 18352
rect 22652 18096 22704 18148
rect 22744 18096 22796 18148
rect 27528 18164 27580 18216
rect 28172 18232 28224 18284
rect 28632 18275 28684 18284
rect 28632 18241 28641 18275
rect 28641 18241 28675 18275
rect 28675 18241 28684 18275
rect 28632 18232 28684 18241
rect 30288 18232 30340 18284
rect 18696 18071 18748 18080
rect 18696 18037 18705 18071
rect 18705 18037 18739 18071
rect 18739 18037 18748 18071
rect 18696 18028 18748 18037
rect 23572 18028 23624 18080
rect 27252 18028 27304 18080
rect 27988 18096 28040 18148
rect 35900 18300 35952 18352
rect 34060 18232 34112 18284
rect 36452 18275 36504 18284
rect 36452 18241 36461 18275
rect 36461 18241 36495 18275
rect 36495 18241 36504 18275
rect 36452 18232 36504 18241
rect 37188 18300 37240 18352
rect 37004 18232 37056 18284
rect 37556 18232 37608 18284
rect 32956 18207 33008 18216
rect 32956 18173 32965 18207
rect 32965 18173 32999 18207
rect 32999 18173 33008 18207
rect 32956 18164 33008 18173
rect 31760 18139 31812 18148
rect 31760 18105 31769 18139
rect 31769 18105 31803 18139
rect 31803 18105 31812 18139
rect 33140 18207 33192 18216
rect 33140 18173 33149 18207
rect 33149 18173 33183 18207
rect 33183 18173 33192 18207
rect 33140 18164 33192 18173
rect 33324 18164 33376 18216
rect 37924 18232 37976 18284
rect 40592 18300 40644 18352
rect 41696 18300 41748 18352
rect 42616 18368 42668 18420
rect 43812 18411 43864 18420
rect 43812 18377 43821 18411
rect 43821 18377 43855 18411
rect 43855 18377 43864 18411
rect 43812 18368 43864 18377
rect 44456 18368 44508 18420
rect 46480 18368 46532 18420
rect 43996 18300 44048 18352
rect 44640 18300 44692 18352
rect 38752 18232 38804 18284
rect 38936 18275 38988 18284
rect 38936 18241 38945 18275
rect 38945 18241 38979 18275
rect 38979 18241 38988 18275
rect 38936 18232 38988 18241
rect 40684 18275 40736 18284
rect 40684 18241 40718 18275
rect 40718 18241 40736 18275
rect 34152 18139 34204 18148
rect 31760 18096 31812 18105
rect 28540 18028 28592 18080
rect 29000 18028 29052 18080
rect 31852 18028 31904 18080
rect 34152 18105 34161 18139
rect 34161 18105 34195 18139
rect 34195 18105 34204 18139
rect 34152 18096 34204 18105
rect 34888 18096 34940 18148
rect 40684 18232 40736 18241
rect 42064 18232 42116 18284
rect 42616 18275 42668 18284
rect 42616 18241 42625 18275
rect 42625 18241 42659 18275
rect 42659 18241 42668 18275
rect 42616 18232 42668 18241
rect 42984 18275 43036 18284
rect 42984 18241 42993 18275
rect 42993 18241 43027 18275
rect 43027 18241 43036 18275
rect 42984 18232 43036 18241
rect 44364 18232 44416 18284
rect 46572 18232 46624 18284
rect 47676 18232 47728 18284
rect 40408 18207 40460 18216
rect 40408 18173 40417 18207
rect 40417 18173 40451 18207
rect 40451 18173 40460 18207
rect 40408 18164 40460 18173
rect 42708 18164 42760 18216
rect 39672 18096 39724 18148
rect 46756 18096 46808 18148
rect 33324 18028 33376 18080
rect 33968 18071 34020 18080
rect 33968 18037 33977 18071
rect 33977 18037 34011 18071
rect 34011 18037 34020 18071
rect 33968 18028 34020 18037
rect 36636 18028 36688 18080
rect 37280 18028 37332 18080
rect 43260 18028 43312 18080
rect 43444 18028 43496 18080
rect 46664 18028 46716 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 2228 17824 2280 17876
rect 12716 17824 12768 17876
rect 23572 17867 23624 17876
rect 23572 17833 23581 17867
rect 23581 17833 23615 17867
rect 23615 17833 23624 17867
rect 23572 17824 23624 17833
rect 28080 17824 28132 17876
rect 30380 17824 30432 17876
rect 32956 17824 33008 17876
rect 34060 17824 34112 17876
rect 18696 17799 18748 17808
rect 18696 17765 18705 17799
rect 18705 17765 18739 17799
rect 18739 17765 18748 17799
rect 18696 17756 18748 17765
rect 28264 17799 28316 17808
rect 28264 17765 28273 17799
rect 28273 17765 28307 17799
rect 28307 17765 28316 17799
rect 28264 17756 28316 17765
rect 11520 17731 11572 17740
rect 11520 17697 11529 17731
rect 11529 17697 11563 17731
rect 11563 17697 11572 17731
rect 11520 17688 11572 17697
rect 2320 17620 2372 17672
rect 15200 17663 15252 17672
rect 15200 17629 15209 17663
rect 15209 17629 15243 17663
rect 15243 17629 15252 17663
rect 15200 17620 15252 17629
rect 18512 17620 18564 17672
rect 18880 17620 18932 17672
rect 27988 17688 28040 17740
rect 29184 17688 29236 17740
rect 22100 17620 22152 17672
rect 22652 17620 22704 17672
rect 25136 17620 25188 17672
rect 27712 17620 27764 17672
rect 29000 17620 29052 17672
rect 31024 17663 31076 17672
rect 31024 17629 31033 17663
rect 31033 17629 31067 17663
rect 31067 17629 31076 17663
rect 31024 17620 31076 17629
rect 31392 17620 31444 17672
rect 31760 17620 31812 17672
rect 34612 17620 34664 17672
rect 35900 17824 35952 17876
rect 39120 17824 39172 17876
rect 40684 17824 40736 17876
rect 12072 17552 12124 17604
rect 22744 17595 22796 17604
rect 22744 17561 22753 17595
rect 22753 17561 22787 17595
rect 22787 17561 22796 17595
rect 22744 17552 22796 17561
rect 28448 17552 28500 17604
rect 28632 17552 28684 17604
rect 15016 17527 15068 17536
rect 15016 17493 15025 17527
rect 15025 17493 15059 17527
rect 15059 17493 15068 17527
rect 15016 17484 15068 17493
rect 19432 17527 19484 17536
rect 19432 17493 19441 17527
rect 19441 17493 19475 17527
rect 19475 17493 19484 17527
rect 19432 17484 19484 17493
rect 28264 17484 28316 17536
rect 35348 17527 35400 17536
rect 35348 17493 35357 17527
rect 35357 17493 35391 17527
rect 35391 17493 35400 17527
rect 35348 17484 35400 17493
rect 36728 17756 36780 17808
rect 37004 17731 37056 17740
rect 37004 17697 37013 17731
rect 37013 17697 37047 17731
rect 37047 17697 37056 17731
rect 37004 17688 37056 17697
rect 35992 17663 36044 17672
rect 35992 17629 36001 17663
rect 36001 17629 36035 17663
rect 36035 17629 36044 17663
rect 35992 17620 36044 17629
rect 35808 17595 35860 17604
rect 35808 17561 35843 17595
rect 35843 17561 35860 17595
rect 35808 17552 35860 17561
rect 36452 17620 36504 17672
rect 36912 17663 36964 17672
rect 36912 17629 36921 17663
rect 36921 17629 36955 17663
rect 36955 17629 36964 17663
rect 36912 17620 36964 17629
rect 37372 17620 37424 17672
rect 37464 17620 37516 17672
rect 38660 17620 38712 17672
rect 41052 17663 41104 17672
rect 41052 17629 41061 17663
rect 41061 17629 41095 17663
rect 41095 17629 41104 17663
rect 41052 17620 41104 17629
rect 41696 17663 41748 17672
rect 41696 17629 41705 17663
rect 41705 17629 41739 17663
rect 41739 17629 41748 17663
rect 41696 17620 41748 17629
rect 40776 17552 40828 17604
rect 42064 17620 42116 17672
rect 43444 17731 43496 17740
rect 43444 17697 43453 17731
rect 43453 17697 43487 17731
rect 43487 17697 43496 17731
rect 43444 17688 43496 17697
rect 46480 17731 46532 17740
rect 46480 17697 46489 17731
rect 46489 17697 46523 17731
rect 46523 17697 46532 17731
rect 46480 17688 46532 17697
rect 46664 17731 46716 17740
rect 46664 17697 46673 17731
rect 46673 17697 46707 17731
rect 46707 17697 46716 17731
rect 46664 17688 46716 17697
rect 48044 17731 48096 17740
rect 48044 17697 48053 17731
rect 48053 17697 48087 17731
rect 48087 17697 48096 17731
rect 48044 17688 48096 17697
rect 43996 17595 44048 17604
rect 36728 17527 36780 17536
rect 36728 17493 36737 17527
rect 36737 17493 36771 17527
rect 36771 17493 36780 17527
rect 36728 17484 36780 17493
rect 41604 17484 41656 17536
rect 42800 17527 42852 17536
rect 42800 17493 42809 17527
rect 42809 17493 42843 17527
rect 42843 17493 42852 17527
rect 42800 17484 42852 17493
rect 43260 17527 43312 17536
rect 43260 17493 43269 17527
rect 43269 17493 43303 17527
rect 43303 17493 43312 17527
rect 43260 17484 43312 17493
rect 43996 17561 44005 17595
rect 44005 17561 44039 17595
rect 44039 17561 44048 17595
rect 43996 17552 44048 17561
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 12072 17323 12124 17332
rect 12072 17289 12081 17323
rect 12081 17289 12115 17323
rect 12115 17289 12124 17323
rect 12072 17280 12124 17289
rect 19064 17280 19116 17332
rect 26240 17323 26292 17332
rect 26240 17289 26249 17323
rect 26249 17289 26283 17323
rect 26283 17289 26292 17323
rect 26240 17280 26292 17289
rect 11520 17212 11572 17264
rect 13912 17212 13964 17264
rect 12716 17144 12768 17196
rect 13176 17144 13228 17196
rect 15016 17212 15068 17264
rect 19432 17212 19484 17264
rect 23480 17212 23532 17264
rect 30196 17212 30248 17264
rect 18328 17144 18380 17196
rect 22192 17187 22244 17196
rect 22192 17153 22201 17187
rect 22201 17153 22235 17187
rect 22235 17153 22244 17187
rect 22192 17144 22244 17153
rect 22560 17144 22612 17196
rect 23848 17144 23900 17196
rect 24400 17144 24452 17196
rect 26148 17187 26200 17196
rect 14096 17076 14148 17128
rect 18420 17119 18472 17128
rect 18420 17085 18429 17119
rect 18429 17085 18463 17119
rect 18463 17085 18472 17119
rect 18420 17076 18472 17085
rect 25320 17119 25372 17128
rect 1584 16940 1636 16992
rect 22100 17008 22152 17060
rect 22744 17008 22796 17060
rect 25320 17085 25329 17119
rect 25329 17085 25363 17119
rect 25363 17085 25372 17119
rect 25320 17076 25372 17085
rect 26148 17153 26157 17187
rect 26157 17153 26191 17187
rect 26191 17153 26200 17187
rect 26148 17144 26200 17153
rect 30748 17144 30800 17196
rect 34612 17255 34664 17264
rect 34612 17221 34621 17255
rect 34621 17221 34655 17255
rect 34655 17221 34664 17255
rect 34612 17212 34664 17221
rect 34796 17255 34848 17264
rect 34796 17221 34821 17255
rect 34821 17221 34848 17255
rect 34796 17212 34848 17221
rect 30932 17076 30984 17128
rect 33324 17144 33376 17196
rect 34520 17144 34572 17196
rect 35532 17212 35584 17264
rect 35992 17144 36044 17196
rect 39120 17280 39172 17332
rect 41052 17280 41104 17332
rect 43444 17280 43496 17332
rect 37372 17212 37424 17264
rect 36820 17144 36872 17196
rect 39488 17187 39540 17196
rect 33692 17076 33744 17128
rect 26240 17008 26292 17060
rect 27436 17008 27488 17060
rect 33416 17008 33468 17060
rect 15016 16940 15068 16992
rect 16856 16983 16908 16992
rect 16856 16949 16865 16983
rect 16865 16949 16899 16983
rect 16899 16949 16908 16983
rect 16856 16940 16908 16949
rect 22008 16983 22060 16992
rect 22008 16949 22017 16983
rect 22017 16949 22051 16983
rect 22051 16949 22060 16983
rect 22008 16940 22060 16949
rect 22560 16940 22612 16992
rect 24400 16983 24452 16992
rect 24400 16949 24409 16983
rect 24409 16949 24443 16983
rect 24443 16949 24452 16983
rect 24400 16940 24452 16949
rect 24860 16983 24912 16992
rect 24860 16949 24869 16983
rect 24869 16949 24903 16983
rect 24903 16949 24912 16983
rect 24860 16940 24912 16949
rect 32496 16940 32548 16992
rect 34060 17008 34112 17060
rect 34428 16940 34480 16992
rect 34704 16940 34756 16992
rect 36912 17119 36964 17128
rect 35808 16940 35860 16992
rect 36912 17085 36921 17119
rect 36921 17085 36955 17119
rect 36955 17085 36964 17119
rect 36912 17076 36964 17085
rect 37464 17119 37516 17128
rect 37464 17085 37473 17119
rect 37473 17085 37507 17119
rect 37507 17085 37516 17119
rect 37464 17076 37516 17085
rect 39488 17153 39497 17187
rect 39497 17153 39531 17187
rect 39531 17153 39540 17187
rect 39488 17144 39540 17153
rect 41604 17187 41656 17196
rect 41604 17153 41613 17187
rect 41613 17153 41647 17187
rect 41647 17153 41656 17187
rect 41604 17144 41656 17153
rect 42892 17144 42944 17196
rect 44364 17212 44416 17264
rect 47124 17212 47176 17264
rect 39948 17076 40000 17128
rect 43260 17076 43312 17128
rect 42708 17008 42760 17060
rect 43628 17144 43680 17196
rect 46388 17076 46440 17128
rect 46848 17119 46900 17128
rect 46848 17085 46857 17119
rect 46857 17085 46891 17119
rect 46891 17085 46900 17119
rect 46848 17076 46900 17085
rect 37648 16940 37700 16992
rect 43812 16940 43864 16992
rect 44180 16940 44232 16992
rect 46480 16940 46532 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 12716 16779 12768 16788
rect 12716 16745 12725 16779
rect 12725 16745 12759 16779
rect 12759 16745 12768 16779
rect 12716 16736 12768 16745
rect 1584 16643 1636 16652
rect 1584 16609 1593 16643
rect 1593 16609 1627 16643
rect 1627 16609 1636 16643
rect 1584 16600 1636 16609
rect 2780 16643 2832 16652
rect 2780 16609 2789 16643
rect 2789 16609 2823 16643
rect 2823 16609 2832 16643
rect 2780 16600 2832 16609
rect 13176 16643 13228 16652
rect 13176 16609 13185 16643
rect 13185 16609 13219 16643
rect 13219 16609 13228 16643
rect 13176 16600 13228 16609
rect 13360 16643 13412 16652
rect 13360 16609 13369 16643
rect 13369 16609 13403 16643
rect 13403 16609 13412 16643
rect 13360 16600 13412 16609
rect 16764 16736 16816 16788
rect 18420 16668 18472 16720
rect 22100 16736 22152 16788
rect 23480 16779 23532 16788
rect 23480 16745 23489 16779
rect 23489 16745 23523 16779
rect 23523 16745 23532 16779
rect 23480 16736 23532 16745
rect 26148 16736 26200 16788
rect 27620 16736 27672 16788
rect 30288 16736 30340 16788
rect 24492 16600 24544 16652
rect 26332 16668 26384 16720
rect 22008 16532 22060 16584
rect 24860 16532 24912 16584
rect 25228 16643 25280 16652
rect 25228 16609 25237 16643
rect 25237 16609 25271 16643
rect 25271 16609 25280 16643
rect 25228 16600 25280 16609
rect 25780 16600 25832 16652
rect 25964 16600 26016 16652
rect 30288 16643 30340 16652
rect 30288 16609 30297 16643
rect 30297 16609 30331 16643
rect 30331 16609 30340 16643
rect 30288 16600 30340 16609
rect 34704 16736 34756 16788
rect 35532 16736 35584 16788
rect 36728 16779 36780 16788
rect 36728 16745 36737 16779
rect 36737 16745 36771 16779
rect 36771 16745 36780 16779
rect 36728 16736 36780 16745
rect 36820 16779 36872 16788
rect 36820 16745 36829 16779
rect 36829 16745 36863 16779
rect 36863 16745 36872 16779
rect 36820 16736 36872 16745
rect 43628 16736 43680 16788
rect 33324 16668 33376 16720
rect 35072 16668 35124 16720
rect 38292 16711 38344 16720
rect 2596 16464 2648 16516
rect 16856 16464 16908 16516
rect 17500 16396 17552 16448
rect 22652 16396 22704 16448
rect 25320 16464 25372 16516
rect 24952 16439 25004 16448
rect 24952 16405 24961 16439
rect 24961 16405 24995 16439
rect 24995 16405 25004 16439
rect 24952 16396 25004 16405
rect 26700 16532 26752 16584
rect 27068 16575 27120 16584
rect 27068 16541 27077 16575
rect 27077 16541 27111 16575
rect 27111 16541 27120 16575
rect 27068 16532 27120 16541
rect 27252 16575 27304 16584
rect 27252 16541 27261 16575
rect 27261 16541 27295 16575
rect 27295 16541 27304 16575
rect 27252 16532 27304 16541
rect 27344 16575 27396 16584
rect 27344 16541 27353 16575
rect 27353 16541 27387 16575
rect 27387 16541 27396 16575
rect 27344 16532 27396 16541
rect 35348 16600 35400 16652
rect 26056 16507 26108 16516
rect 26056 16473 26065 16507
rect 26065 16473 26099 16507
rect 26099 16473 26108 16507
rect 26056 16464 26108 16473
rect 26424 16464 26476 16516
rect 26516 16464 26568 16516
rect 34796 16532 34848 16584
rect 35716 16575 35768 16584
rect 28264 16464 28316 16516
rect 30564 16507 30616 16516
rect 30564 16473 30598 16507
rect 30598 16473 30616 16507
rect 30564 16464 30616 16473
rect 32404 16507 32456 16516
rect 32404 16473 32438 16507
rect 32438 16473 32456 16507
rect 32404 16464 32456 16473
rect 34704 16464 34756 16516
rect 35072 16507 35124 16516
rect 28172 16439 28224 16448
rect 28172 16405 28181 16439
rect 28181 16405 28215 16439
rect 28215 16405 28224 16439
rect 28172 16396 28224 16405
rect 31484 16396 31536 16448
rect 33324 16396 33376 16448
rect 34152 16439 34204 16448
rect 34152 16405 34167 16439
rect 34167 16405 34201 16439
rect 34201 16405 34204 16439
rect 34152 16396 34204 16405
rect 34520 16396 34572 16448
rect 35072 16473 35081 16507
rect 35081 16473 35115 16507
rect 35115 16473 35124 16507
rect 35072 16464 35124 16473
rect 35716 16541 35725 16575
rect 35725 16541 35759 16575
rect 35759 16541 35768 16575
rect 35716 16532 35768 16541
rect 38292 16677 38301 16711
rect 38301 16677 38335 16711
rect 38335 16677 38344 16711
rect 38292 16668 38344 16677
rect 44548 16668 44600 16720
rect 37280 16600 37332 16652
rect 37464 16600 37516 16652
rect 40408 16600 40460 16652
rect 40776 16600 40828 16652
rect 36636 16575 36688 16584
rect 36636 16541 36645 16575
rect 36645 16541 36679 16575
rect 36679 16541 36688 16575
rect 36636 16532 36688 16541
rect 37372 16532 37424 16584
rect 39488 16532 39540 16584
rect 41788 16600 41840 16652
rect 46480 16643 46532 16652
rect 46480 16609 46489 16643
rect 46489 16609 46523 16643
rect 46523 16609 46532 16643
rect 46480 16600 46532 16609
rect 48228 16643 48280 16652
rect 48228 16609 48237 16643
rect 48237 16609 48271 16643
rect 48271 16609 48280 16643
rect 48228 16600 48280 16609
rect 42800 16532 42852 16584
rect 46756 16464 46808 16516
rect 35716 16396 35768 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 2596 16235 2648 16244
rect 2596 16201 2605 16235
rect 2605 16201 2639 16235
rect 2639 16201 2648 16235
rect 2596 16192 2648 16201
rect 13176 16192 13228 16244
rect 17500 16235 17552 16244
rect 17040 16124 17092 16176
rect 17500 16201 17509 16235
rect 17509 16201 17543 16235
rect 17543 16201 17552 16235
rect 17500 16192 17552 16201
rect 18420 16192 18472 16244
rect 22192 16192 22244 16244
rect 26332 16192 26384 16244
rect 26424 16192 26476 16244
rect 2412 16056 2464 16108
rect 12164 16056 12216 16108
rect 12900 16056 12952 16108
rect 15200 16056 15252 16108
rect 18604 16056 18656 16108
rect 18880 16056 18932 16108
rect 22192 16099 22244 16108
rect 22192 16065 22201 16099
rect 22201 16065 22235 16099
rect 22235 16065 22244 16099
rect 22192 16056 22244 16065
rect 22468 16099 22520 16108
rect 22468 16065 22477 16099
rect 22477 16065 22511 16099
rect 22511 16065 22520 16099
rect 22468 16056 22520 16065
rect 22652 16099 22704 16108
rect 22652 16065 22661 16099
rect 22661 16065 22695 16099
rect 22695 16065 22704 16099
rect 24952 16124 25004 16176
rect 24400 16099 24452 16108
rect 22652 16056 22704 16065
rect 24400 16065 24409 16099
rect 24409 16065 24443 16099
rect 24443 16065 24452 16099
rect 24400 16056 24452 16065
rect 24584 16099 24636 16108
rect 24584 16065 24593 16099
rect 24593 16065 24627 16099
rect 24627 16065 24636 16099
rect 24584 16056 24636 16065
rect 24768 16056 24820 16108
rect 13360 15988 13412 16040
rect 15108 15988 15160 16040
rect 17592 16031 17644 16040
rect 17592 15997 17601 16031
rect 17601 15997 17635 16031
rect 17635 15997 17644 16031
rect 17592 15988 17644 15997
rect 17684 16031 17736 16040
rect 17684 15997 17693 16031
rect 17693 15997 17727 16031
rect 17727 15997 17736 16031
rect 17684 15988 17736 15997
rect 26240 16056 26292 16108
rect 28172 16124 28224 16176
rect 27528 16099 27580 16108
rect 27528 16065 27537 16099
rect 27537 16065 27571 16099
rect 27571 16065 27580 16099
rect 27528 16056 27580 16065
rect 31024 16099 31076 16108
rect 25964 16031 26016 16040
rect 25964 15997 25973 16031
rect 25973 15997 26007 16031
rect 26007 15997 26016 16031
rect 25964 15988 26016 15997
rect 27620 16031 27672 16040
rect 24768 15920 24820 15972
rect 27620 15997 27629 16031
rect 27629 15997 27663 16031
rect 27663 15997 27672 16031
rect 27620 15988 27672 15997
rect 27068 15920 27120 15972
rect 31024 16065 31033 16099
rect 31033 16065 31067 16099
rect 31067 16065 31076 16099
rect 31024 16056 31076 16065
rect 31392 16124 31444 16176
rect 32404 16192 32456 16244
rect 34704 16167 34756 16176
rect 34704 16133 34713 16167
rect 34713 16133 34747 16167
rect 34747 16133 34756 16167
rect 34704 16124 34756 16133
rect 35348 16192 35400 16244
rect 41604 16192 41656 16244
rect 47124 16235 47176 16244
rect 47124 16201 47133 16235
rect 47133 16201 47167 16235
rect 47167 16201 47176 16235
rect 47124 16192 47176 16201
rect 39488 16124 39540 16176
rect 31484 16099 31536 16108
rect 31484 16065 31493 16099
rect 31493 16065 31527 16099
rect 31527 16065 31536 16099
rect 32496 16099 32548 16108
rect 31484 16056 31536 16065
rect 27988 16031 28040 16040
rect 27988 15997 27997 16031
rect 27997 15997 28031 16031
rect 28031 15997 28040 16031
rect 27988 15988 28040 15997
rect 13084 15852 13136 15904
rect 19156 15895 19208 15904
rect 19156 15861 19165 15895
rect 19165 15861 19199 15895
rect 19199 15861 19208 15895
rect 19156 15852 19208 15861
rect 26424 15852 26476 15904
rect 26792 15852 26844 15904
rect 30472 15920 30524 15972
rect 32496 16065 32505 16099
rect 32505 16065 32539 16099
rect 32539 16065 32548 16099
rect 32496 16056 32548 16065
rect 32680 16099 32732 16108
rect 32680 16065 32689 16099
rect 32689 16065 32723 16099
rect 32723 16065 32732 16099
rect 32680 16056 32732 16065
rect 33324 16056 33376 16108
rect 33416 16099 33468 16108
rect 33416 16065 33425 16099
rect 33425 16065 33459 16099
rect 33459 16065 33468 16099
rect 33416 16056 33468 16065
rect 33600 16099 33652 16108
rect 33600 16065 33609 16099
rect 33609 16065 33643 16099
rect 33643 16065 33652 16099
rect 33600 16056 33652 16065
rect 34152 16056 34204 16108
rect 39304 16056 39356 16108
rect 39764 16031 39816 16040
rect 30656 15852 30708 15904
rect 33232 15895 33284 15904
rect 33232 15861 33241 15895
rect 33241 15861 33275 15895
rect 33275 15861 33284 15895
rect 33232 15852 33284 15861
rect 34796 15852 34848 15904
rect 35716 15895 35768 15904
rect 35716 15861 35725 15895
rect 35725 15861 35759 15895
rect 35759 15861 35768 15895
rect 39764 15997 39773 16031
rect 39773 15997 39807 16031
rect 39807 15997 39816 16031
rect 39764 15988 39816 15997
rect 41880 16124 41932 16176
rect 41788 16099 41840 16108
rect 41788 16065 41797 16099
rect 41797 16065 41831 16099
rect 41831 16065 41840 16099
rect 41788 16056 41840 16065
rect 46940 16056 46992 16108
rect 46388 15988 46440 16040
rect 42064 15920 42116 15972
rect 35716 15852 35768 15861
rect 40132 15852 40184 15904
rect 41696 15895 41748 15904
rect 41696 15861 41705 15895
rect 41705 15861 41739 15895
rect 41739 15861 41748 15895
rect 41696 15852 41748 15861
rect 41972 15852 42024 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 12900 15691 12952 15700
rect 12900 15657 12909 15691
rect 12909 15657 12943 15691
rect 12943 15657 12952 15691
rect 12900 15648 12952 15657
rect 18880 15691 18932 15700
rect 18880 15657 18889 15691
rect 18889 15657 18923 15691
rect 18923 15657 18932 15691
rect 18880 15648 18932 15657
rect 26240 15691 26292 15700
rect 17500 15580 17552 15632
rect 26240 15657 26249 15691
rect 26249 15657 26283 15691
rect 26283 15657 26292 15691
rect 26240 15648 26292 15657
rect 27068 15580 27120 15632
rect 2780 15555 2832 15564
rect 2780 15521 2789 15555
rect 2789 15521 2823 15555
rect 2823 15521 2832 15555
rect 2780 15512 2832 15521
rect 15016 15555 15068 15564
rect 15016 15521 15025 15555
rect 15025 15521 15059 15555
rect 15059 15521 15068 15555
rect 15016 15512 15068 15521
rect 15108 15555 15160 15564
rect 15108 15521 15117 15555
rect 15117 15521 15151 15555
rect 15151 15521 15160 15555
rect 17684 15555 17736 15564
rect 15108 15512 15160 15521
rect 17684 15521 17693 15555
rect 17693 15521 17727 15555
rect 17727 15521 17736 15555
rect 17684 15512 17736 15521
rect 19340 15512 19392 15564
rect 22100 15512 22152 15564
rect 24768 15512 24820 15564
rect 1584 15487 1636 15496
rect 1584 15453 1593 15487
rect 1593 15453 1627 15487
rect 1627 15453 1636 15487
rect 1584 15444 1636 15453
rect 13084 15487 13136 15496
rect 13084 15453 13093 15487
rect 13093 15453 13127 15487
rect 13127 15453 13136 15487
rect 13084 15444 13136 15453
rect 1952 15376 2004 15428
rect 2412 15376 2464 15428
rect 2872 15308 2924 15360
rect 14096 15308 14148 15360
rect 17040 15444 17092 15496
rect 17408 15487 17460 15496
rect 17408 15453 17417 15487
rect 17417 15453 17451 15487
rect 17451 15453 17460 15487
rect 17408 15444 17460 15453
rect 17132 15308 17184 15360
rect 17500 15351 17552 15360
rect 17500 15317 17509 15351
rect 17509 15317 17543 15351
rect 17543 15317 17552 15351
rect 17500 15308 17552 15317
rect 18604 15376 18656 15428
rect 19984 15376 20036 15428
rect 23204 15376 23256 15428
rect 24584 15444 24636 15496
rect 26516 15512 26568 15564
rect 26424 15487 26476 15496
rect 26424 15453 26433 15487
rect 26433 15453 26467 15487
rect 26467 15453 26476 15487
rect 26424 15444 26476 15453
rect 27252 15512 27304 15564
rect 27068 15487 27120 15496
rect 27068 15453 27077 15487
rect 27077 15453 27111 15487
rect 27111 15453 27120 15487
rect 27068 15444 27120 15453
rect 30564 15648 30616 15700
rect 30840 15691 30892 15700
rect 30840 15657 30849 15691
rect 30849 15657 30883 15691
rect 30883 15657 30892 15691
rect 30840 15648 30892 15657
rect 39304 15691 39356 15700
rect 39304 15657 39313 15691
rect 39313 15657 39347 15691
rect 39347 15657 39356 15691
rect 39304 15648 39356 15657
rect 40776 15648 40828 15700
rect 42708 15648 42760 15700
rect 28264 15580 28316 15632
rect 30932 15555 30984 15564
rect 30932 15521 30941 15555
rect 30941 15521 30975 15555
rect 30975 15521 30984 15555
rect 30932 15512 30984 15521
rect 26792 15376 26844 15428
rect 27344 15376 27396 15428
rect 28632 15444 28684 15496
rect 30656 15487 30708 15496
rect 30656 15453 30665 15487
rect 30665 15453 30699 15487
rect 30699 15453 30708 15487
rect 30656 15444 30708 15453
rect 33232 15444 33284 15496
rect 35716 15512 35768 15564
rect 37096 15444 37148 15496
rect 40776 15555 40828 15564
rect 40776 15521 40785 15555
rect 40785 15521 40819 15555
rect 40819 15521 40828 15555
rect 40776 15512 40828 15521
rect 41788 15555 41840 15564
rect 41788 15521 41797 15555
rect 41797 15521 41831 15555
rect 41831 15521 41840 15555
rect 41788 15512 41840 15521
rect 41880 15555 41932 15564
rect 41880 15521 41889 15555
rect 41889 15521 41923 15555
rect 41923 15521 41932 15555
rect 42708 15555 42760 15564
rect 41880 15512 41932 15521
rect 42708 15521 42717 15555
rect 42717 15521 42751 15555
rect 42751 15521 42760 15555
rect 42708 15512 42760 15521
rect 47952 15512 48004 15564
rect 48228 15555 48280 15564
rect 48228 15521 48237 15555
rect 48237 15521 48271 15555
rect 48271 15521 48280 15555
rect 48228 15512 48280 15521
rect 38936 15444 38988 15496
rect 40500 15444 40552 15496
rect 41604 15487 41656 15496
rect 41604 15453 41613 15487
rect 41613 15453 41647 15487
rect 41647 15453 41656 15487
rect 41604 15444 41656 15453
rect 41972 15444 42024 15496
rect 23664 15308 23716 15360
rect 24584 15308 24636 15360
rect 26700 15308 26752 15360
rect 29276 15376 29328 15428
rect 34520 15376 34572 15428
rect 35716 15376 35768 15428
rect 40040 15419 40092 15428
rect 40040 15385 40049 15419
rect 40049 15385 40083 15419
rect 40083 15385 40092 15419
rect 40040 15376 40092 15385
rect 43076 15376 43128 15428
rect 47124 15376 47176 15428
rect 28540 15308 28592 15360
rect 35440 15351 35492 15360
rect 35440 15317 35449 15351
rect 35449 15317 35483 15351
rect 35483 15317 35492 15351
rect 35440 15308 35492 15317
rect 37372 15308 37424 15360
rect 38936 15308 38988 15360
rect 41420 15351 41472 15360
rect 41420 15317 41429 15351
rect 41429 15317 41463 15351
rect 41463 15317 41472 15351
rect 44088 15351 44140 15360
rect 41420 15308 41472 15317
rect 44088 15317 44097 15351
rect 44097 15317 44131 15351
rect 44131 15317 44140 15351
rect 44088 15308 44140 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 2872 15147 2924 15156
rect 2872 15113 2881 15147
rect 2881 15113 2915 15147
rect 2915 15113 2924 15147
rect 2872 15104 2924 15113
rect 15200 15147 15252 15156
rect 15200 15113 15209 15147
rect 15209 15113 15243 15147
rect 15243 15113 15252 15147
rect 15200 15104 15252 15113
rect 1584 14968 1636 15020
rect 2504 14968 2556 15020
rect 3240 14968 3292 15020
rect 4620 15036 4672 15088
rect 14096 15079 14148 15088
rect 14096 15045 14130 15079
rect 14130 15045 14148 15079
rect 14096 15036 14148 15045
rect 13912 14968 13964 15020
rect 19984 15104 20036 15156
rect 27160 15104 27212 15156
rect 35716 15147 35768 15156
rect 35716 15113 35725 15147
rect 35725 15113 35759 15147
rect 35759 15113 35768 15147
rect 35716 15104 35768 15113
rect 41420 15104 41472 15156
rect 43076 15147 43128 15156
rect 43076 15113 43085 15147
rect 43085 15113 43119 15147
rect 43119 15113 43128 15147
rect 43076 15104 43128 15113
rect 47124 15147 47176 15156
rect 18604 15036 18656 15088
rect 19156 15036 19208 15088
rect 16764 14968 16816 15020
rect 23020 14968 23072 15020
rect 23848 15011 23900 15020
rect 4068 14900 4120 14952
rect 5356 14943 5408 14952
rect 5356 14909 5365 14943
rect 5365 14909 5399 14943
rect 5399 14909 5408 14943
rect 5356 14900 5408 14909
rect 23112 14900 23164 14952
rect 23848 14977 23857 15011
rect 23857 14977 23891 15011
rect 23891 14977 23900 15011
rect 23848 14968 23900 14977
rect 26332 14900 26384 14952
rect 27252 14968 27304 15020
rect 29092 15036 29144 15088
rect 30288 15036 30340 15088
rect 30380 15036 30432 15088
rect 29000 15011 29052 15020
rect 29000 14977 29034 15011
rect 29034 14977 29052 15011
rect 32680 15011 32732 15020
rect 29000 14968 29052 14977
rect 32680 14977 32689 15011
rect 32689 14977 32723 15011
rect 32723 14977 32732 15011
rect 32680 14968 32732 14977
rect 35440 15036 35492 15088
rect 37372 15036 37424 15088
rect 40224 15036 40276 15088
rect 42800 15036 42852 15088
rect 47124 15113 47133 15147
rect 47133 15113 47167 15147
rect 47167 15113 47176 15147
rect 47124 15104 47176 15113
rect 37464 15011 37516 15020
rect 37464 14977 37473 15011
rect 37473 14977 37507 15011
rect 37507 14977 37516 15011
rect 37464 14968 37516 14977
rect 17132 14875 17184 14884
rect 17132 14841 17141 14875
rect 17141 14841 17175 14875
rect 17175 14841 17184 14875
rect 17132 14832 17184 14841
rect 32772 14900 32824 14952
rect 30288 14832 30340 14884
rect 33692 14832 33744 14884
rect 16120 14807 16172 14816
rect 16120 14773 16129 14807
rect 16129 14773 16163 14807
rect 16163 14773 16172 14807
rect 16120 14764 16172 14773
rect 23388 14764 23440 14816
rect 28724 14764 28776 14816
rect 32588 14764 32640 14816
rect 38200 14764 38252 14816
rect 41696 14832 41748 14884
rect 43444 15011 43496 15020
rect 43444 14977 43453 15011
rect 43453 14977 43487 15011
rect 43487 14977 43496 15011
rect 43444 14968 43496 14977
rect 43720 15011 43772 15020
rect 43720 14977 43729 15011
rect 43729 14977 43763 15011
rect 43763 14977 43772 15011
rect 43720 14968 43772 14977
rect 44088 14968 44140 15020
rect 44180 15011 44232 15020
rect 44180 14977 44189 15011
rect 44189 14977 44223 15011
rect 44223 14977 44232 15011
rect 47032 15011 47084 15020
rect 44180 14968 44232 14977
rect 47032 14977 47041 15011
rect 47041 14977 47075 15011
rect 47075 14977 47084 15011
rect 47032 14968 47084 14977
rect 47952 15011 48004 15020
rect 47952 14977 47961 15011
rect 47961 14977 47995 15011
rect 47995 14977 48004 15011
rect 47952 14968 48004 14977
rect 44364 14900 44416 14952
rect 44456 14943 44508 14952
rect 44456 14909 44465 14943
rect 44465 14909 44499 14943
rect 44499 14909 44508 14943
rect 44456 14900 44508 14909
rect 40500 14807 40552 14816
rect 40500 14773 40509 14807
rect 40509 14773 40543 14807
rect 40543 14773 40552 14807
rect 40500 14764 40552 14773
rect 44272 14807 44324 14816
rect 44272 14773 44281 14807
rect 44281 14773 44315 14807
rect 44315 14773 44324 14807
rect 44272 14764 44324 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 4068 14603 4120 14612
rect 4068 14569 4077 14603
rect 4077 14569 4111 14603
rect 4111 14569 4120 14603
rect 4068 14560 4120 14569
rect 17408 14603 17460 14612
rect 17408 14569 17417 14603
rect 17417 14569 17451 14603
rect 17451 14569 17460 14603
rect 17408 14560 17460 14569
rect 23204 14603 23256 14612
rect 23204 14569 23213 14603
rect 23213 14569 23247 14603
rect 23247 14569 23256 14603
rect 23204 14560 23256 14569
rect 25044 14603 25096 14612
rect 25044 14569 25053 14603
rect 25053 14569 25087 14603
rect 25087 14569 25096 14603
rect 25044 14560 25096 14569
rect 27068 14560 27120 14612
rect 29000 14560 29052 14612
rect 29276 14560 29328 14612
rect 38936 14603 38988 14612
rect 22560 14492 22612 14544
rect 23020 14492 23072 14544
rect 2780 14467 2832 14476
rect 2780 14433 2789 14467
rect 2789 14433 2823 14467
rect 2823 14433 2832 14467
rect 2780 14424 2832 14433
rect 23664 14467 23716 14476
rect 23664 14433 23673 14467
rect 23673 14433 23707 14467
rect 23707 14433 23716 14467
rect 23664 14424 23716 14433
rect 27804 14492 27856 14544
rect 29828 14424 29880 14476
rect 30104 14535 30156 14544
rect 30104 14501 30113 14535
rect 30113 14501 30147 14535
rect 30147 14501 30156 14535
rect 30104 14492 30156 14501
rect 30380 14492 30432 14544
rect 38936 14569 38945 14603
rect 38945 14569 38979 14603
rect 38979 14569 38988 14603
rect 38936 14560 38988 14569
rect 41972 14560 42024 14612
rect 44272 14603 44324 14612
rect 44272 14569 44281 14603
rect 44281 14569 44315 14603
rect 44315 14569 44324 14603
rect 44272 14560 44324 14569
rect 44364 14560 44416 14612
rect 37924 14492 37976 14544
rect 33692 14467 33744 14476
rect 1584 14399 1636 14408
rect 1584 14365 1593 14399
rect 1593 14365 1627 14399
rect 1627 14365 1636 14399
rect 1584 14356 1636 14365
rect 3792 14356 3844 14408
rect 16764 14356 16816 14408
rect 23388 14399 23440 14408
rect 23388 14365 23397 14399
rect 23397 14365 23431 14399
rect 23431 14365 23440 14399
rect 23388 14356 23440 14365
rect 24860 14399 24912 14408
rect 24860 14365 24869 14399
rect 24869 14365 24903 14399
rect 24903 14365 24912 14399
rect 24860 14356 24912 14365
rect 25688 14356 25740 14408
rect 27252 14356 27304 14408
rect 1768 14331 1820 14340
rect 1768 14297 1777 14331
rect 1777 14297 1811 14331
rect 1811 14297 1820 14331
rect 1768 14288 1820 14297
rect 16120 14288 16172 14340
rect 26332 14331 26384 14340
rect 26332 14297 26341 14331
rect 26341 14297 26375 14331
rect 26375 14297 26384 14331
rect 26332 14288 26384 14297
rect 24584 14220 24636 14272
rect 27252 14220 27304 14272
rect 27712 14356 27764 14408
rect 28540 14399 28592 14408
rect 28540 14365 28549 14399
rect 28549 14365 28583 14399
rect 28583 14365 28592 14399
rect 28540 14356 28592 14365
rect 28724 14399 28776 14408
rect 28724 14365 28731 14399
rect 28731 14365 28776 14399
rect 28724 14356 28776 14365
rect 29276 14356 29328 14408
rect 31484 14399 31536 14408
rect 27620 14220 27672 14272
rect 28908 14331 28960 14340
rect 28908 14297 28917 14331
rect 28917 14297 28951 14331
rect 28951 14297 28960 14331
rect 28908 14288 28960 14297
rect 29828 14288 29880 14340
rect 31484 14365 31493 14399
rect 31493 14365 31527 14399
rect 31527 14365 31536 14399
rect 31484 14356 31536 14365
rect 31576 14356 31628 14408
rect 33692 14433 33701 14467
rect 33701 14433 33735 14467
rect 33735 14433 33744 14467
rect 33692 14424 33744 14433
rect 43720 14424 43772 14476
rect 31944 14356 31996 14408
rect 32496 14356 32548 14408
rect 38200 14356 38252 14408
rect 38752 14399 38804 14408
rect 38752 14365 38761 14399
rect 38761 14365 38795 14399
rect 38795 14365 38804 14399
rect 38752 14356 38804 14365
rect 38936 14356 38988 14408
rect 42892 14356 42944 14408
rect 44180 14424 44232 14476
rect 44272 14399 44324 14408
rect 44272 14365 44281 14399
rect 44281 14365 44315 14399
rect 44315 14365 44324 14399
rect 44272 14356 44324 14365
rect 44456 14356 44508 14408
rect 30012 14220 30064 14272
rect 30288 14288 30340 14340
rect 37188 14288 37240 14340
rect 40776 14331 40828 14340
rect 40776 14297 40785 14331
rect 40785 14297 40819 14331
rect 40819 14297 40828 14331
rect 40776 14288 40828 14297
rect 30380 14220 30432 14272
rect 32036 14263 32088 14272
rect 32036 14229 32045 14263
rect 32045 14229 32079 14263
rect 32079 14229 32088 14263
rect 32036 14220 32088 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 1768 14016 1820 14068
rect 25688 14059 25740 14068
rect 25688 14025 25697 14059
rect 25697 14025 25731 14059
rect 25731 14025 25740 14059
rect 25688 14016 25740 14025
rect 28264 14016 28316 14068
rect 28908 14016 28960 14068
rect 31024 14016 31076 14068
rect 31576 14016 31628 14068
rect 38016 14016 38068 14068
rect 40776 14059 40828 14068
rect 40776 14025 40785 14059
rect 40785 14025 40819 14059
rect 40819 14025 40828 14059
rect 40776 14016 40828 14025
rect 44180 14016 44232 14068
rect 45468 14016 45520 14068
rect 1584 13880 1636 13932
rect 2964 13880 3016 13932
rect 22560 13948 22612 14000
rect 22192 13923 22244 13932
rect 22192 13889 22201 13923
rect 22201 13889 22235 13923
rect 22235 13889 22244 13923
rect 22192 13880 22244 13889
rect 22468 13923 22520 13932
rect 22468 13889 22477 13923
rect 22477 13889 22511 13923
rect 22511 13889 22520 13923
rect 22468 13880 22520 13889
rect 22652 13923 22704 13932
rect 22652 13889 22661 13923
rect 22661 13889 22695 13923
rect 22695 13889 22704 13923
rect 22652 13880 22704 13889
rect 23296 13812 23348 13864
rect 20996 13719 21048 13728
rect 20996 13685 21005 13719
rect 21005 13685 21039 13719
rect 21039 13685 21048 13719
rect 20996 13676 21048 13685
rect 24584 13923 24636 13932
rect 24584 13889 24618 13923
rect 24618 13889 24636 13923
rect 24584 13880 24636 13889
rect 25780 13880 25832 13932
rect 29092 13948 29144 14000
rect 30012 13991 30064 14000
rect 30012 13957 30046 13991
rect 30046 13957 30064 13991
rect 30012 13948 30064 13957
rect 32588 13991 32640 14000
rect 32588 13957 32622 13991
rect 32622 13957 32640 13991
rect 32588 13948 32640 13957
rect 27252 13880 27304 13932
rect 37556 13880 37608 13932
rect 39764 13948 39816 14000
rect 40868 13948 40920 14000
rect 41512 13948 41564 14000
rect 40132 13880 40184 13932
rect 40224 13880 40276 13932
rect 41604 13923 41656 13932
rect 26516 13855 26568 13864
rect 26516 13821 26525 13855
rect 26525 13821 26559 13855
rect 26559 13821 26568 13855
rect 26516 13812 26568 13821
rect 32312 13855 32364 13864
rect 32312 13821 32321 13855
rect 32321 13821 32355 13855
rect 32355 13821 32364 13855
rect 32312 13812 32364 13821
rect 41604 13889 41613 13923
rect 41613 13889 41647 13923
rect 41647 13889 41656 13923
rect 41604 13880 41656 13889
rect 41972 13880 42024 13932
rect 42892 13880 42944 13932
rect 43720 13923 43772 13932
rect 41788 13812 41840 13864
rect 43720 13889 43729 13923
rect 43729 13889 43763 13923
rect 43763 13889 43772 13923
rect 43720 13880 43772 13889
rect 43628 13812 43680 13864
rect 43536 13744 43588 13796
rect 45744 13880 45796 13932
rect 47032 13923 47084 13932
rect 47032 13889 47041 13923
rect 47041 13889 47075 13923
rect 47075 13889 47084 13923
rect 47032 13880 47084 13889
rect 44640 13812 44692 13864
rect 45100 13812 45152 13864
rect 33784 13676 33836 13728
rect 43628 13676 43680 13728
rect 47124 13719 47176 13728
rect 47124 13685 47133 13719
rect 47133 13685 47167 13719
rect 47167 13685 47176 13719
rect 47124 13676 47176 13685
rect 47952 13719 48004 13728
rect 47952 13685 47961 13719
rect 47961 13685 47995 13719
rect 47995 13685 48004 13719
rect 47952 13676 48004 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 21548 13472 21600 13524
rect 22652 13472 22704 13524
rect 23020 13515 23072 13524
rect 23020 13481 23029 13515
rect 23029 13481 23063 13515
rect 23063 13481 23072 13515
rect 23020 13472 23072 13481
rect 24860 13472 24912 13524
rect 27620 13515 27672 13524
rect 27620 13481 27629 13515
rect 27629 13481 27663 13515
rect 27663 13481 27672 13515
rect 27620 13472 27672 13481
rect 30380 13515 30432 13524
rect 30380 13481 30389 13515
rect 30389 13481 30423 13515
rect 30423 13481 30432 13515
rect 30380 13472 30432 13481
rect 32680 13472 32732 13524
rect 33600 13472 33652 13524
rect 37556 13515 37608 13524
rect 37556 13481 37565 13515
rect 37565 13481 37599 13515
rect 37599 13481 37608 13515
rect 37556 13472 37608 13481
rect 40408 13472 40460 13524
rect 43352 13472 43404 13524
rect 45744 13515 45796 13524
rect 45744 13481 45753 13515
rect 45753 13481 45787 13515
rect 45787 13481 45796 13515
rect 45744 13472 45796 13481
rect 22468 13404 22520 13456
rect 22836 13311 22888 13320
rect 20720 13132 20772 13184
rect 20996 13200 21048 13252
rect 22836 13277 22845 13311
rect 22845 13277 22879 13311
rect 22879 13277 22888 13311
rect 22836 13268 22888 13277
rect 22928 13268 22980 13320
rect 23204 13336 23256 13388
rect 24952 13311 25004 13320
rect 24952 13277 24961 13311
rect 24961 13277 24995 13311
rect 24995 13277 25004 13311
rect 24952 13268 25004 13277
rect 25412 13311 25464 13320
rect 24860 13200 24912 13252
rect 25412 13277 25421 13311
rect 25421 13277 25455 13311
rect 25455 13277 25464 13311
rect 25412 13268 25464 13277
rect 27712 13268 27764 13320
rect 28264 13311 28316 13320
rect 28264 13277 28273 13311
rect 28273 13277 28307 13311
rect 28307 13277 28316 13311
rect 28264 13268 28316 13277
rect 28356 13200 28408 13252
rect 30748 13268 30800 13320
rect 31024 13311 31076 13320
rect 31024 13277 31033 13311
rect 31033 13277 31067 13311
rect 31067 13277 31076 13311
rect 31024 13268 31076 13277
rect 32496 13336 32548 13388
rect 40040 13336 40092 13388
rect 40868 13379 40920 13388
rect 31116 13200 31168 13252
rect 33416 13268 33468 13320
rect 33784 13311 33836 13320
rect 33784 13277 33793 13311
rect 33793 13277 33827 13311
rect 33827 13277 33836 13311
rect 33784 13268 33836 13277
rect 36820 13268 36872 13320
rect 37096 13268 37148 13320
rect 38016 13311 38068 13320
rect 38016 13277 38025 13311
rect 38025 13277 38059 13311
rect 38059 13277 38068 13311
rect 38016 13268 38068 13277
rect 38200 13311 38252 13320
rect 38200 13277 38209 13311
rect 38209 13277 38243 13311
rect 38243 13277 38252 13311
rect 38200 13268 38252 13277
rect 40868 13345 40877 13379
rect 40877 13345 40911 13379
rect 40911 13345 40920 13379
rect 44916 13404 44968 13456
rect 40868 13336 40920 13345
rect 45100 13336 45152 13388
rect 41512 13311 41564 13320
rect 41512 13277 41521 13311
rect 41521 13277 41555 13311
rect 41555 13277 41564 13311
rect 41512 13268 41564 13277
rect 41604 13268 41656 13320
rect 36728 13200 36780 13252
rect 37280 13243 37332 13252
rect 37280 13209 37289 13243
rect 37289 13209 37323 13243
rect 37323 13209 37332 13243
rect 41788 13311 41840 13320
rect 41788 13277 41797 13311
rect 41797 13277 41831 13311
rect 41831 13277 41840 13311
rect 42248 13311 42300 13320
rect 41788 13268 41840 13277
rect 42248 13277 42257 13311
rect 42257 13277 42291 13311
rect 42291 13277 42300 13311
rect 42248 13268 42300 13277
rect 42892 13268 42944 13320
rect 43536 13311 43588 13320
rect 43536 13277 43545 13311
rect 43545 13277 43579 13311
rect 43579 13277 43588 13311
rect 43536 13268 43588 13277
rect 43720 13311 43772 13320
rect 43720 13277 43729 13311
rect 43729 13277 43763 13311
rect 43763 13277 43772 13311
rect 43720 13268 43772 13277
rect 44180 13311 44232 13320
rect 44180 13277 44189 13311
rect 44189 13277 44223 13311
rect 44223 13277 44232 13311
rect 44180 13268 44232 13277
rect 47952 13404 48004 13456
rect 47124 13336 47176 13388
rect 48228 13379 48280 13388
rect 48228 13345 48237 13379
rect 48237 13345 48271 13379
rect 48271 13345 48280 13379
rect 48228 13336 48280 13345
rect 45468 13311 45520 13320
rect 37280 13200 37332 13209
rect 45468 13277 45477 13311
rect 45477 13277 45511 13311
rect 45511 13277 45520 13311
rect 45468 13268 45520 13277
rect 45560 13311 45612 13320
rect 45560 13277 45569 13311
rect 45569 13277 45603 13311
rect 45603 13277 45612 13311
rect 45560 13268 45612 13277
rect 45008 13200 45060 13252
rect 22100 13132 22152 13184
rect 22652 13175 22704 13184
rect 22652 13141 22661 13175
rect 22661 13141 22695 13175
rect 22695 13141 22704 13175
rect 22652 13132 22704 13141
rect 33784 13132 33836 13184
rect 37464 13132 37516 13184
rect 40316 13132 40368 13184
rect 43168 13132 43220 13184
rect 43720 13132 43772 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 22836 12928 22888 12980
rect 40132 12928 40184 12980
rect 40776 12928 40828 12980
rect 22192 12835 22244 12844
rect 22192 12801 22201 12835
rect 22201 12801 22235 12835
rect 22235 12801 22244 12835
rect 23204 12860 23256 12912
rect 32312 12860 32364 12912
rect 33048 12860 33100 12912
rect 40316 12903 40368 12912
rect 22468 12835 22520 12844
rect 22192 12792 22244 12801
rect 22468 12801 22477 12835
rect 22477 12801 22511 12835
rect 22511 12801 22520 12835
rect 22468 12792 22520 12801
rect 22744 12792 22796 12844
rect 32496 12835 32548 12844
rect 32496 12801 32505 12835
rect 32505 12801 32539 12835
rect 32539 12801 32548 12835
rect 32496 12792 32548 12801
rect 40316 12869 40325 12903
rect 40325 12869 40359 12903
rect 40359 12869 40368 12903
rect 40316 12860 40368 12869
rect 41696 12928 41748 12980
rect 45008 12971 45060 12980
rect 34152 12835 34204 12844
rect 34152 12801 34186 12835
rect 34186 12801 34204 12835
rect 36360 12835 36412 12844
rect 34152 12792 34204 12801
rect 36360 12801 36369 12835
rect 36369 12801 36403 12835
rect 36403 12801 36412 12835
rect 36360 12792 36412 12801
rect 37464 12835 37516 12844
rect 37464 12801 37473 12835
rect 37473 12801 37507 12835
rect 37507 12801 37516 12835
rect 37464 12792 37516 12801
rect 37648 12835 37700 12844
rect 37648 12801 37657 12835
rect 37657 12801 37691 12835
rect 37691 12801 37700 12835
rect 37648 12792 37700 12801
rect 40224 12835 40276 12844
rect 40224 12801 40233 12835
rect 40233 12801 40267 12835
rect 40267 12801 40276 12835
rect 40224 12792 40276 12801
rect 40408 12835 40460 12844
rect 40408 12801 40417 12835
rect 40417 12801 40451 12835
rect 40451 12801 40460 12835
rect 40408 12792 40460 12801
rect 41144 12835 41196 12844
rect 36452 12767 36504 12776
rect 36452 12733 36461 12767
rect 36461 12733 36495 12767
rect 36495 12733 36504 12767
rect 36728 12767 36780 12776
rect 36452 12724 36504 12733
rect 36728 12733 36737 12767
rect 36737 12733 36771 12767
rect 36771 12733 36780 12767
rect 36728 12724 36780 12733
rect 40776 12724 40828 12776
rect 34520 12588 34572 12640
rect 36820 12588 36872 12640
rect 40408 12588 40460 12640
rect 41144 12801 41153 12835
rect 41153 12801 41187 12835
rect 41187 12801 41196 12835
rect 41144 12792 41196 12801
rect 41236 12835 41288 12844
rect 41236 12801 41246 12835
rect 41246 12801 41280 12835
rect 41280 12801 41288 12835
rect 42248 12860 42300 12912
rect 45008 12937 45017 12971
rect 45017 12937 45051 12971
rect 45051 12937 45060 12971
rect 45008 12928 45060 12937
rect 41236 12792 41288 12801
rect 42892 12835 42944 12844
rect 41328 12656 41380 12708
rect 42892 12801 42901 12835
rect 42901 12801 42935 12835
rect 42935 12801 42944 12835
rect 42892 12792 42944 12801
rect 42984 12792 43036 12844
rect 43168 12835 43220 12844
rect 43168 12801 43177 12835
rect 43177 12801 43211 12835
rect 43211 12801 43220 12835
rect 43168 12792 43220 12801
rect 44180 12792 44232 12844
rect 43260 12656 43312 12708
rect 42708 12588 42760 12640
rect 42800 12588 42852 12640
rect 44364 12724 44416 12776
rect 47308 12792 47360 12844
rect 47492 12792 47544 12844
rect 44732 12588 44784 12640
rect 47124 12631 47176 12640
rect 47124 12597 47133 12631
rect 47133 12597 47167 12631
rect 47167 12597 47176 12631
rect 47124 12588 47176 12597
rect 47952 12631 48004 12640
rect 47952 12597 47961 12631
rect 47961 12597 47995 12631
rect 47995 12597 48004 12631
rect 47952 12588 48004 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 20720 12291 20772 12300
rect 20720 12257 20729 12291
rect 20729 12257 20763 12291
rect 20763 12257 20772 12291
rect 20720 12248 20772 12257
rect 2044 12180 2096 12232
rect 22652 12180 22704 12232
rect 23020 12316 23072 12368
rect 24308 12248 24360 12300
rect 23020 12223 23072 12232
rect 22468 12112 22520 12164
rect 23020 12189 23029 12223
rect 23029 12189 23063 12223
rect 23063 12189 23072 12223
rect 23020 12180 23072 12189
rect 23296 12180 23348 12232
rect 24952 12180 25004 12232
rect 34152 12384 34204 12436
rect 32680 12248 32732 12300
rect 24860 12112 24912 12164
rect 26148 12180 26200 12232
rect 31760 12180 31812 12232
rect 33784 12223 33836 12232
rect 33784 12189 33793 12223
rect 33793 12189 33827 12223
rect 33827 12189 33836 12223
rect 33784 12180 33836 12189
rect 35716 12180 35768 12232
rect 37648 12384 37700 12436
rect 41788 12384 41840 12436
rect 42800 12427 42852 12436
rect 42800 12393 42809 12427
rect 42809 12393 42843 12427
rect 42843 12393 42852 12427
rect 42800 12384 42852 12393
rect 42892 12384 42944 12436
rect 44180 12384 44232 12436
rect 36452 12359 36504 12368
rect 36452 12325 36461 12359
rect 36461 12325 36495 12359
rect 36495 12325 36504 12359
rect 36452 12316 36504 12325
rect 36360 12248 36412 12300
rect 37280 12248 37332 12300
rect 41236 12248 41288 12300
rect 47952 12316 48004 12368
rect 27804 12112 27856 12164
rect 33968 12155 34020 12164
rect 33968 12121 33977 12155
rect 33977 12121 34011 12155
rect 34011 12121 34020 12155
rect 33968 12112 34020 12121
rect 34520 12112 34572 12164
rect 38752 12180 38804 12232
rect 41144 12223 41196 12232
rect 41144 12189 41153 12223
rect 41153 12189 41187 12223
rect 41187 12189 41196 12223
rect 41144 12180 41196 12189
rect 47124 12248 47176 12300
rect 48228 12291 48280 12300
rect 48228 12257 48237 12291
rect 48237 12257 48271 12291
rect 48271 12257 48280 12291
rect 48228 12248 48280 12257
rect 43260 12223 43312 12232
rect 37096 12112 37148 12164
rect 43260 12189 43269 12223
rect 43269 12189 43303 12223
rect 43303 12189 43312 12223
rect 43260 12180 43312 12189
rect 43720 12155 43772 12164
rect 43720 12121 43729 12155
rect 43729 12121 43763 12155
rect 43763 12121 43772 12155
rect 43720 12112 43772 12121
rect 22100 12087 22152 12096
rect 22100 12053 22109 12087
rect 22109 12053 22143 12087
rect 22143 12053 22152 12087
rect 22100 12044 22152 12053
rect 22560 12087 22612 12096
rect 22560 12053 22569 12087
rect 22569 12053 22603 12087
rect 22603 12053 22612 12087
rect 22560 12044 22612 12053
rect 25596 12044 25648 12096
rect 27528 12044 27580 12096
rect 35440 12044 35492 12096
rect 41328 12087 41380 12096
rect 41328 12053 41337 12087
rect 41337 12053 41371 12087
rect 41371 12053 41380 12087
rect 41328 12044 41380 12053
rect 42892 12044 42944 12096
rect 45008 12044 45060 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 22100 11840 22152 11892
rect 22744 11840 22796 11892
rect 2044 11747 2096 11756
rect 2044 11713 2053 11747
rect 2053 11713 2087 11747
rect 2087 11713 2096 11747
rect 2044 11704 2096 11713
rect 22468 11747 22520 11756
rect 22468 11713 22477 11747
rect 22477 11713 22511 11747
rect 22511 11713 22520 11747
rect 22468 11704 22520 11713
rect 23020 11772 23072 11824
rect 22928 11747 22980 11756
rect 22928 11713 22937 11747
rect 22937 11713 22971 11747
rect 22971 11713 22980 11747
rect 22928 11704 22980 11713
rect 24860 11772 24912 11824
rect 25872 11772 25924 11824
rect 2320 11636 2372 11688
rect 2780 11679 2832 11688
rect 2780 11645 2789 11679
rect 2789 11645 2823 11679
rect 2823 11645 2832 11679
rect 2780 11636 2832 11645
rect 25136 11704 25188 11756
rect 25596 11747 25648 11756
rect 25596 11713 25605 11747
rect 25605 11713 25639 11747
rect 25639 11713 25648 11747
rect 25596 11704 25648 11713
rect 27160 11747 27212 11756
rect 27160 11713 27169 11747
rect 27169 11713 27203 11747
rect 27203 11713 27212 11747
rect 27160 11704 27212 11713
rect 27252 11704 27304 11756
rect 27528 11772 27580 11824
rect 27988 11840 28040 11892
rect 30012 11840 30064 11892
rect 31944 11840 31996 11892
rect 33968 11883 34020 11892
rect 33968 11849 33977 11883
rect 33977 11849 34011 11883
rect 34011 11849 34020 11883
rect 33968 11840 34020 11849
rect 37280 11840 37332 11892
rect 27804 11704 27856 11756
rect 28632 11747 28684 11756
rect 28632 11713 28641 11747
rect 28641 11713 28675 11747
rect 28675 11713 28684 11747
rect 28632 11704 28684 11713
rect 28816 11747 28868 11756
rect 28816 11713 28825 11747
rect 28825 11713 28859 11747
rect 28859 11713 28868 11747
rect 28816 11704 28868 11713
rect 29000 11747 29052 11756
rect 29000 11713 29009 11747
rect 29009 11713 29043 11747
rect 29043 11713 29052 11747
rect 29000 11704 29052 11713
rect 29092 11747 29144 11756
rect 29092 11713 29101 11747
rect 29101 11713 29135 11747
rect 29135 11713 29144 11747
rect 29092 11704 29144 11713
rect 29736 11747 29788 11756
rect 29736 11713 29745 11747
rect 29745 11713 29779 11747
rect 29779 11713 29788 11747
rect 29736 11704 29788 11713
rect 29920 11704 29972 11756
rect 30656 11747 30708 11756
rect 30656 11713 30665 11747
rect 30665 11713 30699 11747
rect 30699 11713 30708 11747
rect 30656 11704 30708 11713
rect 24860 11636 24912 11688
rect 33600 11772 33652 11824
rect 32036 11704 32088 11756
rect 33784 11747 33836 11756
rect 33784 11713 33793 11747
rect 33793 11713 33827 11747
rect 33827 11713 33836 11747
rect 33784 11704 33836 11713
rect 36360 11772 36412 11824
rect 41144 11840 41196 11892
rect 35900 11704 35952 11756
rect 25044 11568 25096 11620
rect 31852 11636 31904 11688
rect 25964 11568 26016 11620
rect 32404 11568 32456 11620
rect 36728 11636 36780 11688
rect 38016 11704 38068 11756
rect 38384 11747 38436 11756
rect 38384 11713 38393 11747
rect 38393 11713 38427 11747
rect 38427 11713 38436 11747
rect 38384 11704 38436 11713
rect 43076 11704 43128 11756
rect 43628 11747 43680 11756
rect 38936 11636 38988 11688
rect 42800 11679 42852 11688
rect 42800 11645 42809 11679
rect 42809 11645 42843 11679
rect 42843 11645 42852 11679
rect 42800 11636 42852 11645
rect 43260 11636 43312 11688
rect 43628 11713 43637 11747
rect 43637 11713 43671 11747
rect 43671 11713 43680 11747
rect 43628 11704 43680 11713
rect 44732 11772 44784 11824
rect 44456 11704 44508 11756
rect 44916 11704 44968 11756
rect 22652 11500 22704 11552
rect 24768 11500 24820 11552
rect 25412 11543 25464 11552
rect 25412 11509 25421 11543
rect 25421 11509 25455 11543
rect 25455 11509 25464 11543
rect 25412 11500 25464 11509
rect 25780 11543 25832 11552
rect 25780 11509 25789 11543
rect 25789 11509 25823 11543
rect 25823 11509 25832 11543
rect 25780 11500 25832 11509
rect 25872 11500 25924 11552
rect 27712 11500 27764 11552
rect 32128 11500 32180 11552
rect 32312 11543 32364 11552
rect 32312 11509 32321 11543
rect 32321 11509 32355 11543
rect 32355 11509 32364 11543
rect 32312 11500 32364 11509
rect 32588 11500 32640 11552
rect 36452 11500 36504 11552
rect 37832 11543 37884 11552
rect 37832 11509 37841 11543
rect 37841 11509 37875 11543
rect 37875 11509 37884 11543
rect 37832 11500 37884 11509
rect 38292 11500 38344 11552
rect 38568 11543 38620 11552
rect 38568 11509 38577 11543
rect 38577 11509 38611 11543
rect 38611 11509 38620 11543
rect 44732 11611 44784 11620
rect 44732 11577 44741 11611
rect 44741 11577 44775 11611
rect 44775 11577 44784 11611
rect 44732 11568 44784 11577
rect 38568 11500 38620 11509
rect 44180 11500 44232 11552
rect 45100 11500 45152 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 2320 11339 2372 11348
rect 2320 11305 2329 11339
rect 2329 11305 2363 11339
rect 2363 11305 2372 11339
rect 2320 11296 2372 11305
rect 23296 11296 23348 11348
rect 25964 11228 26016 11280
rect 20720 11160 20772 11212
rect 21824 11160 21876 11212
rect 2228 11135 2280 11144
rect 2228 11101 2237 11135
rect 2237 11101 2271 11135
rect 2271 11101 2280 11135
rect 2228 11092 2280 11101
rect 3056 11135 3108 11144
rect 3056 11101 3065 11135
rect 3065 11101 3099 11135
rect 3099 11101 3108 11135
rect 3056 11092 3108 11101
rect 3792 11092 3844 11144
rect 12624 11092 12676 11144
rect 26148 11092 26200 11144
rect 27528 11135 27580 11144
rect 27528 11101 27537 11135
rect 27537 11101 27571 11135
rect 27571 11101 27580 11135
rect 27528 11092 27580 11101
rect 29000 11296 29052 11348
rect 31668 11296 31720 11348
rect 36360 11296 36412 11348
rect 32128 11228 32180 11280
rect 22468 11024 22520 11076
rect 25412 11024 25464 11076
rect 2872 10956 2924 11008
rect 12532 10956 12584 11008
rect 23296 10999 23348 11008
rect 23296 10965 23305 10999
rect 23305 10965 23339 10999
rect 23339 10965 23348 10999
rect 23296 10956 23348 10965
rect 28724 11160 28776 11212
rect 29184 11135 29236 11144
rect 29184 11101 29193 11135
rect 29193 11101 29227 11135
rect 29227 11101 29236 11135
rect 29736 11135 29788 11144
rect 29184 11092 29236 11101
rect 29736 11101 29745 11135
rect 29745 11101 29779 11135
rect 29779 11101 29788 11135
rect 29736 11092 29788 11101
rect 30012 11135 30064 11144
rect 30012 11101 30021 11135
rect 30021 11101 30055 11135
rect 30055 11101 30064 11135
rect 30012 11092 30064 11101
rect 31760 11092 31812 11144
rect 32864 11092 32916 11144
rect 34520 11160 34572 11212
rect 29920 11067 29972 11076
rect 29920 11033 29929 11067
rect 29929 11033 29963 11067
rect 29963 11033 29972 11067
rect 29920 11024 29972 11033
rect 32312 11024 32364 11076
rect 32404 11024 32456 11076
rect 35808 11228 35860 11280
rect 39120 11296 39172 11348
rect 43076 11339 43128 11348
rect 43076 11305 43085 11339
rect 43085 11305 43119 11339
rect 43119 11305 43128 11339
rect 43076 11296 43128 11305
rect 44456 11296 44508 11348
rect 35440 11203 35492 11212
rect 35440 11169 35449 11203
rect 35449 11169 35483 11203
rect 35483 11169 35492 11203
rect 35440 11160 35492 11169
rect 35900 11092 35952 11144
rect 41328 11228 41380 11280
rect 38108 11160 38160 11212
rect 40316 11160 40368 11212
rect 40868 11160 40920 11212
rect 43904 11160 43956 11212
rect 45652 11160 45704 11212
rect 37924 11092 37976 11144
rect 38016 11135 38068 11144
rect 38016 11101 38025 11135
rect 38025 11101 38059 11135
rect 38059 11101 38068 11135
rect 38476 11135 38528 11144
rect 38016 11092 38068 11101
rect 38476 11101 38485 11135
rect 38485 11101 38519 11135
rect 38519 11101 38528 11135
rect 38476 11092 38528 11101
rect 39120 11135 39172 11144
rect 39120 11101 39129 11135
rect 39129 11101 39163 11135
rect 39163 11101 39172 11135
rect 39120 11092 39172 11101
rect 42984 11092 43036 11144
rect 44456 11135 44508 11144
rect 44456 11101 44465 11135
rect 44465 11101 44499 11135
rect 44499 11101 44508 11135
rect 44456 11092 44508 11101
rect 45100 11092 45152 11144
rect 45560 11135 45612 11144
rect 45560 11101 45569 11135
rect 45569 11101 45603 11135
rect 45603 11101 45612 11135
rect 45560 11092 45612 11101
rect 30564 10956 30616 11008
rect 32772 10956 32824 11008
rect 33140 10956 33192 11008
rect 34060 10956 34112 11008
rect 35532 10956 35584 11008
rect 38660 10956 38712 11008
rect 42800 10956 42852 11008
rect 44180 11024 44232 11076
rect 44916 10956 44968 11008
rect 45744 10999 45796 11008
rect 45744 10965 45753 10999
rect 45753 10965 45787 10999
rect 45787 10965 45796 10999
rect 45744 10956 45796 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 22468 10795 22520 10804
rect 22468 10761 22477 10795
rect 22477 10761 22511 10795
rect 22511 10761 22520 10795
rect 22468 10752 22520 10761
rect 2872 10727 2924 10736
rect 2872 10693 2881 10727
rect 2881 10693 2915 10727
rect 2915 10693 2924 10727
rect 2872 10684 2924 10693
rect 12532 10727 12584 10736
rect 12532 10693 12541 10727
rect 12541 10693 12575 10727
rect 12575 10693 12584 10727
rect 12532 10684 12584 10693
rect 25044 10684 25096 10736
rect 30656 10752 30708 10804
rect 30932 10752 30984 10804
rect 35808 10752 35860 10804
rect 22652 10659 22704 10668
rect 22652 10625 22661 10659
rect 22661 10625 22695 10659
rect 22695 10625 22704 10659
rect 22652 10616 22704 10625
rect 3056 10548 3108 10600
rect 3148 10591 3200 10600
rect 3148 10557 3157 10591
rect 3157 10557 3191 10591
rect 3191 10557 3200 10591
rect 3148 10548 3200 10557
rect 12624 10548 12676 10600
rect 14188 10591 14240 10600
rect 14188 10557 14197 10591
rect 14197 10557 14231 10591
rect 14231 10557 14240 10591
rect 14188 10548 14240 10557
rect 21824 10548 21876 10600
rect 24584 10616 24636 10668
rect 26516 10616 26568 10668
rect 27528 10659 27580 10668
rect 23296 10548 23348 10600
rect 27528 10625 27537 10659
rect 27537 10625 27571 10659
rect 27571 10625 27580 10659
rect 27528 10616 27580 10625
rect 27712 10659 27764 10668
rect 27712 10625 27721 10659
rect 27721 10625 27755 10659
rect 27755 10625 27764 10659
rect 27712 10616 27764 10625
rect 29000 10616 29052 10668
rect 29184 10616 29236 10668
rect 30564 10616 30616 10668
rect 31484 10684 31536 10736
rect 30932 10659 30984 10668
rect 30932 10625 30941 10659
rect 30941 10625 30975 10659
rect 30975 10625 30984 10659
rect 34060 10684 34112 10736
rect 35532 10727 35584 10736
rect 35532 10693 35541 10727
rect 35541 10693 35575 10727
rect 35575 10693 35584 10727
rect 35532 10684 35584 10693
rect 30932 10616 30984 10625
rect 32772 10616 32824 10668
rect 33140 10616 33192 10668
rect 35624 10659 35676 10668
rect 28816 10548 28868 10600
rect 29736 10591 29788 10600
rect 29736 10557 29745 10591
rect 29745 10557 29779 10591
rect 29779 10557 29788 10591
rect 29736 10548 29788 10557
rect 29920 10548 29972 10600
rect 28908 10480 28960 10532
rect 31944 10480 31996 10532
rect 35624 10625 35633 10659
rect 35633 10625 35667 10659
rect 35667 10625 35676 10659
rect 35624 10616 35676 10625
rect 35716 10659 35768 10668
rect 35716 10625 35725 10659
rect 35725 10625 35759 10659
rect 35759 10625 35768 10659
rect 38568 10752 38620 10804
rect 38660 10795 38712 10804
rect 38660 10761 38669 10795
rect 38669 10761 38703 10795
rect 38703 10761 38712 10795
rect 38660 10752 38712 10761
rect 37832 10684 37884 10736
rect 38384 10684 38436 10736
rect 35716 10616 35768 10625
rect 38936 10659 38988 10668
rect 36728 10548 36780 10600
rect 38936 10625 38945 10659
rect 38945 10625 38979 10659
rect 38979 10625 38988 10659
rect 38936 10616 38988 10625
rect 40132 10752 40184 10804
rect 41052 10752 41104 10804
rect 41604 10752 41656 10804
rect 44916 10752 44968 10804
rect 38476 10548 38528 10600
rect 39212 10548 39264 10600
rect 44640 10684 44692 10736
rect 40316 10659 40368 10668
rect 40316 10625 40325 10659
rect 40325 10625 40359 10659
rect 40359 10625 40368 10659
rect 40316 10616 40368 10625
rect 38200 10480 38252 10532
rect 40868 10616 40920 10668
rect 44180 10659 44232 10668
rect 41052 10480 41104 10532
rect 44180 10625 44189 10659
rect 44189 10625 44223 10659
rect 44223 10625 44232 10659
rect 44180 10616 44232 10625
rect 44548 10616 44600 10668
rect 44916 10659 44968 10668
rect 44916 10625 44925 10659
rect 44925 10625 44959 10659
rect 44959 10625 44968 10659
rect 44916 10616 44968 10625
rect 45376 10684 45428 10736
rect 45744 10684 45796 10736
rect 45192 10616 45244 10668
rect 44088 10591 44140 10600
rect 44088 10557 44097 10591
rect 44097 10557 44131 10591
rect 44131 10557 44140 10591
rect 44088 10548 44140 10557
rect 44456 10548 44508 10600
rect 44824 10548 44876 10600
rect 42616 10480 42668 10532
rect 22744 10412 22796 10464
rect 27896 10455 27948 10464
rect 27896 10421 27905 10455
rect 27905 10421 27939 10455
rect 27939 10421 27948 10455
rect 27896 10412 27948 10421
rect 29000 10455 29052 10464
rect 29000 10421 29009 10455
rect 29009 10421 29043 10455
rect 29043 10421 29052 10455
rect 29000 10412 29052 10421
rect 29828 10455 29880 10464
rect 29828 10421 29837 10455
rect 29837 10421 29871 10455
rect 29871 10421 29880 10455
rect 29828 10412 29880 10421
rect 32128 10412 32180 10464
rect 35900 10455 35952 10464
rect 35900 10421 35909 10455
rect 35909 10421 35943 10455
rect 35943 10421 35952 10455
rect 35900 10412 35952 10421
rect 36912 10455 36964 10464
rect 36912 10421 36921 10455
rect 36921 10421 36955 10455
rect 36955 10421 36964 10455
rect 36912 10412 36964 10421
rect 38292 10412 38344 10464
rect 40408 10412 40460 10464
rect 41144 10455 41196 10464
rect 41144 10421 41153 10455
rect 41153 10421 41187 10455
rect 41187 10421 41196 10455
rect 41144 10412 41196 10421
rect 43536 10412 43588 10464
rect 44824 10412 44876 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 24584 10251 24636 10260
rect 24584 10217 24593 10251
rect 24593 10217 24627 10251
rect 24627 10217 24636 10251
rect 24584 10208 24636 10217
rect 27712 10208 27764 10260
rect 29092 10208 29144 10260
rect 29920 10208 29972 10260
rect 32588 10208 32640 10260
rect 33784 10208 33836 10260
rect 35624 10208 35676 10260
rect 38292 10208 38344 10260
rect 40868 10208 40920 10260
rect 45652 10208 45704 10260
rect 22836 10140 22888 10192
rect 25780 10140 25832 10192
rect 21824 10115 21876 10124
rect 21824 10081 21833 10115
rect 21833 10081 21867 10115
rect 21867 10081 21876 10115
rect 21824 10072 21876 10081
rect 25044 10115 25096 10124
rect 25044 10081 25053 10115
rect 25053 10081 25087 10115
rect 25087 10081 25096 10115
rect 25044 10072 25096 10081
rect 26148 10115 26200 10124
rect 26148 10081 26157 10115
rect 26157 10081 26191 10115
rect 26191 10081 26200 10115
rect 26148 10072 26200 10081
rect 30840 10183 30892 10192
rect 30840 10149 30849 10183
rect 30849 10149 30883 10183
rect 30883 10149 30892 10183
rect 30840 10140 30892 10149
rect 2044 10004 2096 10056
rect 24768 10047 24820 10056
rect 24768 10013 24777 10047
rect 24777 10013 24811 10047
rect 24811 10013 24820 10047
rect 24768 10004 24820 10013
rect 27896 10004 27948 10056
rect 29736 10072 29788 10124
rect 32036 10140 32088 10192
rect 32864 10140 32916 10192
rect 34060 10183 34112 10192
rect 28172 10047 28224 10056
rect 28172 10013 28181 10047
rect 28181 10013 28215 10047
rect 28215 10013 28224 10047
rect 28172 10004 28224 10013
rect 30196 10047 30248 10056
rect 30196 10013 30205 10047
rect 30205 10013 30239 10047
rect 30239 10013 30248 10047
rect 30196 10004 30248 10013
rect 34060 10149 34069 10183
rect 34069 10149 34103 10183
rect 34103 10149 34112 10183
rect 34060 10140 34112 10149
rect 41604 10183 41656 10192
rect 41604 10149 41613 10183
rect 41613 10149 41647 10183
rect 41647 10149 41656 10183
rect 41604 10140 41656 10149
rect 36912 10072 36964 10124
rect 31944 10047 31996 10056
rect 22376 9936 22428 9988
rect 28724 9936 28776 9988
rect 23204 9911 23256 9920
rect 23204 9877 23213 9911
rect 23213 9877 23247 9911
rect 23247 9877 23256 9911
rect 23204 9868 23256 9877
rect 29184 9936 29236 9988
rect 30840 9936 30892 9988
rect 31392 9936 31444 9988
rect 31944 10013 31953 10047
rect 31953 10013 31987 10047
rect 31987 10013 31996 10047
rect 31944 10004 31996 10013
rect 32404 9868 32456 9920
rect 33140 10004 33192 10056
rect 35900 10004 35952 10056
rect 38200 10047 38252 10056
rect 38200 10013 38209 10047
rect 38209 10013 38243 10047
rect 38243 10013 38252 10047
rect 38200 10004 38252 10013
rect 38568 10004 38620 10056
rect 38752 10004 38804 10056
rect 39212 9936 39264 9988
rect 38016 9911 38068 9920
rect 38016 9877 38025 9911
rect 38025 9877 38059 9911
rect 38059 9877 38068 9911
rect 38016 9868 38068 9877
rect 39396 9868 39448 9920
rect 40224 10047 40276 10056
rect 40224 10013 40233 10047
rect 40233 10013 40267 10047
rect 40267 10013 40276 10047
rect 42616 10072 42668 10124
rect 43904 10115 43956 10124
rect 43904 10081 43913 10115
rect 43913 10081 43947 10115
rect 43947 10081 43956 10115
rect 43904 10072 43956 10081
rect 44180 10072 44232 10124
rect 42064 10047 42116 10056
rect 40224 10004 40276 10013
rect 42064 10013 42073 10047
rect 42073 10013 42107 10047
rect 42107 10013 42116 10047
rect 42064 10004 42116 10013
rect 43536 10047 43588 10056
rect 43536 10013 43545 10047
rect 43545 10013 43579 10047
rect 43579 10013 43588 10047
rect 43812 10047 43864 10056
rect 43536 10004 43588 10013
rect 43812 10013 43821 10047
rect 43821 10013 43855 10047
rect 43855 10013 43864 10047
rect 43812 10004 43864 10013
rect 44088 10004 44140 10056
rect 44916 10004 44968 10056
rect 40316 9936 40368 9988
rect 45376 9979 45428 9988
rect 45376 9945 45385 9979
rect 45385 9945 45419 9979
rect 45419 9945 45428 9979
rect 45376 9936 45428 9945
rect 40592 9868 40644 9920
rect 43260 9911 43312 9920
rect 43260 9877 43269 9911
rect 43269 9877 43303 9911
rect 43303 9877 43312 9911
rect 43260 9868 43312 9877
rect 44824 9868 44876 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 22376 9707 22428 9716
rect 22376 9673 22385 9707
rect 22385 9673 22419 9707
rect 22419 9673 22428 9707
rect 22376 9664 22428 9673
rect 23204 9664 23256 9716
rect 2044 9571 2096 9580
rect 2044 9537 2053 9571
rect 2053 9537 2087 9571
rect 2087 9537 2096 9571
rect 2044 9528 2096 9537
rect 22560 9571 22612 9580
rect 22560 9537 22569 9571
rect 22569 9537 22603 9571
rect 22603 9537 22612 9571
rect 22560 9528 22612 9537
rect 22744 9571 22796 9580
rect 22744 9537 22753 9571
rect 22753 9537 22787 9571
rect 22787 9537 22796 9571
rect 22744 9528 22796 9537
rect 23204 9528 23256 9580
rect 27712 9528 27764 9580
rect 28172 9664 28224 9716
rect 29828 9664 29880 9716
rect 32772 9664 32824 9716
rect 35716 9664 35768 9716
rect 38568 9664 38620 9716
rect 40684 9664 40736 9716
rect 2320 9460 2372 9512
rect 2780 9503 2832 9512
rect 2780 9469 2789 9503
rect 2789 9469 2823 9503
rect 2823 9469 2832 9503
rect 2780 9460 2832 9469
rect 29092 9596 29144 9648
rect 29000 9528 29052 9580
rect 30196 9596 30248 9648
rect 32036 9528 32088 9580
rect 32404 9571 32456 9580
rect 32404 9537 32413 9571
rect 32413 9537 32447 9571
rect 32447 9537 32456 9571
rect 32404 9528 32456 9537
rect 40224 9596 40276 9648
rect 41144 9596 41196 9648
rect 29828 9460 29880 9512
rect 35992 9503 36044 9512
rect 31852 9392 31904 9444
rect 35624 9392 35676 9444
rect 35992 9469 36001 9503
rect 36001 9469 36035 9503
rect 36035 9469 36044 9503
rect 35992 9460 36044 9469
rect 28908 9324 28960 9376
rect 29736 9367 29788 9376
rect 29736 9333 29745 9367
rect 29745 9333 29779 9367
rect 29779 9333 29788 9367
rect 29736 9324 29788 9333
rect 31392 9367 31444 9376
rect 31392 9333 31401 9367
rect 31401 9333 31435 9367
rect 31435 9333 31444 9367
rect 31392 9324 31444 9333
rect 32036 9324 32088 9376
rect 38016 9528 38068 9580
rect 39396 9528 39448 9580
rect 39488 9571 39540 9580
rect 39488 9537 39497 9571
rect 39497 9537 39531 9571
rect 39531 9537 39540 9571
rect 39488 9528 39540 9537
rect 40132 9528 40184 9580
rect 40408 9571 40460 9580
rect 40408 9537 40417 9571
rect 40417 9537 40451 9571
rect 40451 9537 40460 9571
rect 40408 9528 40460 9537
rect 40592 9571 40644 9580
rect 40592 9537 40601 9571
rect 40601 9537 40635 9571
rect 40635 9537 40644 9571
rect 40592 9528 40644 9537
rect 40684 9571 40736 9580
rect 40684 9537 40719 9571
rect 40719 9537 40736 9571
rect 40684 9528 40736 9537
rect 41604 9596 41656 9648
rect 43812 9664 43864 9716
rect 43904 9664 43956 9716
rect 43260 9596 43312 9648
rect 45652 9596 45704 9648
rect 40316 9460 40368 9512
rect 42616 9571 42668 9580
rect 38476 9392 38528 9444
rect 41328 9392 41380 9444
rect 42616 9537 42625 9571
rect 42625 9537 42659 9571
rect 42659 9537 42668 9571
rect 42616 9528 42668 9537
rect 44088 9528 44140 9580
rect 42064 9460 42116 9512
rect 45008 9435 45060 9444
rect 45008 9401 45017 9435
rect 45017 9401 45051 9435
rect 45051 9401 45060 9435
rect 45008 9392 45060 9401
rect 38752 9324 38804 9376
rect 39212 9324 39264 9376
rect 44824 9367 44876 9376
rect 44824 9333 44833 9367
rect 44833 9333 44867 9367
rect 44867 9333 44876 9367
rect 44824 9324 44876 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 2320 9163 2372 9172
rect 2320 9129 2329 9163
rect 2329 9129 2363 9163
rect 2363 9129 2372 9163
rect 2320 9120 2372 9129
rect 32036 9163 32088 9172
rect 32036 9129 32045 9163
rect 32045 9129 32079 9163
rect 32079 9129 32088 9163
rect 32036 9120 32088 9129
rect 39488 9120 39540 9172
rect 39672 9120 39724 9172
rect 44088 9095 44140 9104
rect 44088 9061 44097 9095
rect 44097 9061 44131 9095
rect 44131 9061 44140 9095
rect 44088 9052 44140 9061
rect 38752 8984 38804 9036
rect 2228 8959 2280 8968
rect 2228 8925 2237 8959
rect 2237 8925 2271 8959
rect 2271 8925 2280 8959
rect 2228 8916 2280 8925
rect 8300 8916 8352 8968
rect 31944 8959 31996 8968
rect 31944 8925 31953 8959
rect 31953 8925 31987 8959
rect 31987 8925 31996 8959
rect 31944 8916 31996 8925
rect 32128 8959 32180 8968
rect 32128 8925 32137 8959
rect 32137 8925 32171 8959
rect 32171 8925 32180 8959
rect 32128 8916 32180 8925
rect 39212 8959 39264 8968
rect 39212 8925 39221 8959
rect 39221 8925 39255 8959
rect 39255 8925 39264 8959
rect 39212 8916 39264 8925
rect 43904 8984 43956 9036
rect 41328 8916 41380 8968
rect 45376 8916 45428 8968
rect 47952 8891 48004 8900
rect 47952 8857 47961 8891
rect 47961 8857 47995 8891
rect 47995 8857 48004 8891
rect 47952 8848 48004 8857
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 47860 8483 47912 8492
rect 47860 8449 47869 8483
rect 47869 8449 47903 8483
rect 47903 8449 47912 8483
rect 47860 8440 47912 8449
rect 32220 8372 32272 8424
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 2044 7828 2096 7880
rect 3240 7828 3292 7880
rect 5632 7828 5684 7880
rect 2228 7692 2280 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 2228 7463 2280 7472
rect 2228 7429 2237 7463
rect 2237 7429 2271 7463
rect 2271 7429 2280 7463
rect 2228 7420 2280 7429
rect 2044 7395 2096 7404
rect 2044 7361 2053 7395
rect 2053 7361 2087 7395
rect 2087 7361 2096 7395
rect 2044 7352 2096 7361
rect 2780 7327 2832 7336
rect 2780 7293 2789 7327
rect 2789 7293 2823 7327
rect 2823 7293 2832 7327
rect 2780 7284 2832 7293
rect 47952 7191 48004 7200
rect 47952 7157 47961 7191
rect 47961 7157 47995 7191
rect 47995 7157 48004 7191
rect 47952 7148 48004 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 2780 6851 2832 6860
rect 2780 6817 2789 6851
rect 2789 6817 2823 6851
rect 2823 6817 2832 6851
rect 2780 6808 2832 6817
rect 47952 6808 48004 6860
rect 48228 6851 48280 6860
rect 48228 6817 48237 6851
rect 48237 6817 48271 6851
rect 48271 6817 48280 6851
rect 48228 6808 48280 6817
rect 1584 6783 1636 6792
rect 1584 6749 1593 6783
rect 1593 6749 1627 6783
rect 1627 6749 1636 6783
rect 1584 6740 1636 6749
rect 1768 6715 1820 6724
rect 1768 6681 1777 6715
rect 1777 6681 1811 6715
rect 1811 6681 1820 6715
rect 1768 6672 1820 6681
rect 47860 6672 47912 6724
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 1768 6400 1820 6452
rect 47860 6443 47912 6452
rect 47860 6409 47869 6443
rect 47869 6409 47903 6443
rect 47903 6409 47912 6443
rect 47860 6400 47912 6409
rect 1584 6264 1636 6316
rect 2872 6264 2924 6316
rect 47032 6264 47084 6316
rect 47768 6307 47820 6316
rect 47768 6273 47777 6307
rect 47777 6273 47811 6307
rect 47811 6273 47820 6307
rect 47768 6264 47820 6273
rect 39212 6060 39264 6112
rect 43076 6060 43128 6112
rect 46480 6103 46532 6112
rect 46480 6069 46489 6103
rect 46489 6069 46523 6103
rect 46523 6069 46532 6103
rect 46480 6060 46532 6069
rect 47216 6103 47268 6112
rect 47216 6069 47225 6103
rect 47225 6069 47259 6103
rect 47259 6069 47268 6103
rect 47216 6060 47268 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 47216 5720 47268 5772
rect 48228 5763 48280 5772
rect 48228 5729 48237 5763
rect 48237 5729 48271 5763
rect 48271 5729 48280 5763
rect 48228 5720 48280 5729
rect 1860 5695 1912 5704
rect 1860 5661 1869 5695
rect 1869 5661 1903 5695
rect 1903 5661 1912 5695
rect 1860 5652 1912 5661
rect 2688 5652 2740 5704
rect 3148 5695 3200 5704
rect 3148 5661 3157 5695
rect 3157 5661 3191 5695
rect 3191 5661 3200 5695
rect 3148 5652 3200 5661
rect 9772 5695 9824 5704
rect 9772 5661 9781 5695
rect 9781 5661 9815 5695
rect 9815 5661 9824 5695
rect 9772 5652 9824 5661
rect 16120 5652 16172 5704
rect 39028 5652 39080 5704
rect 46020 5695 46072 5704
rect 46020 5661 46029 5695
rect 46029 5661 46063 5695
rect 46063 5661 46072 5695
rect 46020 5652 46072 5661
rect 47584 5584 47636 5636
rect 1768 5516 1820 5568
rect 10048 5516 10100 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 39212 5287 39264 5296
rect 39212 5253 39221 5287
rect 39221 5253 39255 5287
rect 39255 5253 39264 5287
rect 39212 5244 39264 5253
rect 39028 5219 39080 5228
rect 39028 5185 39037 5219
rect 39037 5185 39071 5219
rect 39071 5185 39080 5219
rect 39028 5176 39080 5185
rect 47492 5312 47544 5364
rect 47768 5219 47820 5228
rect 47768 5185 47777 5219
rect 47777 5185 47811 5219
rect 47811 5185 47820 5219
rect 47768 5176 47820 5185
rect 2872 5108 2924 5160
rect 2964 5151 3016 5160
rect 2964 5117 2973 5151
rect 2973 5117 3007 5151
rect 3007 5117 3016 5151
rect 40040 5151 40092 5160
rect 2964 5108 3016 5117
rect 40040 5117 40049 5151
rect 40049 5117 40083 5151
rect 40083 5117 40092 5151
rect 40040 5108 40092 5117
rect 46020 5108 46072 5160
rect 47216 5151 47268 5160
rect 47216 5117 47225 5151
rect 47225 5117 47259 5151
rect 47259 5117 47268 5151
rect 47216 5108 47268 5117
rect 44272 5015 44324 5024
rect 44272 4981 44281 5015
rect 44281 4981 44315 5015
rect 44315 4981 44324 5015
rect 44272 4972 44324 4981
rect 45376 4972 45428 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 47584 4811 47636 4820
rect 47584 4777 47593 4811
rect 47593 4777 47627 4811
rect 47627 4777 47636 4811
rect 47584 4768 47636 4777
rect 3148 4700 3200 4752
rect 1768 4675 1820 4684
rect 1768 4641 1777 4675
rect 1777 4641 1811 4675
rect 1811 4641 1820 4675
rect 1768 4632 1820 4641
rect 2780 4675 2832 4684
rect 2780 4641 2789 4675
rect 2789 4641 2823 4675
rect 2823 4641 2832 4675
rect 2780 4632 2832 4641
rect 3516 4632 3568 4684
rect 9772 4632 9824 4684
rect 10048 4675 10100 4684
rect 10048 4641 10057 4675
rect 10057 4641 10091 4675
rect 10091 4641 10100 4675
rect 10048 4632 10100 4641
rect 4620 4564 4672 4616
rect 4988 4607 5040 4616
rect 4988 4573 4997 4607
rect 4997 4573 5031 4607
rect 5031 4573 5040 4607
rect 4988 4564 5040 4573
rect 5540 4607 5592 4616
rect 5540 4573 5549 4607
rect 5549 4573 5583 4607
rect 5583 4573 5592 4607
rect 5540 4564 5592 4573
rect 47676 4700 47728 4752
rect 44272 4632 44324 4684
rect 45376 4675 45428 4684
rect 45376 4641 45385 4675
rect 45385 4641 45419 4675
rect 45419 4641 45428 4675
rect 45376 4632 45428 4641
rect 45652 4675 45704 4684
rect 45652 4641 45661 4675
rect 45661 4641 45695 4675
rect 45695 4641 45704 4675
rect 45652 4632 45704 4641
rect 44640 4607 44692 4616
rect 44640 4573 44649 4607
rect 44649 4573 44683 4607
rect 44683 4573 44692 4607
rect 44640 4564 44692 4573
rect 47492 4607 47544 4616
rect 47492 4573 47501 4607
rect 47501 4573 47535 4607
rect 47535 4573 47544 4607
rect 47492 4564 47544 4573
rect 48136 4607 48188 4616
rect 48136 4573 48145 4607
rect 48145 4573 48179 4607
rect 48179 4573 48188 4607
rect 48136 4564 48188 4573
rect 6276 4539 6328 4548
rect 6276 4505 6285 4539
rect 6285 4505 6319 4539
rect 6319 4505 6328 4539
rect 6276 4496 6328 4505
rect 39948 4428 40000 4480
rect 43260 4428 43312 4480
rect 46940 4428 46992 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 43260 4199 43312 4208
rect 2872 4131 2924 4140
rect 2872 4097 2881 4131
rect 2881 4097 2915 4131
rect 2915 4097 2924 4131
rect 2872 4088 2924 4097
rect 2964 4020 3016 4072
rect 3976 4063 4028 4072
rect 3976 4029 3985 4063
rect 3985 4029 4019 4063
rect 4019 4029 4028 4063
rect 3976 4020 4028 4029
rect 43260 4165 43269 4199
rect 43269 4165 43303 4199
rect 43303 4165 43312 4199
rect 43260 4156 43312 4165
rect 48136 4224 48188 4276
rect 5540 4088 5592 4140
rect 2044 3884 2096 3936
rect 3240 3952 3292 4004
rect 6552 4020 6604 4072
rect 9864 4088 9916 4140
rect 13268 4020 13320 4072
rect 19432 4088 19484 4140
rect 39948 4131 40000 4140
rect 39948 4097 39957 4131
rect 39957 4097 39991 4131
rect 39991 4097 40000 4131
rect 39948 4088 40000 4097
rect 43076 4131 43128 4140
rect 17132 4020 17184 4072
rect 19708 4020 19760 4072
rect 22192 4063 22244 4072
rect 10140 3952 10192 4004
rect 22192 4029 22201 4063
rect 22201 4029 22235 4063
rect 22235 4029 22244 4063
rect 22192 4020 22244 4029
rect 22560 4063 22612 4072
rect 22560 4029 22569 4063
rect 22569 4029 22603 4063
rect 22603 4029 22612 4063
rect 22560 4020 22612 4029
rect 43076 4097 43085 4131
rect 43085 4097 43119 4131
rect 43119 4097 43128 4131
rect 43076 4088 43128 4097
rect 41604 4020 41656 4072
rect 44916 4063 44968 4072
rect 44916 4029 44925 4063
rect 44925 4029 44959 4063
rect 44959 4029 44968 4063
rect 44916 4020 44968 4029
rect 47400 4088 47452 4140
rect 46940 4020 46992 4072
rect 47676 4020 47728 4072
rect 47952 3952 48004 4004
rect 5632 3884 5684 3936
rect 6276 3884 6328 3936
rect 6736 3927 6788 3936
rect 6736 3893 6745 3927
rect 6745 3893 6779 3927
rect 6779 3893 6788 3927
rect 6736 3884 6788 3893
rect 7288 3884 7340 3936
rect 10692 3884 10744 3936
rect 12992 3884 13044 3936
rect 16764 3884 16816 3936
rect 17316 3884 17368 3936
rect 19892 3884 19944 3936
rect 20168 3927 20220 3936
rect 20168 3893 20177 3927
rect 20177 3893 20211 3927
rect 20211 3893 20220 3927
rect 20168 3884 20220 3893
rect 24768 3884 24820 3936
rect 25964 3884 26016 3936
rect 27160 3884 27212 3936
rect 40132 3884 40184 3936
rect 40776 3884 40828 3936
rect 41420 3884 41472 3936
rect 46112 3884 46164 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 2964 3680 3016 3732
rect 3976 3680 4028 3732
rect 9588 3680 9640 3732
rect 12900 3680 12952 3732
rect 14188 3680 14240 3732
rect 1952 3519 2004 3528
rect 1952 3485 1961 3519
rect 1961 3485 1995 3519
rect 1995 3485 2004 3519
rect 1952 3476 2004 3485
rect 5172 3612 5224 3664
rect 9864 3612 9916 3664
rect 5448 3544 5500 3596
rect 6460 3587 6512 3596
rect 6460 3553 6469 3587
rect 6469 3553 6503 3587
rect 6503 3553 6512 3587
rect 6460 3544 6512 3553
rect 6552 3544 6604 3596
rect 10692 3587 10744 3596
rect 10692 3553 10701 3587
rect 10701 3553 10735 3587
rect 10735 3553 10744 3587
rect 10692 3544 10744 3553
rect 10968 3587 11020 3596
rect 10968 3553 10977 3587
rect 10977 3553 11011 3587
rect 11011 3553 11020 3587
rect 10968 3544 11020 3553
rect 4160 3476 4212 3528
rect 8300 3519 8352 3528
rect 4344 3340 4396 3392
rect 8300 3485 8309 3519
rect 8309 3485 8343 3519
rect 8343 3485 8352 3519
rect 8300 3476 8352 3485
rect 10508 3519 10560 3528
rect 10508 3485 10517 3519
rect 10517 3485 10551 3519
rect 10551 3485 10560 3519
rect 10508 3476 10560 3485
rect 9588 3408 9640 3460
rect 22008 3680 22060 3732
rect 22192 3723 22244 3732
rect 22192 3689 22201 3723
rect 22201 3689 22235 3723
rect 22235 3689 22244 3723
rect 22192 3680 22244 3689
rect 22284 3680 22336 3732
rect 16120 3612 16172 3664
rect 16764 3587 16816 3596
rect 16764 3553 16773 3587
rect 16773 3553 16807 3587
rect 16807 3553 16816 3587
rect 16764 3544 16816 3553
rect 17408 3587 17460 3596
rect 17408 3553 17417 3587
rect 17417 3553 17451 3587
rect 17451 3553 17460 3587
rect 17408 3544 17460 3553
rect 19708 3587 19760 3596
rect 19708 3553 19717 3587
rect 19717 3553 19751 3587
rect 19751 3553 19760 3587
rect 19708 3544 19760 3553
rect 19892 3587 19944 3596
rect 19892 3553 19901 3587
rect 19901 3553 19935 3587
rect 19935 3553 19944 3587
rect 19892 3544 19944 3553
rect 20628 3587 20680 3596
rect 20628 3553 20637 3587
rect 20637 3553 20671 3587
rect 20671 3553 20680 3587
rect 20628 3544 20680 3553
rect 25964 3587 26016 3596
rect 25964 3553 25973 3587
rect 25973 3553 26007 3587
rect 26007 3553 26016 3587
rect 25964 3544 26016 3553
rect 26424 3587 26476 3596
rect 26424 3553 26433 3587
rect 26433 3553 26467 3587
rect 26467 3553 26476 3587
rect 26424 3544 26476 3553
rect 16120 3519 16172 3528
rect 16120 3485 16129 3519
rect 16129 3485 16163 3519
rect 16163 3485 16172 3519
rect 16120 3476 16172 3485
rect 22008 3476 22060 3528
rect 25320 3519 25372 3528
rect 17132 3408 17184 3460
rect 25320 3485 25329 3519
rect 25329 3485 25363 3519
rect 25363 3485 25372 3519
rect 25320 3476 25372 3485
rect 39304 3612 39356 3664
rect 40040 3612 40092 3664
rect 41236 3612 41288 3664
rect 40776 3587 40828 3596
rect 40776 3553 40785 3587
rect 40785 3553 40819 3587
rect 40819 3553 40828 3587
rect 40776 3544 40828 3553
rect 41420 3544 41472 3596
rect 32312 3476 32364 3528
rect 39948 3476 40000 3528
rect 42616 3476 42668 3528
rect 40960 3408 41012 3460
rect 44916 3680 44968 3732
rect 48320 3680 48372 3732
rect 46112 3587 46164 3596
rect 46112 3553 46121 3587
rect 46121 3553 46155 3587
rect 46155 3553 46164 3587
rect 46112 3544 46164 3553
rect 47032 3587 47084 3596
rect 47032 3553 47041 3587
rect 47041 3553 47075 3587
rect 47075 3553 47084 3587
rect 47032 3544 47084 3553
rect 44916 3476 44968 3528
rect 46572 3408 46624 3460
rect 5540 3340 5592 3392
rect 7472 3340 7524 3392
rect 13176 3340 13228 3392
rect 13268 3340 13320 3392
rect 18420 3340 18472 3392
rect 24952 3340 25004 3392
rect 27344 3340 27396 3392
rect 32496 3340 32548 3392
rect 45100 3340 45152 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 1952 3136 2004 3188
rect 5172 3136 5224 3188
rect 8300 3136 8352 3188
rect 19432 3136 19484 3188
rect 2044 3111 2096 3120
rect 2044 3077 2053 3111
rect 2053 3077 2087 3111
rect 2087 3077 2096 3111
rect 2044 3068 2096 3077
rect 4344 3111 4396 3120
rect 4344 3077 4353 3111
rect 4353 3077 4387 3111
rect 4387 3077 4396 3111
rect 4344 3068 4396 3077
rect 7472 3111 7524 3120
rect 7472 3077 7481 3111
rect 7481 3077 7515 3111
rect 7515 3077 7524 3111
rect 7472 3068 7524 3077
rect 13176 3111 13228 3120
rect 13176 3077 13185 3111
rect 13185 3077 13219 3111
rect 13219 3077 13228 3111
rect 13176 3068 13228 3077
rect 1860 3043 1912 3052
rect 1860 3009 1869 3043
rect 1869 3009 1903 3043
rect 1903 3009 1912 3043
rect 1860 3000 1912 3009
rect 7288 3043 7340 3052
rect 7288 3009 7297 3043
rect 7297 3009 7331 3043
rect 7331 3009 7340 3043
rect 7288 3000 7340 3009
rect 10508 3000 10560 3052
rect 12992 3043 13044 3052
rect 12992 3009 13001 3043
rect 13001 3009 13035 3043
rect 13035 3009 13044 3043
rect 12992 3000 13044 3009
rect 17316 3043 17368 3052
rect 17316 3009 17325 3043
rect 17325 3009 17359 3043
rect 17359 3009 17368 3043
rect 17316 3000 17368 3009
rect 20168 3068 20220 3120
rect 24952 3111 25004 3120
rect 24952 3077 24961 3111
rect 24961 3077 24995 3111
rect 24995 3077 25004 3111
rect 24952 3068 25004 3077
rect 27344 3111 27396 3120
rect 27344 3077 27353 3111
rect 27353 3077 27387 3111
rect 27387 3077 27396 3111
rect 27344 3068 27396 3077
rect 32496 3111 32548 3120
rect 32496 3077 32505 3111
rect 32505 3077 32539 3111
rect 32539 3077 32548 3111
rect 32496 3068 32548 3077
rect 40132 3111 40184 3120
rect 40132 3077 40141 3111
rect 40141 3077 40175 3111
rect 40175 3077 40184 3111
rect 40132 3068 40184 3077
rect 24768 3043 24820 3052
rect 24768 3009 24777 3043
rect 24777 3009 24811 3043
rect 24811 3009 24820 3043
rect 24768 3000 24820 3009
rect 27160 3043 27212 3052
rect 27160 3009 27169 3043
rect 27169 3009 27203 3043
rect 27203 3009 27212 3043
rect 27160 3000 27212 3009
rect 32312 3043 32364 3052
rect 32312 3009 32321 3043
rect 32321 3009 32355 3043
rect 32355 3009 32364 3043
rect 32312 3000 32364 3009
rect 39948 3043 40000 3052
rect 39948 3009 39957 3043
rect 39957 3009 39991 3043
rect 39991 3009 40000 3043
rect 39948 3000 40000 3009
rect 2780 2975 2832 2984
rect 2780 2941 2789 2975
rect 2789 2941 2823 2975
rect 2823 2941 2832 2975
rect 2780 2932 2832 2941
rect 4988 2932 5040 2984
rect 5172 2975 5224 2984
rect 5172 2941 5181 2975
rect 5181 2941 5215 2975
rect 5215 2941 5224 2975
rect 5172 2932 5224 2941
rect 7748 2975 7800 2984
rect 7748 2941 7757 2975
rect 7757 2941 7791 2975
rect 7791 2941 7800 2975
rect 7748 2932 7800 2941
rect 13544 2975 13596 2984
rect 13544 2941 13553 2975
rect 13553 2941 13587 2975
rect 13587 2941 13596 2975
rect 13544 2932 13596 2941
rect 18512 2932 18564 2984
rect 19340 2932 19392 2984
rect 19800 2975 19852 2984
rect 19800 2941 19809 2975
rect 19809 2941 19843 2975
rect 19843 2941 19852 2975
rect 19800 2932 19852 2941
rect 25780 2975 25832 2984
rect 25780 2941 25789 2975
rect 25789 2941 25823 2975
rect 25823 2941 25832 2975
rect 25780 2932 25832 2941
rect 27712 2975 27764 2984
rect 27712 2941 27721 2975
rect 27721 2941 27755 2975
rect 27755 2941 27764 2975
rect 27712 2932 27764 2941
rect 32220 2932 32272 2984
rect 40592 2975 40644 2984
rect 40592 2941 40601 2975
rect 40601 2941 40635 2975
rect 40635 2941 40644 2975
rect 40592 2932 40644 2941
rect 48964 3136 49016 3188
rect 45100 3111 45152 3120
rect 45100 3077 45109 3111
rect 45109 3077 45143 3111
rect 45143 3077 45152 3111
rect 45100 3068 45152 3077
rect 42616 3043 42668 3052
rect 42616 3009 42625 3043
rect 42625 3009 42659 3043
rect 42659 3009 42668 3043
rect 42616 3000 42668 3009
rect 44916 3043 44968 3052
rect 44916 3009 44925 3043
rect 44925 3009 44959 3043
rect 44959 3009 44968 3043
rect 44916 3000 44968 3009
rect 48044 3043 48096 3052
rect 48044 3009 48053 3043
rect 48053 3009 48087 3043
rect 48087 3009 48096 3043
rect 48044 3000 48096 3009
rect 42892 2932 42944 2984
rect 45744 2975 45796 2984
rect 41880 2864 41932 2916
rect 45744 2941 45753 2975
rect 45753 2941 45787 2975
rect 45787 2941 45796 2975
rect 45744 2932 45796 2941
rect 45100 2864 45152 2916
rect 45652 2864 45704 2916
rect 6828 2839 6880 2848
rect 6828 2805 6837 2839
rect 6837 2805 6871 2839
rect 6871 2805 6880 2839
rect 6828 2796 6880 2805
rect 28356 2796 28408 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 4620 2524 4672 2576
rect 4160 2499 4212 2508
rect 4160 2465 4169 2499
rect 4169 2465 4203 2499
rect 4203 2465 4212 2499
rect 4160 2456 4212 2465
rect 4528 2499 4580 2508
rect 4528 2465 4537 2499
rect 4537 2465 4571 2499
rect 4571 2465 4580 2499
rect 4528 2456 4580 2465
rect 6828 2456 6880 2508
rect 7104 2499 7156 2508
rect 7104 2465 7113 2499
rect 7113 2465 7147 2499
rect 7147 2465 7156 2499
rect 7104 2456 7156 2465
rect 17592 2592 17644 2644
rect 18512 2635 18564 2644
rect 18512 2601 18521 2635
rect 18521 2601 18555 2635
rect 18555 2601 18564 2635
rect 18512 2592 18564 2601
rect 19800 2592 19852 2644
rect 42892 2592 42944 2644
rect 47952 2635 48004 2644
rect 47952 2601 47961 2635
rect 47961 2601 47995 2635
rect 47995 2601 48004 2635
rect 47952 2592 48004 2601
rect 17776 2524 17828 2576
rect 25044 2524 25096 2576
rect 39580 2524 39632 2576
rect 26056 2456 26108 2508
rect 44640 2456 44692 2508
rect 46480 2456 46532 2508
rect 46848 2499 46900 2508
rect 46848 2465 46857 2499
rect 46857 2465 46891 2499
rect 46891 2465 46900 2499
rect 46848 2456 46900 2465
rect 11612 2388 11664 2440
rect 14188 2388 14240 2440
rect 18420 2431 18472 2440
rect 18420 2397 18429 2431
rect 18429 2397 18463 2431
rect 18463 2397 18472 2431
rect 18420 2388 18472 2397
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 19984 2388 20036 2440
rect 38660 2388 38712 2440
rect 41604 2431 41656 2440
rect 41604 2397 41613 2431
rect 41613 2397 41647 2431
rect 41647 2397 41656 2431
rect 41604 2388 41656 2397
rect 1308 2320 1360 2372
rect 2780 2320 2832 2372
rect 6828 2363 6880 2372
rect 6828 2329 6837 2363
rect 6837 2329 6871 2363
rect 6871 2329 6880 2363
rect 6828 2320 6880 2329
rect 25320 2320 25372 2372
rect 29000 2320 29052 2372
rect 43812 2320 43864 2372
rect 2872 2295 2924 2304
rect 2872 2261 2881 2295
rect 2881 2261 2915 2295
rect 2915 2261 2924 2295
rect 2872 2252 2924 2261
rect 23848 2252 23900 2304
rect 32864 2252 32916 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 2872 1980 2924 2032
rect 17500 1980 17552 2032
rect 2872 1844 2924 1896
rect 5356 1844 5408 1896
<< metal2 >>
rect -10 49200 102 49800
rect 1278 49314 1390 49800
rect 216 49286 1390 49314
rect 216 45554 244 49286
rect 1278 49200 1390 49286
rect 1922 49314 2034 49800
rect 1922 49286 2360 49314
rect 1922 49200 2034 49286
rect 2136 47048 2188 47054
rect 2136 46990 2188 46996
rect 2044 46504 2096 46510
rect 2044 46446 2096 46452
rect 2056 46170 2084 46446
rect 2044 46164 2096 46170
rect 2044 46106 2096 46112
rect 32 45526 244 45554
rect 32 44878 60 45526
rect 20 44872 72 44878
rect 20 44814 72 44820
rect 1768 44736 1820 44742
rect 1768 44678 1820 44684
rect 1584 43784 1636 43790
rect 1584 43726 1636 43732
rect 1596 43314 1624 43726
rect 1584 43308 1636 43314
rect 1584 43250 1636 43256
rect 1584 38956 1636 38962
rect 1584 38898 1636 38904
rect 1596 38865 1624 38898
rect 1582 38856 1638 38865
rect 1582 38791 1638 38800
rect 1584 37256 1636 37262
rect 1584 37198 1636 37204
rect 1596 36825 1624 37198
rect 1780 36922 1808 44678
rect 2148 42566 2176 46990
rect 2332 46510 2360 49286
rect 2566 49200 2678 49800
rect 3854 49200 3966 49800
rect 4498 49314 4610 49800
rect 4498 49286 4936 49314
rect 4498 49200 4610 49286
rect 2608 46646 2636 49200
rect 2778 48376 2834 48385
rect 2778 48311 2834 48320
rect 2596 46640 2648 46646
rect 2596 46582 2648 46588
rect 2320 46504 2372 46510
rect 2320 46446 2372 46452
rect 2792 46034 2820 48311
rect 2962 47696 3018 47705
rect 2962 47631 3018 47640
rect 2870 46336 2926 46345
rect 2870 46271 2926 46280
rect 2780 46028 2832 46034
rect 2780 45970 2832 45976
rect 2778 45656 2834 45665
rect 2778 45591 2834 45600
rect 2792 44334 2820 45591
rect 2320 44328 2372 44334
rect 2320 44270 2372 44276
rect 2780 44328 2832 44334
rect 2780 44270 2832 44276
rect 2332 42770 2360 44270
rect 2780 43852 2832 43858
rect 2780 43794 2832 43800
rect 2412 43716 2464 43722
rect 2412 43658 2464 43664
rect 2424 43450 2452 43658
rect 2792 43625 2820 43794
rect 2778 43616 2834 43625
rect 2778 43551 2834 43560
rect 2412 43444 2464 43450
rect 2412 43386 2464 43392
rect 2688 43308 2740 43314
rect 2688 43250 2740 43256
rect 2320 42764 2372 42770
rect 2320 42706 2372 42712
rect 2412 42696 2464 42702
rect 2412 42638 2464 42644
rect 2136 42560 2188 42566
rect 2136 42502 2188 42508
rect 2044 41608 2096 41614
rect 2044 41550 2096 41556
rect 2056 41138 2084 41550
rect 2044 41132 2096 41138
rect 2044 41074 2096 41080
rect 2320 41064 2372 41070
rect 2320 41006 2372 41012
rect 2332 40730 2360 41006
rect 2320 40724 2372 40730
rect 2320 40666 2372 40672
rect 1860 38752 1912 38758
rect 1860 38694 1912 38700
rect 1768 36916 1820 36922
rect 1768 36858 1820 36864
rect 1582 36816 1638 36825
rect 1582 36751 1638 36760
rect 1584 34604 1636 34610
rect 1584 34546 1636 34552
rect 1596 34105 1624 34546
rect 1768 34400 1820 34406
rect 1768 34342 1820 34348
rect 1780 34202 1808 34342
rect 1768 34196 1820 34202
rect 1768 34138 1820 34144
rect 1582 34096 1638 34105
rect 1582 34031 1638 34040
rect 1582 32056 1638 32065
rect 1582 31991 1638 32000
rect 1596 31890 1624 31991
rect 1584 31884 1636 31890
rect 1584 31826 1636 31832
rect 1872 30666 1900 38694
rect 2136 32904 2188 32910
rect 2136 32846 2188 32852
rect 2148 32434 2176 32846
rect 2320 32768 2372 32774
rect 2320 32710 2372 32716
rect 2332 32502 2360 32710
rect 2320 32496 2372 32502
rect 2320 32438 2372 32444
rect 2136 32428 2188 32434
rect 2136 32370 2188 32376
rect 1860 30660 1912 30666
rect 1860 30602 1912 30608
rect 2424 26234 2452 42638
rect 2596 40520 2648 40526
rect 2596 40462 2648 40468
rect 2504 32904 2556 32910
rect 2504 32846 2556 32852
rect 2240 26206 2452 26234
rect 2240 25906 2268 26206
rect 2228 25900 2280 25906
rect 2228 25842 2280 25848
rect 1768 25696 1820 25702
rect 1768 25638 1820 25644
rect 1780 25362 1808 25638
rect 1768 25356 1820 25362
rect 1768 25298 1820 25304
rect 1584 25288 1636 25294
rect 1584 25230 1636 25236
rect 1596 24818 1624 25230
rect 1584 24812 1636 24818
rect 1584 24754 1636 24760
rect 2044 22024 2096 22030
rect 2044 21966 2096 21972
rect 2056 21554 2084 21966
rect 2044 21548 2096 21554
rect 2044 21490 2096 21496
rect 2240 21026 2268 25842
rect 2516 21570 2544 32846
rect 2424 21542 2544 21570
rect 2320 21480 2372 21486
rect 2320 21422 2372 21428
rect 2332 21146 2360 21422
rect 2320 21140 2372 21146
rect 2320 21082 2372 21088
rect 2240 20998 2360 21026
rect 2332 20942 2360 20998
rect 2320 20936 2372 20942
rect 2320 20878 2372 20884
rect 204 19780 256 19786
rect 204 19722 256 19728
rect 216 16574 244 19722
rect 2044 18760 2096 18766
rect 2044 18702 2096 18708
rect 2056 18290 2084 18702
rect 2044 18284 2096 18290
rect 2044 18226 2096 18232
rect 2228 18216 2280 18222
rect 2228 18158 2280 18164
rect 2240 17882 2268 18158
rect 2228 17876 2280 17882
rect 2228 17818 2280 17824
rect 2332 17678 2360 20878
rect 2320 17672 2372 17678
rect 2320 17614 2372 17620
rect 1584 16992 1636 16998
rect 1584 16934 1636 16940
rect 1596 16658 1624 16934
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 2332 16574 2360 17614
rect 216 16546 704 16574
rect 676 800 704 16546
rect 2240 16546 2360 16574
rect 1584 15496 1636 15502
rect 1584 15438 1636 15444
rect 1596 15026 1624 15438
rect 1952 15428 2004 15434
rect 1952 15370 2004 15376
rect 1584 15020 1636 15026
rect 1584 14962 1636 14968
rect 1584 14408 1636 14414
rect 1584 14350 1636 14356
rect 1596 13938 1624 14350
rect 1768 14340 1820 14346
rect 1768 14282 1820 14288
rect 1780 14074 1808 14282
rect 1768 14068 1820 14074
rect 1768 14010 1820 14016
rect 1584 13932 1636 13938
rect 1584 13874 1636 13880
rect 1584 6792 1636 6798
rect 1584 6734 1636 6740
rect 1596 6322 1624 6734
rect 1768 6724 1820 6730
rect 1768 6666 1820 6672
rect 1780 6458 1808 6666
rect 1768 6452 1820 6458
rect 1768 6394 1820 6400
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 1860 5704 1912 5710
rect 1860 5646 1912 5652
rect 1768 5568 1820 5574
rect 1768 5510 1820 5516
rect 1780 4690 1808 5510
rect 1768 4684 1820 4690
rect 1768 4626 1820 4632
rect 1872 3058 1900 5646
rect 1964 3534 1992 15370
rect 2044 12232 2096 12238
rect 2044 12174 2096 12180
rect 2056 11762 2084 12174
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 2240 11150 2268 16546
rect 2424 16114 2452 21542
rect 2608 21434 2636 40462
rect 2516 21406 2636 21434
rect 2412 16108 2464 16114
rect 2412 16050 2464 16056
rect 2424 15434 2452 16050
rect 2412 15428 2464 15434
rect 2412 15370 2464 15376
rect 2516 15026 2544 21406
rect 2596 16516 2648 16522
rect 2596 16458 2648 16464
rect 2608 16250 2636 16458
rect 2596 16244 2648 16250
rect 2596 16186 2648 16192
rect 2504 15020 2556 15026
rect 2504 14962 2556 14968
rect 2320 11688 2372 11694
rect 2320 11630 2372 11636
rect 2332 11354 2360 11630
rect 2320 11348 2372 11354
rect 2320 11290 2372 11296
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2044 10056 2096 10062
rect 2044 9998 2096 10004
rect 2056 9586 2084 9998
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 2240 8974 2268 11086
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2332 9178 2360 9454
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 2056 7410 2084 7822
rect 2228 7744 2280 7750
rect 2228 7686 2280 7692
rect 2240 7478 2268 7686
rect 2228 7472 2280 7478
rect 2228 7414 2280 7420
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 2700 5710 2728 43250
rect 2884 42634 2912 46271
rect 2976 45422 3004 47631
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4160 47116 4212 47122
rect 4160 47058 4212 47064
rect 4068 47048 4120 47054
rect 4068 46990 4120 46996
rect 4080 45966 4108 46990
rect 4172 46578 4200 47058
rect 4804 46980 4856 46986
rect 4804 46922 4856 46928
rect 4160 46572 4212 46578
rect 4160 46514 4212 46520
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4068 45960 4120 45966
rect 4068 45902 4120 45908
rect 2964 45416 3016 45422
rect 2964 45358 3016 45364
rect 4080 44878 4108 45902
rect 4620 45892 4672 45898
rect 4620 45834 4672 45840
rect 4632 45626 4660 45834
rect 4620 45620 4672 45626
rect 4620 45562 4672 45568
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4068 44872 4120 44878
rect 4068 44814 4120 44820
rect 3792 44804 3844 44810
rect 3792 44746 3844 44752
rect 3056 44260 3108 44266
rect 3056 44202 3108 44208
rect 3068 42770 3096 44202
rect 3700 43784 3752 43790
rect 3700 43726 3752 43732
rect 3712 43314 3740 43726
rect 3700 43308 3752 43314
rect 3700 43250 3752 43256
rect 3148 43240 3200 43246
rect 3148 43182 3200 43188
rect 3056 42764 3108 42770
rect 3056 42706 3108 42712
rect 2872 42628 2924 42634
rect 2872 42570 2924 42576
rect 2778 41576 2834 41585
rect 2778 41511 2834 41520
rect 2792 41070 2820 41511
rect 2780 41064 2832 41070
rect 2780 41006 2832 41012
rect 2778 32736 2834 32745
rect 2778 32671 2834 32680
rect 2792 32366 2820 32671
rect 2780 32360 2832 32366
rect 2780 32302 2832 32308
rect 2780 25356 2832 25362
rect 2780 25298 2832 25304
rect 2792 25265 2820 25298
rect 2778 25256 2834 25265
rect 2778 25191 2834 25200
rect 2778 21856 2834 21865
rect 2778 21791 2834 21800
rect 2792 21486 2820 21791
rect 2780 21480 2832 21486
rect 2780 21422 2832 21428
rect 2962 20496 3018 20505
rect 2962 20431 3018 20440
rect 2976 20330 3004 20431
rect 2964 20324 3016 20330
rect 2964 20266 3016 20272
rect 2778 18456 2834 18465
rect 2778 18391 2834 18400
rect 2792 18222 2820 18391
rect 2780 18216 2832 18222
rect 2780 18158 2832 18164
rect 2778 17096 2834 17105
rect 2778 17031 2834 17040
rect 2792 16658 2820 17031
rect 2780 16652 2832 16658
rect 2780 16594 2832 16600
rect 3160 16574 3188 43182
rect 3514 40896 3570 40905
rect 3514 40831 3570 40840
rect 3528 20874 3556 40831
rect 3516 20868 3568 20874
rect 3516 20810 3568 20816
rect 2976 16546 3188 16574
rect 2780 15564 2832 15570
rect 2780 15506 2832 15512
rect 2792 15065 2820 15506
rect 2872 15360 2924 15366
rect 2872 15302 2924 15308
rect 2884 15162 2912 15302
rect 2872 15156 2924 15162
rect 2872 15098 2924 15104
rect 2778 15056 2834 15065
rect 2778 14991 2834 15000
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 2792 14385 2820 14418
rect 2778 14376 2834 14385
rect 2778 14311 2834 14320
rect 2976 13938 3004 16546
rect 3240 15020 3292 15026
rect 3240 14962 3292 14968
rect 2964 13932 3016 13938
rect 2964 13874 3016 13880
rect 2780 11688 2832 11694
rect 2778 11656 2780 11665
rect 2832 11656 2834 11665
rect 2778 11591 2834 11600
rect 2872 11008 2924 11014
rect 2872 10950 2924 10956
rect 2884 10742 2912 10950
rect 2872 10736 2924 10742
rect 2872 10678 2924 10684
rect 2778 9616 2834 9625
rect 2778 9551 2834 9560
rect 2792 9518 2820 9551
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 2778 7576 2834 7585
rect 2778 7511 2834 7520
rect 2792 7342 2820 7511
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 2976 6914 3004 13874
rect 3056 11144 3108 11150
rect 3056 11086 3108 11092
rect 3068 10606 3096 11086
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 3160 10305 3188 10542
rect 3146 10296 3202 10305
rect 3146 10231 3202 10240
rect 3252 7886 3280 14962
rect 3804 14414 3832 44746
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 3884 43988 3936 43994
rect 3884 43930 3936 43936
rect 3896 43246 3924 43930
rect 3884 43240 3936 43246
rect 3884 43182 3936 43188
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4632 42702 4660 45562
rect 4816 44418 4844 46922
rect 4908 45898 4936 49286
rect 5786 49200 5898 49800
rect 6430 49200 6542 49800
rect 7718 49200 7830 49800
rect 8362 49200 8474 49800
rect 9006 49200 9118 49800
rect 10294 49200 10406 49800
rect 10938 49200 11050 49800
rect 12226 49200 12338 49800
rect 12870 49200 12982 49800
rect 14158 49200 14270 49800
rect 14802 49200 14914 49800
rect 15446 49200 15558 49800
rect 16734 49200 16846 49800
rect 17378 49200 17490 49800
rect 18666 49200 18778 49800
rect 19310 49200 19422 49800
rect 20598 49200 20710 49800
rect 21242 49200 21354 49800
rect 21886 49200 21998 49800
rect 23174 49200 23286 49800
rect 23818 49200 23930 49800
rect 25106 49200 25218 49800
rect 25750 49200 25862 49800
rect 27038 49200 27150 49800
rect 27682 49200 27794 49800
rect 28970 49200 29082 49800
rect 29614 49200 29726 49800
rect 30258 49200 30370 49800
rect 31546 49200 31658 49800
rect 32190 49200 32302 49800
rect 33478 49200 33590 49800
rect 34122 49200 34234 49800
rect 35410 49200 35522 49800
rect 36054 49200 36166 49800
rect 36698 49200 36810 49800
rect 37986 49200 38098 49800
rect 38630 49200 38742 49800
rect 39918 49200 40030 49800
rect 40562 49200 40674 49800
rect 41850 49200 41962 49800
rect 42494 49200 42606 49800
rect 43138 49200 43250 49800
rect 44426 49200 44538 49800
rect 45070 49200 45182 49800
rect 46358 49200 46470 49800
rect 47002 49314 47114 49800
rect 47002 49286 47624 49314
rect 47002 49200 47114 49286
rect 5356 47048 5408 47054
rect 5356 46990 5408 46996
rect 5264 46368 5316 46374
rect 5264 46310 5316 46316
rect 5276 46034 5304 46310
rect 5264 46028 5316 46034
rect 5264 45970 5316 45976
rect 4896 45892 4948 45898
rect 4896 45834 4948 45840
rect 4896 45484 4948 45490
rect 4896 45426 4948 45432
rect 4908 44878 4936 45426
rect 4896 44872 4948 44878
rect 4896 44814 4948 44820
rect 4724 44390 4844 44418
rect 4908 44402 4936 44814
rect 5368 44810 5396 46990
rect 5632 46980 5684 46986
rect 5632 46922 5684 46928
rect 5540 46912 5592 46918
rect 5540 46854 5592 46860
rect 5552 46034 5580 46854
rect 5540 46028 5592 46034
rect 5540 45970 5592 45976
rect 5540 45892 5592 45898
rect 5540 45834 5592 45840
rect 5448 45416 5500 45422
rect 5448 45358 5500 45364
rect 5356 44804 5408 44810
rect 5356 44746 5408 44752
rect 5264 44736 5316 44742
rect 5264 44678 5316 44684
rect 4896 44396 4948 44402
rect 4724 43382 4752 44390
rect 4896 44338 4948 44344
rect 4804 44328 4856 44334
rect 4804 44270 4856 44276
rect 4712 43376 4764 43382
rect 4712 43318 4764 43324
rect 4620 42696 4672 42702
rect 4620 42638 4672 42644
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4712 31136 4764 31142
rect 4712 31078 4764 31084
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4724 29578 4752 31078
rect 4712 29572 4764 29578
rect 4712 29514 4764 29520
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4724 28218 4752 29514
rect 4712 28212 4764 28218
rect 4712 28154 4764 28160
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4066 23896 4122 23905
rect 4066 23831 4122 23840
rect 4080 23526 4108 23831
rect 4068 23520 4120 23526
rect 4068 23462 4120 23468
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4620 22160 4672 22166
rect 4620 22102 4672 22108
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4160 20936 4212 20942
rect 4160 20878 4212 20884
rect 4172 20466 4200 20878
rect 4160 20460 4212 20466
rect 4160 20402 4212 20408
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4632 15094 4660 22102
rect 4816 19854 4844 44270
rect 4908 43790 4936 44338
rect 4988 43852 5040 43858
rect 4988 43794 5040 43800
rect 4896 43784 4948 43790
rect 4896 43726 4948 43732
rect 5000 42226 5028 43794
rect 5080 42628 5132 42634
rect 5080 42570 5132 42576
rect 5092 42362 5120 42570
rect 5080 42356 5132 42362
rect 5080 42298 5132 42304
rect 4988 42220 5040 42226
rect 4988 42162 5040 42168
rect 5000 35894 5028 42162
rect 5000 35866 5120 35894
rect 4896 30048 4948 30054
rect 4896 29990 4948 29996
rect 4908 29646 4936 29990
rect 4896 29640 4948 29646
rect 4896 29582 4948 29588
rect 4988 28416 5040 28422
rect 4988 28358 5040 28364
rect 5000 28150 5028 28358
rect 4988 28144 5040 28150
rect 4988 28086 5040 28092
rect 4988 27872 5040 27878
rect 4988 27814 5040 27820
rect 5000 27674 5028 27814
rect 4988 27668 5040 27674
rect 4988 27610 5040 27616
rect 5092 20602 5120 35866
rect 5276 32910 5304 44678
rect 5368 44402 5396 44746
rect 5356 44396 5408 44402
rect 5356 44338 5408 44344
rect 5264 32904 5316 32910
rect 5264 32846 5316 32852
rect 5356 31136 5408 31142
rect 5356 31078 5408 31084
rect 5368 30938 5396 31078
rect 5356 30932 5408 30938
rect 5356 30874 5408 30880
rect 5172 30728 5224 30734
rect 5172 30670 5224 30676
rect 5184 30258 5212 30670
rect 5172 30252 5224 30258
rect 5172 30194 5224 30200
rect 5184 29170 5212 30194
rect 5172 29164 5224 29170
rect 5172 29106 5224 29112
rect 5184 27470 5212 29106
rect 5172 27464 5224 27470
rect 5172 27406 5224 27412
rect 5172 26988 5224 26994
rect 5224 26948 5304 26976
rect 5172 26930 5224 26936
rect 5276 26382 5304 26948
rect 5264 26376 5316 26382
rect 5264 26318 5316 26324
rect 5276 22166 5304 26318
rect 5264 22160 5316 22166
rect 5264 22102 5316 22108
rect 5080 20596 5132 20602
rect 5080 20538 5132 20544
rect 4896 20392 4948 20398
rect 4896 20334 4948 20340
rect 4908 20058 4936 20334
rect 4896 20052 4948 20058
rect 4896 19994 4948 20000
rect 4804 19848 4856 19854
rect 4804 19790 4856 19796
rect 4620 15088 4672 15094
rect 4620 15030 4672 15036
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 5356 14952 5408 14958
rect 5356 14894 5408 14900
rect 4080 14618 4108 14894
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 3792 14408 3844 14414
rect 3792 14350 3844 14356
rect 3804 11150 3832 14350
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 3792 11144 3844 11150
rect 3792 11086 3844 11092
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 2778 6896 2834 6905
rect 2778 6831 2780 6840
rect 2832 6831 2834 6840
rect 2884 6886 3004 6914
rect 2780 6802 2832 6808
rect 2884 6322 2912 6886
rect 2872 6316 2924 6322
rect 2872 6258 2924 6264
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 2688 5704 2740 5710
rect 2688 5646 2740 5652
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 2964 5160 3016 5166
rect 2964 5102 3016 5108
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 2044 3936 2096 3942
rect 2044 3878 2096 3884
rect 1952 3528 2004 3534
rect 1952 3470 2004 3476
rect 1964 3194 1992 3470
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 2056 3126 2084 3878
rect 2792 3505 2820 4626
rect 2884 4146 2912 5102
rect 2976 4865 3004 5102
rect 2962 4856 3018 4865
rect 2962 4791 3018 4800
rect 3160 4758 3188 5646
rect 3514 5536 3570 5545
rect 3514 5471 3570 5480
rect 3148 4752 3200 4758
rect 3148 4694 3200 4700
rect 3528 4690 3556 5471
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 3516 4684 3568 4690
rect 3516 4626 3568 4632
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4988 4616 5040 4622
rect 4988 4558 5040 4564
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 3976 4072 4028 4078
rect 3976 4014 4028 4020
rect 2976 3738 3004 4014
rect 3240 4004 3292 4010
rect 3240 3946 3292 3952
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 2778 3496 2834 3505
rect 2778 3431 2834 3440
rect 2044 3120 2096 3126
rect 2044 3062 2096 3068
rect 1860 3052 1912 3058
rect 1860 2994 1912 3000
rect 2780 2984 2832 2990
rect 2780 2926 2832 2932
rect 2792 2825 2820 2926
rect 2778 2816 2834 2825
rect 2778 2751 2834 2760
rect 1308 2372 1360 2378
rect 1308 2314 1360 2320
rect 2780 2372 2832 2378
rect 2780 2314 2832 2320
rect 1320 800 1348 2314
rect -10 200 102 800
rect 634 200 746 800
rect 1278 200 1390 800
rect 2566 200 2678 800
rect 2792 785 2820 2314
rect 2872 2304 2924 2310
rect 2872 2246 2924 2252
rect 2884 2038 2912 2246
rect 2872 2032 2924 2038
rect 2872 1974 2924 1980
rect 2872 1896 2924 1902
rect 2872 1838 2924 1844
rect 2884 1465 2912 1838
rect 2870 1456 2926 1465
rect 2870 1391 2926 1400
rect 3252 800 3280 3946
rect 3988 3738 4016 4014
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4172 2938 4200 3470
rect 4344 3392 4396 3398
rect 4344 3334 4396 3340
rect 4356 3126 4384 3334
rect 4344 3120 4396 3126
rect 4344 3062 4396 3068
rect 4080 2910 4200 2938
rect 4080 2530 4108 2910
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2582 4660 4558
rect 5000 2990 5028 4558
rect 5172 3664 5224 3670
rect 5172 3606 5224 3612
rect 5184 3194 5212 3606
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 4620 2576 4672 2582
rect 4080 2514 4200 2530
rect 4620 2518 4672 2524
rect 4080 2508 4212 2514
rect 4080 2502 4160 2508
rect 4160 2450 4212 2456
rect 4528 2508 4580 2514
rect 4528 2450 4580 2456
rect 4540 800 4568 2450
rect 5184 800 5212 2926
rect 5368 1902 5396 14894
rect 5460 3602 5488 45358
rect 5552 42770 5580 45834
rect 5644 45558 5672 46922
rect 5828 46034 5856 49200
rect 9048 47122 9076 49200
rect 7196 47116 7248 47122
rect 7196 47058 7248 47064
rect 9036 47116 9088 47122
rect 9036 47058 9088 47064
rect 6552 47048 6604 47054
rect 6552 46990 6604 46996
rect 5908 46504 5960 46510
rect 5908 46446 5960 46452
rect 5816 46028 5868 46034
rect 5816 45970 5868 45976
rect 5920 45558 5948 46446
rect 5632 45552 5684 45558
rect 5632 45494 5684 45500
rect 5908 45552 5960 45558
rect 5908 45494 5960 45500
rect 6564 43994 6592 46990
rect 6920 45960 6972 45966
rect 6920 45902 6972 45908
rect 6932 45506 6960 45902
rect 6840 45478 6960 45506
rect 7208 45490 7236 47058
rect 7380 47048 7432 47054
rect 7380 46990 7432 46996
rect 8852 47048 8904 47054
rect 8852 46990 8904 46996
rect 7288 45824 7340 45830
rect 7288 45766 7340 45772
rect 7300 45558 7328 45766
rect 7288 45552 7340 45558
rect 7288 45494 7340 45500
rect 7196 45484 7248 45490
rect 6840 44946 6868 45478
rect 7196 45426 7248 45432
rect 7392 45354 7420 46990
rect 8024 46368 8076 46374
rect 8024 46310 8076 46316
rect 8036 46102 8064 46310
rect 8024 46096 8076 46102
rect 8024 46038 8076 46044
rect 7380 45348 7432 45354
rect 7380 45290 7432 45296
rect 6828 44940 6880 44946
rect 6828 44882 6880 44888
rect 6552 43988 6604 43994
rect 6552 43930 6604 43936
rect 5540 42764 5592 42770
rect 5540 42706 5592 42712
rect 6644 31816 6696 31822
rect 6644 31758 6696 31764
rect 6000 31340 6052 31346
rect 6000 31282 6052 31288
rect 6012 30938 6040 31282
rect 6000 30932 6052 30938
rect 6000 30874 6052 30880
rect 6184 30728 6236 30734
rect 6184 30670 6236 30676
rect 5540 30592 5592 30598
rect 5540 30534 5592 30540
rect 5552 30394 5580 30534
rect 6196 30394 6224 30670
rect 5540 30388 5592 30394
rect 5540 30330 5592 30336
rect 6184 30388 6236 30394
rect 6184 30330 6236 30336
rect 6656 30326 6684 31758
rect 6644 30320 6696 30326
rect 6644 30262 6696 30268
rect 5724 29504 5776 29510
rect 5724 29446 5776 29452
rect 5736 29034 5764 29446
rect 5724 29028 5776 29034
rect 5724 28970 5776 28976
rect 5632 28960 5684 28966
rect 5632 28902 5684 28908
rect 5644 28558 5672 28902
rect 5632 28552 5684 28558
rect 5632 28494 5684 28500
rect 5724 27668 5776 27674
rect 5724 27610 5776 27616
rect 5736 27130 5764 27610
rect 5908 27328 5960 27334
rect 5908 27270 5960 27276
rect 6368 27328 6420 27334
rect 6368 27270 6420 27276
rect 5724 27124 5776 27130
rect 5724 27066 5776 27072
rect 5920 26994 5948 27270
rect 6380 27062 6408 27270
rect 6368 27056 6420 27062
rect 6368 26998 6420 27004
rect 5908 26988 5960 26994
rect 5908 26930 5960 26936
rect 6552 26784 6604 26790
rect 6552 26726 6604 26732
rect 6564 26382 6592 26726
rect 6552 26376 6604 26382
rect 6552 26318 6604 26324
rect 5540 19848 5592 19854
rect 5540 19790 5592 19796
rect 5552 4622 5580 19790
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5552 4146 5580 4558
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 5552 3398 5580 4082
rect 5644 3942 5672 7822
rect 6840 6914 6868 44882
rect 8392 31340 8444 31346
rect 8392 31282 8444 31288
rect 8208 31136 8260 31142
rect 8208 31078 8260 31084
rect 6920 30796 6972 30802
rect 6920 30738 6972 30744
rect 6932 29714 6960 30738
rect 8220 30734 8248 31078
rect 8208 30728 8260 30734
rect 8208 30670 8260 30676
rect 7840 30592 7892 30598
rect 7840 30534 7892 30540
rect 7392 30258 7788 30274
rect 7852 30258 7880 30534
rect 8404 30394 8432 31282
rect 8392 30388 8444 30394
rect 8392 30330 8444 30336
rect 7380 30252 7788 30258
rect 7432 30246 7788 30252
rect 7380 30194 7432 30200
rect 7760 30190 7788 30246
rect 7840 30252 7892 30258
rect 7840 30194 7892 30200
rect 8668 30252 8720 30258
rect 8668 30194 8720 30200
rect 7748 30184 7800 30190
rect 7748 30126 7800 30132
rect 7472 30116 7524 30122
rect 7472 30058 7524 30064
rect 6920 29708 6972 29714
rect 6920 29650 6972 29656
rect 6932 29578 6960 29650
rect 6920 29572 6972 29578
rect 6920 29514 6972 29520
rect 7288 29572 7340 29578
rect 7288 29514 7340 29520
rect 6932 28150 6960 29514
rect 7300 29306 7328 29514
rect 7288 29300 7340 29306
rect 7288 29242 7340 29248
rect 7484 29170 7512 30058
rect 7760 29186 7788 30126
rect 7852 29306 7880 30194
rect 8392 30048 8444 30054
rect 8392 29990 8444 29996
rect 8300 29504 8352 29510
rect 8300 29446 8352 29452
rect 7840 29300 7892 29306
rect 7840 29242 7892 29248
rect 7760 29170 7880 29186
rect 7472 29164 7524 29170
rect 7760 29164 7892 29170
rect 7760 29158 7840 29164
rect 7472 29106 7524 29112
rect 7840 29106 7892 29112
rect 8312 28966 8340 29446
rect 8404 29102 8432 29990
rect 8680 29306 8708 30194
rect 8668 29300 8720 29306
rect 8668 29242 8720 29248
rect 8392 29096 8444 29102
rect 8392 29038 8444 29044
rect 8300 28960 8352 28966
rect 8300 28902 8352 28908
rect 6920 28144 6972 28150
rect 6920 28086 6972 28092
rect 8864 28014 8892 46990
rect 10048 45620 10100 45626
rect 10048 45562 10100 45568
rect 10060 44402 10088 45562
rect 10980 45554 11008 49200
rect 12716 47048 12768 47054
rect 12716 46990 12768 46996
rect 12728 46646 12756 46990
rect 12716 46640 12768 46646
rect 12716 46582 12768 46588
rect 12912 46510 12940 49200
rect 14200 47122 14228 49200
rect 14188 47116 14240 47122
rect 14188 47058 14240 47064
rect 13820 46980 13872 46986
rect 13820 46922 13872 46928
rect 12532 46504 12584 46510
rect 12532 46446 12584 46452
rect 12900 46504 12952 46510
rect 12900 46446 12952 46452
rect 12544 46170 12572 46446
rect 13832 46170 13860 46922
rect 14844 46510 14872 49200
rect 14280 46504 14332 46510
rect 14280 46446 14332 46452
rect 14464 46504 14516 46510
rect 14464 46446 14516 46452
rect 14832 46504 14884 46510
rect 14832 46446 14884 46452
rect 12532 46164 12584 46170
rect 12532 46106 12584 46112
rect 13820 46164 13872 46170
rect 13820 46106 13872 46112
rect 12440 45960 12492 45966
rect 12440 45902 12492 45908
rect 10980 45526 11100 45554
rect 10508 45280 10560 45286
rect 10508 45222 10560 45228
rect 10520 44946 10548 45222
rect 11072 44946 11100 45526
rect 10508 44940 10560 44946
rect 10508 44882 10560 44888
rect 11060 44940 11112 44946
rect 11060 44882 11112 44888
rect 10692 44804 10744 44810
rect 10692 44746 10744 44752
rect 10704 44538 10732 44746
rect 12452 44742 12480 45902
rect 14292 45490 14320 46446
rect 14476 46170 14504 46446
rect 15016 46368 15068 46374
rect 15016 46310 15068 46316
rect 14464 46164 14516 46170
rect 14464 46106 14516 46112
rect 15028 46034 15056 46310
rect 15488 46034 15516 49200
rect 17420 47054 17448 49200
rect 17960 47184 18012 47190
rect 17960 47126 18012 47132
rect 17408 47048 17460 47054
rect 17408 46990 17460 46996
rect 15016 46028 15068 46034
rect 15016 45970 15068 45976
rect 15476 46028 15528 46034
rect 15476 45970 15528 45976
rect 15200 45892 15252 45898
rect 15200 45834 15252 45840
rect 15212 45626 15240 45834
rect 15200 45620 15252 45626
rect 15200 45562 15252 45568
rect 14280 45484 14332 45490
rect 14280 45426 14332 45432
rect 15200 45484 15252 45490
rect 15200 45426 15252 45432
rect 15212 45354 15240 45426
rect 15200 45348 15252 45354
rect 15200 45290 15252 45296
rect 12440 44736 12492 44742
rect 12440 44678 12492 44684
rect 10692 44532 10744 44538
rect 10692 44474 10744 44480
rect 10048 44396 10100 44402
rect 10048 44338 10100 44344
rect 15212 43994 15240 45290
rect 15200 43988 15252 43994
rect 15200 43930 15252 43936
rect 17132 43240 17184 43246
rect 17132 43182 17184 43188
rect 17408 43240 17460 43246
rect 17408 43182 17460 43188
rect 14004 42696 14056 42702
rect 14004 42638 14056 42644
rect 14016 42294 14044 42638
rect 15200 42560 15252 42566
rect 15200 42502 15252 42508
rect 16120 42560 16172 42566
rect 16120 42502 16172 42508
rect 14004 42288 14056 42294
rect 14004 42230 14056 42236
rect 14924 42016 14976 42022
rect 14924 41958 14976 41964
rect 14936 41614 14964 41958
rect 14924 41608 14976 41614
rect 14924 41550 14976 41556
rect 14740 41472 14792 41478
rect 14740 41414 14792 41420
rect 14752 41206 14780 41414
rect 15212 41274 15240 42502
rect 16132 42362 16160 42502
rect 16120 42356 16172 42362
rect 16120 42298 16172 42304
rect 16132 42158 16160 42298
rect 17144 42226 17172 43182
rect 17420 42906 17448 43182
rect 17408 42900 17460 42906
rect 17408 42842 17460 42848
rect 17132 42220 17184 42226
rect 17132 42162 17184 42168
rect 16028 42152 16080 42158
rect 16028 42094 16080 42100
rect 16120 42152 16172 42158
rect 16120 42094 16172 42100
rect 15476 42084 15528 42090
rect 15476 42026 15528 42032
rect 15488 41682 15516 42026
rect 15476 41676 15528 41682
rect 15476 41618 15528 41624
rect 15936 41540 15988 41546
rect 15936 41482 15988 41488
rect 15200 41268 15252 41274
rect 15200 41210 15252 41216
rect 14740 41200 14792 41206
rect 14740 41142 14792 41148
rect 14096 41064 14148 41070
rect 14096 41006 14148 41012
rect 14108 39506 14136 41006
rect 15948 40730 15976 41482
rect 16040 41138 16068 42094
rect 17144 41818 17172 42162
rect 17684 42152 17736 42158
rect 17684 42094 17736 42100
rect 17696 41818 17724 42094
rect 17132 41812 17184 41818
rect 17132 41754 17184 41760
rect 17500 41812 17552 41818
rect 17500 41754 17552 41760
rect 17684 41812 17736 41818
rect 17684 41754 17736 41760
rect 17144 41546 17172 41754
rect 17408 41744 17460 41750
rect 17408 41686 17460 41692
rect 17132 41540 17184 41546
rect 17132 41482 17184 41488
rect 17144 41414 17172 41482
rect 17420 41478 17448 41686
rect 17408 41472 17460 41478
rect 17408 41414 17460 41420
rect 17052 41386 17172 41414
rect 17328 41386 17448 41414
rect 17052 41138 17080 41386
rect 17328 41138 17356 41386
rect 16028 41132 16080 41138
rect 16028 41074 16080 41080
rect 17040 41132 17092 41138
rect 17040 41074 17092 41080
rect 17316 41132 17368 41138
rect 17316 41074 17368 41080
rect 16040 40730 16068 41074
rect 16120 40928 16172 40934
rect 16120 40870 16172 40876
rect 15936 40724 15988 40730
rect 15936 40666 15988 40672
rect 16028 40724 16080 40730
rect 16028 40666 16080 40672
rect 16132 40526 16160 40870
rect 16948 40588 17000 40594
rect 16948 40530 17000 40536
rect 16120 40520 16172 40526
rect 16120 40462 16172 40468
rect 14096 39500 14148 39506
rect 14096 39442 14148 39448
rect 14280 39500 14332 39506
rect 14280 39442 14332 39448
rect 13912 39364 13964 39370
rect 13912 39306 13964 39312
rect 13924 39098 13952 39306
rect 13912 39092 13964 39098
rect 13912 39034 13964 39040
rect 14292 38962 14320 39442
rect 15200 39296 15252 39302
rect 15200 39238 15252 39244
rect 14096 38956 14148 38962
rect 14096 38898 14148 38904
rect 14280 38956 14332 38962
rect 14280 38898 14332 38904
rect 14108 38554 14136 38898
rect 14372 38888 14424 38894
rect 14372 38830 14424 38836
rect 14096 38548 14148 38554
rect 14096 38490 14148 38496
rect 12900 37868 12952 37874
rect 12900 37810 12952 37816
rect 12624 37664 12676 37670
rect 12624 37606 12676 37612
rect 12636 37262 12664 37606
rect 12348 37256 12400 37262
rect 12348 37198 12400 37204
rect 12624 37256 12676 37262
rect 12624 37198 12676 37204
rect 12360 36174 12388 37198
rect 12440 37188 12492 37194
rect 12440 37130 12492 37136
rect 11796 36168 11848 36174
rect 11796 36110 11848 36116
rect 12348 36168 12400 36174
rect 12348 36110 12400 36116
rect 11808 34066 11836 36110
rect 11796 34060 11848 34066
rect 11796 34002 11848 34008
rect 11808 33590 11836 34002
rect 12072 33924 12124 33930
rect 12072 33866 12124 33872
rect 12084 33658 12112 33866
rect 12072 33652 12124 33658
rect 12072 33594 12124 33600
rect 11796 33584 11848 33590
rect 11796 33526 11848 33532
rect 11808 31346 11836 33526
rect 12164 33516 12216 33522
rect 12164 33458 12216 33464
rect 12176 33114 12204 33458
rect 12452 33454 12480 37130
rect 12912 36922 12940 37810
rect 13636 37120 13688 37126
rect 13636 37062 13688 37068
rect 13648 36922 13676 37062
rect 12900 36916 12952 36922
rect 12900 36858 12952 36864
rect 13636 36916 13688 36922
rect 13636 36858 13688 36864
rect 12808 36100 12860 36106
rect 12808 36042 12860 36048
rect 12820 35834 12848 36042
rect 12808 35828 12860 35834
rect 12808 35770 12860 35776
rect 13648 35766 13676 36858
rect 14096 36712 14148 36718
rect 14096 36654 14148 36660
rect 13820 36032 13872 36038
rect 13820 35974 13872 35980
rect 13832 35834 13860 35974
rect 13820 35828 13872 35834
rect 13820 35770 13872 35776
rect 13636 35760 13688 35766
rect 13636 35702 13688 35708
rect 13648 35086 13676 35702
rect 13728 35692 13780 35698
rect 13728 35634 13780 35640
rect 13740 35086 13768 35634
rect 13832 35154 13860 35770
rect 14108 35630 14136 36654
rect 14096 35624 14148 35630
rect 14096 35566 14148 35572
rect 13820 35148 13872 35154
rect 13820 35090 13872 35096
rect 13636 35080 13688 35086
rect 13636 35022 13688 35028
rect 13728 35080 13780 35086
rect 13728 35022 13780 35028
rect 13740 34202 13768 35022
rect 12992 34196 13044 34202
rect 12992 34138 13044 34144
rect 13728 34196 13780 34202
rect 13728 34138 13780 34144
rect 12440 33448 12492 33454
rect 12440 33390 12492 33396
rect 12808 33448 12860 33454
rect 12808 33390 12860 33396
rect 12532 33312 12584 33318
rect 12532 33254 12584 33260
rect 12164 33108 12216 33114
rect 12164 33050 12216 33056
rect 12440 31680 12492 31686
rect 12440 31622 12492 31628
rect 12452 31414 12480 31622
rect 12440 31408 12492 31414
rect 12440 31350 12492 31356
rect 11796 31340 11848 31346
rect 11796 31282 11848 31288
rect 12544 30938 12572 33254
rect 12624 32904 12676 32910
rect 12624 32846 12676 32852
rect 12636 31754 12664 32846
rect 12636 31726 12756 31754
rect 12624 31408 12676 31414
rect 12624 31350 12676 31356
rect 12532 30932 12584 30938
rect 12532 30874 12584 30880
rect 9128 30796 9180 30802
rect 9128 30738 9180 30744
rect 9140 30598 9168 30738
rect 12636 30734 12664 31350
rect 12440 30728 12492 30734
rect 12440 30670 12492 30676
rect 12624 30728 12676 30734
rect 12624 30670 12676 30676
rect 9496 30660 9548 30666
rect 9496 30602 9548 30608
rect 9128 30592 9180 30598
rect 9128 30534 9180 30540
rect 9508 30394 9536 30602
rect 10508 30592 10560 30598
rect 10508 30534 10560 30540
rect 12256 30592 12308 30598
rect 12256 30534 12308 30540
rect 9496 30388 9548 30394
rect 9496 30330 9548 30336
rect 10520 30054 10548 30534
rect 11888 30320 11940 30326
rect 11888 30262 11940 30268
rect 10508 30048 10560 30054
rect 10508 29990 10560 29996
rect 9220 29096 9272 29102
rect 9220 29038 9272 29044
rect 9232 28762 9260 29038
rect 9220 28756 9272 28762
rect 9220 28698 9272 28704
rect 9404 28552 9456 28558
rect 9404 28494 9456 28500
rect 9416 28082 9444 28494
rect 9404 28076 9456 28082
rect 9404 28018 9456 28024
rect 8852 28008 8904 28014
rect 8852 27950 8904 27956
rect 8024 27872 8076 27878
rect 8024 27814 8076 27820
rect 7012 27396 7064 27402
rect 7012 27338 7064 27344
rect 6920 26512 6972 26518
rect 6920 26454 6972 26460
rect 6932 25702 6960 26454
rect 7024 25906 7052 27338
rect 7564 27328 7616 27334
rect 7564 27270 7616 27276
rect 7576 26994 7604 27270
rect 7564 26988 7616 26994
rect 7564 26930 7616 26936
rect 8036 26926 8064 27814
rect 8392 27668 8444 27674
rect 8392 27610 8444 27616
rect 7104 26920 7156 26926
rect 7104 26862 7156 26868
rect 8024 26920 8076 26926
rect 8024 26862 8076 26868
rect 7116 26382 7144 26862
rect 8404 26586 8432 27610
rect 9416 27130 9444 28018
rect 9588 27940 9640 27946
rect 9588 27882 9640 27888
rect 9404 27124 9456 27130
rect 9404 27066 9456 27072
rect 8392 26580 8444 26586
rect 8392 26522 8444 26528
rect 7104 26376 7156 26382
rect 7104 26318 7156 26324
rect 7748 26308 7800 26314
rect 7748 26250 7800 26256
rect 7760 26042 7788 26250
rect 7748 26036 7800 26042
rect 7748 25978 7800 25984
rect 7012 25900 7064 25906
rect 7012 25842 7064 25848
rect 6920 25696 6972 25702
rect 6920 25638 6972 25644
rect 9600 21554 9628 27882
rect 11900 23798 11928 30262
rect 12268 30258 12296 30534
rect 12256 30252 12308 30258
rect 12256 30194 12308 30200
rect 11980 30184 12032 30190
rect 11980 30126 12032 30132
rect 11992 27538 12020 30126
rect 12452 29850 12480 30670
rect 12440 29844 12492 29850
rect 12440 29786 12492 29792
rect 11980 27532 12032 27538
rect 11980 27474 12032 27480
rect 11992 25362 12020 27474
rect 12532 27396 12584 27402
rect 12532 27338 12584 27344
rect 12544 27130 12572 27338
rect 12532 27124 12584 27130
rect 12532 27066 12584 27072
rect 12532 25696 12584 25702
rect 12532 25638 12584 25644
rect 11980 25356 12032 25362
rect 11980 25298 12032 25304
rect 12348 25220 12400 25226
rect 12348 25162 12400 25168
rect 12360 24954 12388 25162
rect 12348 24948 12400 24954
rect 12348 24890 12400 24896
rect 12544 24818 12572 25638
rect 12532 24812 12584 24818
rect 12532 24754 12584 24760
rect 11888 23792 11940 23798
rect 11888 23734 11940 23740
rect 11060 23520 11112 23526
rect 11060 23462 11112 23468
rect 11072 23186 11100 23462
rect 11060 23180 11112 23186
rect 11060 23122 11112 23128
rect 10140 23112 10192 23118
rect 10140 23054 10192 23060
rect 9588 21548 9640 21554
rect 9588 21490 9640 21496
rect 10048 21412 10100 21418
rect 10048 21354 10100 21360
rect 10060 20942 10088 21354
rect 10048 20936 10100 20942
rect 10048 20878 10100 20884
rect 9588 20596 9640 20602
rect 9588 20538 9640 20544
rect 9600 19854 9628 20538
rect 9588 19848 9640 19854
rect 9588 19790 9640 19796
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 6564 6886 6868 6914
rect 6276 4548 6328 4554
rect 6276 4490 6328 4496
rect 6288 3942 6316 4490
rect 6564 4078 6592 6886
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 6564 3602 6592 4014
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 6552 3596 6604 3602
rect 6552 3538 6604 3544
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5356 1896 5408 1902
rect 5356 1838 5408 1844
rect 6472 800 6500 3538
rect 6748 2394 6776 3878
rect 7300 3058 7328 3878
rect 8312 3534 8340 8910
rect 9600 3738 9628 19790
rect 9956 19372 10008 19378
rect 9956 19314 10008 19320
rect 9968 18698 9996 19314
rect 10060 19310 10088 20878
rect 10152 20398 10180 23054
rect 10508 23044 10560 23050
rect 10508 22986 10560 22992
rect 10520 22778 10548 22986
rect 10508 22772 10560 22778
rect 10508 22714 10560 22720
rect 10416 22636 10468 22642
rect 10416 22578 10468 22584
rect 12532 22636 12584 22642
rect 12532 22578 12584 22584
rect 10428 21593 10456 22578
rect 12164 22568 12216 22574
rect 12164 22510 12216 22516
rect 11520 22160 11572 22166
rect 11520 22102 11572 22108
rect 10414 21584 10470 21593
rect 10414 21519 10416 21528
rect 10468 21519 10470 21528
rect 10416 21490 10468 21496
rect 10324 21480 10376 21486
rect 10324 21422 10376 21428
rect 10232 21344 10284 21350
rect 10232 21286 10284 21292
rect 10244 21010 10272 21286
rect 10232 21004 10284 21010
rect 10232 20946 10284 20952
rect 10336 20398 10364 21422
rect 10140 20392 10192 20398
rect 10140 20334 10192 20340
rect 10324 20392 10376 20398
rect 10324 20334 10376 20340
rect 10048 19304 10100 19310
rect 10048 19246 10100 19252
rect 9956 18692 10008 18698
rect 9956 18634 10008 18640
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9784 4690 9812 5646
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 10060 4690 10088 5510
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7484 3126 7512 3334
rect 8312 3194 8340 3470
rect 9600 3466 9628 3674
rect 9876 3670 9904 4082
rect 10152 4010 10180 20334
rect 10232 19848 10284 19854
rect 10232 19790 10284 19796
rect 10244 19310 10272 19790
rect 11532 19378 11560 22102
rect 12176 21350 12204 22510
rect 12544 22234 12572 22578
rect 12532 22228 12584 22234
rect 12532 22170 12584 22176
rect 12440 21548 12492 21554
rect 12440 21490 12492 21496
rect 12164 21344 12216 21350
rect 12164 21286 12216 21292
rect 12176 20942 12204 21286
rect 12164 20936 12216 20942
rect 12164 20878 12216 20884
rect 11520 19372 11572 19378
rect 11520 19314 11572 19320
rect 11796 19372 11848 19378
rect 11796 19314 11848 19320
rect 10232 19304 10284 19310
rect 10232 19246 10284 19252
rect 11532 17746 11560 19314
rect 11808 18970 11836 19314
rect 11796 18964 11848 18970
rect 11796 18906 11848 18912
rect 11520 17740 11572 17746
rect 11520 17682 11572 17688
rect 11532 17270 11560 17682
rect 12072 17604 12124 17610
rect 12072 17546 12124 17552
rect 12084 17338 12112 17546
rect 12072 17332 12124 17338
rect 12072 17274 12124 17280
rect 11520 17264 11572 17270
rect 11520 17206 11572 17212
rect 12176 16114 12204 20878
rect 12452 20602 12480 21490
rect 12440 20596 12492 20602
rect 12440 20538 12492 20544
rect 12532 20460 12584 20466
rect 12532 20402 12584 20408
rect 12544 19514 12572 20402
rect 12532 19508 12584 19514
rect 12532 19450 12584 19456
rect 12544 18766 12572 19450
rect 12256 18760 12308 18766
rect 12256 18702 12308 18708
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12268 18426 12296 18702
rect 12256 18420 12308 18426
rect 12256 18362 12308 18368
rect 12636 18154 12664 30670
rect 12728 29646 12756 31726
rect 12716 29640 12768 29646
rect 12716 29582 12768 29588
rect 12728 27962 12756 29582
rect 12820 28082 12848 33390
rect 13004 32910 13032 34138
rect 13820 33312 13872 33318
rect 13820 33254 13872 33260
rect 12992 32904 13044 32910
rect 12992 32846 13044 32852
rect 13832 32842 13860 33254
rect 12900 32836 12952 32842
rect 12900 32778 12952 32784
rect 13820 32836 13872 32842
rect 13820 32778 13872 32784
rect 12912 32570 12940 32778
rect 12900 32564 12952 32570
rect 12900 32506 12952 32512
rect 12912 29646 12940 32506
rect 13820 31816 13872 31822
rect 13820 31758 13872 31764
rect 13832 31482 13860 31758
rect 13820 31476 13872 31482
rect 13820 31418 13872 31424
rect 14108 31278 14136 35566
rect 14280 33516 14332 33522
rect 14280 33458 14332 33464
rect 14292 33114 14320 33458
rect 14280 33108 14332 33114
rect 14280 33050 14332 33056
rect 14384 32978 14412 38830
rect 15212 38350 15240 39238
rect 15476 38956 15528 38962
rect 15476 38898 15528 38904
rect 15200 38344 15252 38350
rect 15200 38286 15252 38292
rect 15212 36174 15240 38286
rect 15384 38208 15436 38214
rect 15384 38150 15436 38156
rect 15396 37874 15424 38150
rect 15488 38010 15516 38898
rect 15568 38752 15620 38758
rect 15568 38694 15620 38700
rect 16120 38752 16172 38758
rect 16120 38694 16172 38700
rect 15476 38004 15528 38010
rect 15476 37946 15528 37952
rect 15580 37874 15608 38694
rect 16132 38350 16160 38694
rect 16120 38344 16172 38350
rect 16120 38286 16172 38292
rect 16856 38344 16908 38350
rect 16856 38286 16908 38292
rect 15384 37868 15436 37874
rect 15384 37810 15436 37816
rect 15568 37868 15620 37874
rect 15568 37810 15620 37816
rect 15660 37800 15712 37806
rect 15660 37742 15712 37748
rect 15672 37330 15700 37742
rect 15660 37324 15712 37330
rect 15660 37266 15712 37272
rect 16132 36922 16160 38286
rect 16868 37466 16896 38286
rect 16856 37460 16908 37466
rect 16856 37402 16908 37408
rect 16960 37126 16988 40530
rect 17052 40458 17080 41074
rect 17328 40594 17356 41074
rect 17512 41070 17540 41754
rect 17500 41064 17552 41070
rect 17500 41006 17552 41012
rect 17316 40588 17368 40594
rect 17316 40530 17368 40536
rect 17040 40452 17092 40458
rect 17040 40394 17092 40400
rect 17500 38956 17552 38962
rect 17500 38898 17552 38904
rect 17132 38548 17184 38554
rect 17132 38490 17184 38496
rect 17144 38282 17172 38490
rect 17132 38276 17184 38282
rect 17132 38218 17184 38224
rect 16948 37120 17000 37126
rect 16948 37062 17000 37068
rect 16120 36916 16172 36922
rect 16120 36858 16172 36864
rect 17144 36786 17172 38218
rect 17512 38010 17540 38898
rect 17592 38276 17644 38282
rect 17592 38218 17644 38224
rect 17500 38004 17552 38010
rect 17500 37946 17552 37952
rect 17224 37800 17276 37806
rect 17224 37742 17276 37748
rect 17132 36780 17184 36786
rect 17132 36722 17184 36728
rect 16028 36712 16080 36718
rect 16028 36654 16080 36660
rect 16120 36712 16172 36718
rect 16120 36654 16172 36660
rect 16040 36378 16068 36654
rect 16028 36372 16080 36378
rect 16028 36314 16080 36320
rect 16132 36242 16160 36654
rect 16120 36236 16172 36242
rect 16120 36178 16172 36184
rect 16948 36236 17000 36242
rect 16948 36178 17000 36184
rect 15200 36168 15252 36174
rect 15200 36110 15252 36116
rect 14832 36032 14884 36038
rect 14832 35974 14884 35980
rect 15292 36032 15344 36038
rect 15292 35974 15344 35980
rect 14844 35834 14872 35974
rect 14832 35828 14884 35834
rect 14832 35770 14884 35776
rect 15304 35290 15332 35974
rect 15384 35760 15436 35766
rect 15384 35702 15436 35708
rect 15292 35284 15344 35290
rect 15292 35226 15344 35232
rect 15396 35222 15424 35702
rect 15660 35488 15712 35494
rect 15660 35430 15712 35436
rect 15384 35216 15436 35222
rect 15384 35158 15436 35164
rect 14556 35080 14608 35086
rect 14556 35022 14608 35028
rect 14740 35080 14792 35086
rect 14740 35022 14792 35028
rect 14568 34610 14596 35022
rect 14752 34610 14780 35022
rect 15016 34944 15068 34950
rect 15016 34886 15068 34892
rect 14556 34604 14608 34610
rect 14556 34546 14608 34552
rect 14740 34604 14792 34610
rect 14740 34546 14792 34552
rect 14752 33590 14780 34546
rect 15028 34406 15056 34886
rect 15200 34536 15252 34542
rect 15200 34478 15252 34484
rect 15016 34400 15068 34406
rect 15016 34342 15068 34348
rect 15028 33998 15056 34342
rect 15212 33998 15240 34478
rect 15396 33998 15424 35158
rect 15672 35154 15700 35430
rect 15660 35148 15712 35154
rect 15660 35090 15712 35096
rect 15844 35080 15896 35086
rect 15844 35022 15896 35028
rect 15856 34746 15884 35022
rect 15844 34740 15896 34746
rect 15844 34682 15896 34688
rect 15016 33992 15068 33998
rect 15016 33934 15068 33940
rect 15200 33992 15252 33998
rect 15200 33934 15252 33940
rect 15384 33992 15436 33998
rect 15384 33934 15436 33940
rect 15752 33856 15804 33862
rect 15752 33798 15804 33804
rect 14740 33584 14792 33590
rect 14740 33526 14792 33532
rect 14924 33516 14976 33522
rect 14924 33458 14976 33464
rect 14464 33312 14516 33318
rect 14464 33254 14516 33260
rect 14372 32972 14424 32978
rect 14372 32914 14424 32920
rect 14476 32910 14504 33254
rect 14936 33046 14964 33458
rect 15200 33380 15252 33386
rect 15200 33322 15252 33328
rect 14924 33040 14976 33046
rect 14924 32982 14976 32988
rect 14464 32904 14516 32910
rect 14464 32846 14516 32852
rect 14936 32434 14964 32982
rect 15016 32972 15068 32978
rect 15016 32914 15068 32920
rect 14924 32428 14976 32434
rect 14924 32370 14976 32376
rect 14096 31272 14148 31278
rect 14096 31214 14148 31220
rect 14464 31272 14516 31278
rect 14464 31214 14516 31220
rect 13636 31204 13688 31210
rect 13636 31146 13688 31152
rect 13544 31136 13596 31142
rect 13544 31078 13596 31084
rect 13556 30734 13584 31078
rect 13544 30728 13596 30734
rect 13544 30670 13596 30676
rect 13648 30666 13676 31146
rect 13728 30728 13780 30734
rect 13728 30670 13780 30676
rect 13636 30660 13688 30666
rect 13636 30602 13688 30608
rect 13084 30048 13136 30054
rect 13084 29990 13136 29996
rect 13096 29646 13124 29990
rect 12900 29640 12952 29646
rect 12900 29582 12952 29588
rect 13084 29640 13136 29646
rect 13084 29582 13136 29588
rect 12808 28076 12860 28082
rect 12808 28018 12860 28024
rect 12728 27934 12848 27962
rect 12716 27872 12768 27878
rect 12716 27814 12768 27820
rect 12728 26994 12756 27814
rect 12716 26988 12768 26994
rect 12716 26930 12768 26936
rect 12820 25906 12848 27934
rect 12912 25974 12940 29582
rect 13648 28948 13676 30602
rect 13740 30054 13768 30670
rect 13728 30048 13780 30054
rect 13728 29990 13780 29996
rect 13648 28920 13952 28948
rect 13820 28756 13872 28762
rect 13820 28698 13872 28704
rect 13452 28552 13504 28558
rect 13452 28494 13504 28500
rect 13636 28552 13688 28558
rect 13636 28494 13688 28500
rect 13464 28218 13492 28494
rect 13544 28416 13596 28422
rect 13544 28358 13596 28364
rect 13452 28212 13504 28218
rect 13452 28154 13504 28160
rect 12992 28076 13044 28082
rect 12992 28018 13044 28024
rect 12900 25968 12952 25974
rect 12900 25910 12952 25916
rect 12808 25900 12860 25906
rect 12808 25842 12860 25848
rect 12808 24744 12860 24750
rect 12808 24686 12860 24692
rect 12820 24138 12848 24686
rect 12808 24132 12860 24138
rect 12808 24074 12860 24080
rect 13004 23322 13032 28018
rect 13464 27334 13492 28154
rect 13556 27334 13584 28358
rect 13452 27328 13504 27334
rect 13452 27270 13504 27276
rect 13544 27328 13596 27334
rect 13544 27270 13596 27276
rect 13464 26382 13492 27270
rect 13556 26994 13584 27270
rect 13544 26988 13596 26994
rect 13544 26930 13596 26936
rect 13648 26382 13676 28494
rect 13832 28014 13860 28698
rect 13820 28008 13872 28014
rect 13820 27950 13872 27956
rect 13452 26376 13504 26382
rect 13452 26318 13504 26324
rect 13636 26376 13688 26382
rect 13636 26318 13688 26324
rect 13648 25906 13676 26318
rect 13636 25900 13688 25906
rect 13636 25842 13688 25848
rect 13648 25498 13676 25842
rect 13636 25492 13688 25498
rect 13636 25434 13688 25440
rect 13820 25288 13872 25294
rect 13820 25230 13872 25236
rect 13832 24818 13860 25230
rect 13820 24812 13872 24818
rect 13820 24754 13872 24760
rect 13360 23520 13412 23526
rect 13360 23462 13412 23468
rect 12992 23316 13044 23322
rect 12992 23258 13044 23264
rect 13176 22432 13228 22438
rect 13176 22374 13228 22380
rect 13188 22030 13216 22374
rect 13268 22092 13320 22098
rect 13268 22034 13320 22040
rect 12808 22024 12860 22030
rect 12808 21966 12860 21972
rect 13176 22024 13228 22030
rect 13176 21966 13228 21972
rect 12820 21146 12848 21966
rect 13188 21622 13216 21966
rect 13280 21690 13308 22034
rect 13268 21684 13320 21690
rect 13268 21626 13320 21632
rect 13176 21616 13228 21622
rect 13176 21558 13228 21564
rect 12808 21140 12860 21146
rect 12808 21082 12860 21088
rect 13280 21010 13308 21626
rect 13372 21486 13400 23462
rect 13924 23186 13952 28920
rect 14476 28762 14504 31214
rect 14464 28756 14516 28762
rect 14464 28698 14516 28704
rect 14556 28620 14608 28626
rect 14556 28562 14608 28568
rect 14568 28150 14596 28562
rect 14832 28484 14884 28490
rect 14832 28426 14884 28432
rect 14556 28144 14608 28150
rect 14556 28086 14608 28092
rect 14372 28076 14424 28082
rect 14372 28018 14424 28024
rect 14384 27606 14412 28018
rect 14568 27962 14596 28086
rect 14844 28082 14872 28426
rect 14832 28076 14884 28082
rect 14832 28018 14884 28024
rect 14568 27934 14688 27962
rect 14556 27872 14608 27878
rect 14556 27814 14608 27820
rect 14372 27600 14424 27606
rect 14372 27542 14424 27548
rect 14568 27470 14596 27814
rect 14556 27464 14608 27470
rect 14556 27406 14608 27412
rect 14660 27130 14688 27934
rect 14648 27124 14700 27130
rect 14648 27066 14700 27072
rect 14188 26920 14240 26926
rect 14188 26862 14240 26868
rect 14200 26586 14228 26862
rect 14188 26580 14240 26586
rect 14188 26522 14240 26528
rect 14832 26240 14884 26246
rect 14832 26182 14884 26188
rect 14844 25294 14872 26182
rect 14832 25288 14884 25294
rect 14832 25230 14884 25236
rect 14372 24812 14424 24818
rect 14372 24754 14424 24760
rect 14384 24410 14412 24754
rect 14372 24404 14424 24410
rect 14372 24346 14424 24352
rect 13912 23180 13964 23186
rect 13912 23122 13964 23128
rect 14556 23112 14608 23118
rect 14556 23054 14608 23060
rect 14568 22710 14596 23054
rect 14556 22704 14608 22710
rect 14556 22646 14608 22652
rect 14280 22636 14332 22642
rect 14280 22578 14332 22584
rect 14292 22234 14320 22578
rect 14280 22228 14332 22234
rect 14280 22170 14332 22176
rect 14924 22160 14976 22166
rect 14924 22102 14976 22108
rect 13912 22024 13964 22030
rect 13912 21966 13964 21972
rect 13924 21690 13952 21966
rect 13912 21684 13964 21690
rect 13912 21626 13964 21632
rect 13360 21480 13412 21486
rect 13360 21422 13412 21428
rect 13372 21010 13400 21422
rect 13820 21344 13872 21350
rect 13820 21286 13872 21292
rect 13268 21004 13320 21010
rect 13268 20946 13320 20952
rect 13360 21004 13412 21010
rect 13360 20946 13412 20952
rect 13176 20800 13228 20806
rect 13176 20742 13228 20748
rect 13188 20534 13216 20742
rect 13176 20528 13228 20534
rect 13176 20470 13228 20476
rect 12716 18828 12768 18834
rect 12716 18770 12768 18776
rect 12728 18222 12756 18770
rect 13372 18222 13400 20946
rect 13832 20466 13860 21286
rect 13820 20460 13872 20466
rect 13820 20402 13872 20408
rect 14936 19378 14964 22102
rect 13912 19372 13964 19378
rect 13912 19314 13964 19320
rect 14924 19372 14976 19378
rect 14924 19314 14976 19320
rect 13924 18902 13952 19314
rect 15028 19310 15056 32914
rect 15212 32570 15240 33322
rect 15200 32564 15252 32570
rect 15200 32506 15252 32512
rect 15384 32224 15436 32230
rect 15384 32166 15436 32172
rect 15396 31482 15424 32166
rect 15384 31476 15436 31482
rect 15384 31418 15436 31424
rect 15568 31272 15620 31278
rect 15568 31214 15620 31220
rect 15580 30938 15608 31214
rect 15568 30932 15620 30938
rect 15568 30874 15620 30880
rect 15476 30728 15528 30734
rect 15476 30670 15528 30676
rect 15200 30592 15252 30598
rect 15200 30534 15252 30540
rect 15212 30258 15240 30534
rect 15488 30258 15516 30670
rect 15200 30252 15252 30258
rect 15200 30194 15252 30200
rect 15476 30252 15528 30258
rect 15476 30194 15528 30200
rect 15764 30138 15792 33798
rect 16132 32366 16160 36178
rect 16304 36168 16356 36174
rect 16304 36110 16356 36116
rect 16316 35630 16344 36110
rect 16960 35834 16988 36178
rect 16948 35828 17000 35834
rect 16948 35770 17000 35776
rect 16304 35624 16356 35630
rect 16304 35566 16356 35572
rect 16960 35290 16988 35770
rect 16948 35284 17000 35290
rect 16948 35226 17000 35232
rect 16672 34944 16724 34950
rect 16672 34886 16724 34892
rect 15844 32360 15896 32366
rect 15844 32302 15896 32308
rect 16120 32360 16172 32366
rect 16120 32302 16172 32308
rect 15856 31278 15884 32302
rect 15844 31272 15896 31278
rect 15844 31214 15896 31220
rect 15936 30864 15988 30870
rect 15936 30806 15988 30812
rect 15764 30110 15884 30138
rect 15752 30048 15804 30054
rect 15752 29990 15804 29996
rect 15764 29850 15792 29990
rect 15752 29844 15804 29850
rect 15752 29786 15804 29792
rect 15384 29164 15436 29170
rect 15384 29106 15436 29112
rect 15200 28416 15252 28422
rect 15200 28358 15252 28364
rect 15212 27402 15240 28358
rect 15396 27606 15424 29106
rect 15856 28558 15884 30110
rect 15948 30054 15976 30806
rect 15936 30048 15988 30054
rect 15936 29990 15988 29996
rect 15936 29640 15988 29646
rect 15936 29582 15988 29588
rect 16028 29640 16080 29646
rect 16028 29582 16080 29588
rect 15948 29170 15976 29582
rect 16040 29170 16068 29582
rect 15936 29164 15988 29170
rect 15936 29106 15988 29112
rect 16028 29164 16080 29170
rect 16028 29106 16080 29112
rect 15752 28552 15804 28558
rect 15752 28494 15804 28500
rect 15844 28552 15896 28558
rect 15844 28494 15896 28500
rect 15476 28144 15528 28150
rect 15476 28086 15528 28092
rect 15384 27600 15436 27606
rect 15384 27542 15436 27548
rect 15292 27464 15344 27470
rect 15292 27406 15344 27412
rect 15200 27396 15252 27402
rect 15200 27338 15252 27344
rect 15304 24682 15332 27406
rect 15488 27334 15516 28086
rect 15764 27946 15792 28494
rect 15856 28014 15884 28494
rect 16040 28218 16068 29106
rect 16028 28212 16080 28218
rect 16028 28154 16080 28160
rect 15844 28008 15896 28014
rect 15844 27950 15896 27956
rect 15752 27940 15804 27946
rect 15752 27882 15804 27888
rect 15568 27872 15620 27878
rect 15568 27814 15620 27820
rect 15580 27470 15608 27814
rect 15568 27464 15620 27470
rect 15568 27406 15620 27412
rect 15660 27464 15712 27470
rect 15660 27406 15712 27412
rect 15476 27328 15528 27334
rect 15476 27270 15528 27276
rect 15580 26926 15608 27406
rect 15672 27130 15700 27406
rect 15764 27334 15792 27882
rect 16132 27606 16160 32302
rect 16488 31816 16540 31822
rect 16488 31758 16540 31764
rect 16500 31142 16528 31758
rect 16580 31272 16632 31278
rect 16580 31214 16632 31220
rect 16488 31136 16540 31142
rect 16488 31078 16540 31084
rect 16304 30864 16356 30870
rect 16304 30806 16356 30812
rect 16316 30598 16344 30806
rect 16500 30734 16528 31078
rect 16592 30870 16620 31214
rect 16580 30864 16632 30870
rect 16580 30806 16632 30812
rect 16488 30728 16540 30734
rect 16488 30670 16540 30676
rect 16304 30592 16356 30598
rect 16304 30534 16356 30540
rect 16684 29510 16712 34886
rect 16856 33924 16908 33930
rect 16856 33866 16908 33872
rect 16868 33658 16896 33866
rect 17132 33856 17184 33862
rect 17132 33798 17184 33804
rect 16856 33652 16908 33658
rect 16856 33594 16908 33600
rect 17040 33516 17092 33522
rect 17040 33458 17092 33464
rect 17052 33114 17080 33458
rect 17040 33108 17092 33114
rect 17040 33050 17092 33056
rect 17144 32910 17172 33798
rect 17236 33522 17264 37742
rect 17500 33992 17552 33998
rect 17500 33934 17552 33940
rect 17512 33590 17540 33934
rect 17500 33584 17552 33590
rect 17500 33526 17552 33532
rect 17224 33516 17276 33522
rect 17224 33458 17276 33464
rect 16856 32904 16908 32910
rect 16856 32846 16908 32852
rect 17132 32904 17184 32910
rect 17132 32846 17184 32852
rect 16868 32366 16896 32846
rect 17144 32570 17172 32846
rect 17132 32564 17184 32570
rect 17132 32506 17184 32512
rect 16856 32360 16908 32366
rect 16856 32302 16908 32308
rect 17132 31884 17184 31890
rect 17132 31826 17184 31832
rect 16764 31680 16816 31686
rect 16764 31622 16816 31628
rect 16776 30870 16804 31622
rect 16856 31340 16908 31346
rect 16856 31282 16908 31288
rect 17040 31340 17092 31346
rect 17040 31282 17092 31288
rect 16764 30864 16816 30870
rect 16764 30806 16816 30812
rect 16776 30122 16804 30806
rect 16868 30258 16896 31282
rect 16948 30728 17000 30734
rect 16948 30670 17000 30676
rect 16960 30394 16988 30670
rect 16948 30388 17000 30394
rect 16948 30330 17000 30336
rect 16856 30252 16908 30258
rect 16856 30194 16908 30200
rect 16764 30116 16816 30122
rect 16764 30058 16816 30064
rect 16672 29504 16724 29510
rect 16672 29446 16724 29452
rect 16580 29300 16632 29306
rect 16580 29242 16632 29248
rect 16592 28558 16620 29242
rect 16684 29238 16712 29446
rect 16672 29232 16724 29238
rect 16672 29174 16724 29180
rect 16580 28552 16632 28558
rect 16580 28494 16632 28500
rect 16212 28416 16264 28422
rect 16212 28358 16264 28364
rect 16224 27878 16252 28358
rect 16212 27872 16264 27878
rect 16212 27814 16264 27820
rect 16592 27606 16620 28494
rect 16684 28422 16712 29174
rect 16960 29102 16988 30330
rect 17052 30326 17080 31282
rect 17144 30326 17172 31826
rect 17040 30320 17092 30326
rect 17040 30262 17092 30268
rect 17132 30320 17184 30326
rect 17132 30262 17184 30268
rect 16948 29096 17000 29102
rect 16948 29038 17000 29044
rect 16948 28960 17000 28966
rect 16948 28902 17000 28908
rect 16960 28558 16988 28902
rect 16948 28552 17000 28558
rect 16948 28494 17000 28500
rect 16672 28416 16724 28422
rect 16672 28358 16724 28364
rect 16120 27600 16172 27606
rect 16120 27542 16172 27548
rect 16580 27600 16632 27606
rect 16580 27542 16632 27548
rect 16856 27532 16908 27538
rect 16856 27474 16908 27480
rect 16580 27464 16632 27470
rect 16580 27406 16632 27412
rect 15752 27328 15804 27334
rect 15752 27270 15804 27276
rect 15660 27124 15712 27130
rect 15660 27066 15712 27072
rect 16592 26994 16620 27406
rect 16868 27130 16896 27474
rect 16856 27124 16908 27130
rect 16856 27066 16908 27072
rect 16580 26988 16632 26994
rect 16580 26930 16632 26936
rect 15568 26920 15620 26926
rect 15568 26862 15620 26868
rect 17052 25906 17080 30262
rect 17236 29050 17264 33458
rect 17316 33448 17368 33454
rect 17316 33390 17368 33396
rect 17328 31414 17356 33390
rect 17512 32978 17540 33526
rect 17500 32972 17552 32978
rect 17500 32914 17552 32920
rect 17604 32366 17632 38218
rect 17684 38208 17736 38214
rect 17684 38150 17736 38156
rect 17696 37874 17724 38150
rect 17972 37874 18000 47126
rect 19352 47054 19380 49200
rect 19340 47048 19392 47054
rect 22468 47048 22520 47054
rect 19340 46990 19392 46996
rect 19706 47016 19762 47025
rect 22468 46990 22520 46996
rect 19706 46951 19708 46960
rect 19760 46951 19762 46960
rect 19708 46922 19760 46928
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 22480 46578 22508 46990
rect 22468 46572 22520 46578
rect 22468 46514 22520 46520
rect 23216 46510 23244 49200
rect 23860 47054 23888 49200
rect 23848 47048 23900 47054
rect 23848 46990 23900 46996
rect 22744 46504 22796 46510
rect 22744 46446 22796 46452
rect 23204 46504 23256 46510
rect 23204 46446 23256 46452
rect 24952 46504 25004 46510
rect 24952 46446 25004 46452
rect 22756 46170 22784 46446
rect 22744 46164 22796 46170
rect 22744 46106 22796 46112
rect 19064 46028 19116 46034
rect 19064 45970 19116 45976
rect 19076 43382 19104 45970
rect 22652 45960 22704 45966
rect 22652 45902 22704 45908
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 22664 45626 22692 45902
rect 24860 45892 24912 45898
rect 24860 45834 24912 45840
rect 24872 45626 24900 45834
rect 24964 45626 24992 46446
rect 25148 45898 25176 49200
rect 25688 47048 25740 47054
rect 25688 46990 25740 46996
rect 25412 46980 25464 46986
rect 25412 46922 25464 46928
rect 25136 45892 25188 45898
rect 25136 45834 25188 45840
rect 22652 45620 22704 45626
rect 22652 45562 22704 45568
rect 24860 45620 24912 45626
rect 24860 45562 24912 45568
rect 24952 45620 25004 45626
rect 24952 45562 25004 45568
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 20536 44192 20588 44198
rect 20536 44134 20588 44140
rect 20548 43858 20576 44134
rect 20536 43852 20588 43858
rect 20536 43794 20588 43800
rect 20352 43784 20404 43790
rect 20352 43726 20404 43732
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 19064 43376 19116 43382
rect 19064 43318 19116 43324
rect 19524 42696 19576 42702
rect 19444 42644 19524 42650
rect 19444 42638 19576 42644
rect 19444 42622 19564 42638
rect 20364 42634 20392 43726
rect 22560 42764 22612 42770
rect 22560 42706 22612 42712
rect 20628 42696 20680 42702
rect 20628 42638 20680 42644
rect 20352 42628 20404 42634
rect 19340 42560 19392 42566
rect 19340 42502 19392 42508
rect 19352 41682 19380 42502
rect 19444 42362 19472 42622
rect 20352 42570 20404 42576
rect 20168 42560 20220 42566
rect 20168 42502 20220 42508
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 19432 42356 19484 42362
rect 19432 42298 19484 42304
rect 19984 42356 20036 42362
rect 19984 42298 20036 42304
rect 19432 42220 19484 42226
rect 19432 42162 19484 42168
rect 19444 41818 19472 42162
rect 19432 41812 19484 41818
rect 19432 41754 19484 41760
rect 19340 41676 19392 41682
rect 19340 41618 19392 41624
rect 19432 41472 19484 41478
rect 19432 41414 19484 41420
rect 19248 41064 19300 41070
rect 19248 41006 19300 41012
rect 18420 39976 18472 39982
rect 18420 39918 18472 39924
rect 18432 39506 18460 39918
rect 18420 39500 18472 39506
rect 18420 39442 18472 39448
rect 18432 39030 18460 39442
rect 18420 39024 18472 39030
rect 18420 38966 18472 38972
rect 18420 38752 18472 38758
rect 18420 38694 18472 38700
rect 18432 38350 18460 38694
rect 18420 38344 18472 38350
rect 18420 38286 18472 38292
rect 17684 37868 17736 37874
rect 17684 37810 17736 37816
rect 17960 37868 18012 37874
rect 17960 37810 18012 37816
rect 17868 37256 17920 37262
rect 17788 37216 17868 37244
rect 17788 37126 17816 37216
rect 17868 37198 17920 37204
rect 17776 37120 17828 37126
rect 17776 37062 17828 37068
rect 17684 35692 17736 35698
rect 17684 35634 17736 35640
rect 17696 35222 17724 35634
rect 17684 35216 17736 35222
rect 17684 35158 17736 35164
rect 17592 32360 17644 32366
rect 17592 32302 17644 32308
rect 17316 31408 17368 31414
rect 17316 31350 17368 31356
rect 17592 31340 17644 31346
rect 17592 31282 17644 31288
rect 17604 30870 17632 31282
rect 17592 30864 17644 30870
rect 17592 30806 17644 30812
rect 17684 30728 17736 30734
rect 17684 30670 17736 30676
rect 17696 30258 17724 30670
rect 17684 30252 17736 30258
rect 17684 30194 17736 30200
rect 17696 30122 17724 30194
rect 17684 30116 17736 30122
rect 17684 30058 17736 30064
rect 17236 29022 17356 29050
rect 17224 28960 17276 28966
rect 17224 28902 17276 28908
rect 17236 28082 17264 28902
rect 17224 28076 17276 28082
rect 17224 28018 17276 28024
rect 17224 27396 17276 27402
rect 17224 27338 17276 27344
rect 17236 26994 17264 27338
rect 17224 26988 17276 26994
rect 17224 26930 17276 26936
rect 17236 26586 17264 26930
rect 17224 26580 17276 26586
rect 17224 26522 17276 26528
rect 16580 25900 16632 25906
rect 16580 25842 16632 25848
rect 17040 25900 17092 25906
rect 17040 25842 17092 25848
rect 16592 25498 16620 25842
rect 16856 25696 16908 25702
rect 16856 25638 16908 25644
rect 17040 25696 17092 25702
rect 17040 25638 17092 25644
rect 16580 25492 16632 25498
rect 16580 25434 16632 25440
rect 16868 25294 16896 25638
rect 17052 25294 17080 25638
rect 17328 25498 17356 29022
rect 17408 28552 17460 28558
rect 17408 28494 17460 28500
rect 17420 28014 17448 28494
rect 17500 28416 17552 28422
rect 17500 28358 17552 28364
rect 17408 28008 17460 28014
rect 17408 27950 17460 27956
rect 17420 26382 17448 27950
rect 17512 27470 17540 28358
rect 17500 27464 17552 27470
rect 17500 27406 17552 27412
rect 17408 26376 17460 26382
rect 17408 26318 17460 26324
rect 17316 25492 17368 25498
rect 17316 25434 17368 25440
rect 16856 25288 16908 25294
rect 16856 25230 16908 25236
rect 17040 25288 17092 25294
rect 17040 25230 17092 25236
rect 15844 24812 15896 24818
rect 15844 24754 15896 24760
rect 15292 24676 15344 24682
rect 15292 24618 15344 24624
rect 15660 24608 15712 24614
rect 15660 24550 15712 24556
rect 15672 24274 15700 24550
rect 15856 24410 15884 24754
rect 17052 24682 17080 25230
rect 17040 24676 17092 24682
rect 17040 24618 17092 24624
rect 15844 24404 15896 24410
rect 15844 24346 15896 24352
rect 17328 24342 17356 25434
rect 17592 25288 17644 25294
rect 17592 25230 17644 25236
rect 17604 24954 17632 25230
rect 17592 24948 17644 24954
rect 17592 24890 17644 24896
rect 17316 24336 17368 24342
rect 17316 24278 17368 24284
rect 15660 24268 15712 24274
rect 15660 24210 15712 24216
rect 17500 24200 17552 24206
rect 17500 24142 17552 24148
rect 17408 24132 17460 24138
rect 17408 24074 17460 24080
rect 16948 24064 17000 24070
rect 16948 24006 17000 24012
rect 16856 23792 16908 23798
rect 16856 23734 16908 23740
rect 16868 22710 16896 23734
rect 16960 23050 16988 24006
rect 16948 23044 17000 23050
rect 16948 22986 17000 22992
rect 17316 22976 17368 22982
rect 17316 22918 17368 22924
rect 16856 22704 16908 22710
rect 16856 22646 16908 22652
rect 15568 22432 15620 22438
rect 15568 22374 15620 22380
rect 15580 22098 15608 22374
rect 15568 22092 15620 22098
rect 15568 22034 15620 22040
rect 15844 22092 15896 22098
rect 15844 22034 15896 22040
rect 15856 21486 15884 22034
rect 17328 22030 17356 22918
rect 17316 22024 17368 22030
rect 17316 21966 17368 21972
rect 15936 21888 15988 21894
rect 15936 21830 15988 21836
rect 15844 21480 15896 21486
rect 15844 21422 15896 21428
rect 15200 20868 15252 20874
rect 15200 20810 15252 20816
rect 15212 20058 15240 20810
rect 15856 20398 15884 21422
rect 15292 20392 15344 20398
rect 15292 20334 15344 20340
rect 15844 20392 15896 20398
rect 15844 20334 15896 20340
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 14096 19304 14148 19310
rect 14096 19246 14148 19252
rect 15016 19304 15068 19310
rect 15304 19258 15332 20334
rect 15384 20256 15436 20262
rect 15384 20198 15436 20204
rect 15396 19854 15424 20198
rect 15384 19848 15436 19854
rect 15384 19790 15436 19796
rect 15476 19712 15528 19718
rect 15476 19654 15528 19660
rect 15016 19246 15068 19252
rect 13912 18896 13964 18902
rect 13912 18838 13964 18844
rect 13912 18760 13964 18766
rect 13912 18702 13964 18708
rect 12716 18216 12768 18222
rect 12716 18158 12768 18164
rect 13360 18216 13412 18222
rect 13360 18158 13412 18164
rect 12624 18148 12676 18154
rect 12624 18090 12676 18096
rect 12728 17882 12756 18158
rect 12716 17876 12768 17882
rect 12716 17818 12768 17824
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 12728 16794 12756 17138
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 13188 16658 13216 17138
rect 13372 16658 13400 18158
rect 13924 17270 13952 18702
rect 13912 17264 13964 17270
rect 13912 17206 13964 17212
rect 13176 16652 13228 16658
rect 13176 16594 13228 16600
rect 13360 16652 13412 16658
rect 13360 16594 13412 16600
rect 13188 16250 13216 16594
rect 13176 16244 13228 16250
rect 13176 16186 13228 16192
rect 12164 16108 12216 16114
rect 12164 16050 12216 16056
rect 12900 16108 12952 16114
rect 12900 16050 12952 16056
rect 12912 15706 12940 16050
rect 13372 16046 13400 16594
rect 13360 16040 13412 16046
rect 13360 15982 13412 15988
rect 13084 15904 13136 15910
rect 13084 15846 13136 15852
rect 12900 15700 12952 15706
rect 12900 15642 12952 15648
rect 13096 15502 13124 15846
rect 13084 15496 13136 15502
rect 13084 15438 13136 15444
rect 13924 15026 13952 17206
rect 14108 17134 14136 19246
rect 15212 19230 15332 19258
rect 15212 19174 15240 19230
rect 15200 19168 15252 19174
rect 15200 19110 15252 19116
rect 15488 18766 15516 19654
rect 15476 18760 15528 18766
rect 15476 18702 15528 18708
rect 15856 18154 15884 20334
rect 15948 19854 15976 21830
rect 16028 21480 16080 21486
rect 16028 21422 16080 21428
rect 16040 21146 16068 21422
rect 16028 21140 16080 21146
rect 16028 21082 16080 21088
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 16396 18692 16448 18698
rect 16396 18634 16448 18640
rect 16028 18624 16080 18630
rect 16028 18566 16080 18572
rect 16040 18222 16068 18566
rect 16408 18426 16436 18634
rect 16396 18420 16448 18426
rect 16396 18362 16448 18368
rect 16028 18216 16080 18222
rect 16028 18158 16080 18164
rect 15844 18148 15896 18154
rect 15844 18090 15896 18096
rect 15200 18080 15252 18086
rect 15200 18022 15252 18028
rect 15212 17678 15240 18022
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 15016 17536 15068 17542
rect 15016 17478 15068 17484
rect 15028 17270 15056 17478
rect 15016 17264 15068 17270
rect 15016 17206 15068 17212
rect 14096 17128 14148 17134
rect 14096 17070 14148 17076
rect 15016 16992 15068 16998
rect 15016 16934 15068 16940
rect 15028 15570 15056 16934
rect 16776 16794 16804 18702
rect 16856 16992 16908 16998
rect 16856 16934 16908 16940
rect 16764 16788 16816 16794
rect 16764 16730 16816 16736
rect 15200 16108 15252 16114
rect 15200 16050 15252 16056
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 15120 15570 15148 15982
rect 15016 15564 15068 15570
rect 15016 15506 15068 15512
rect 15108 15564 15160 15570
rect 15108 15506 15160 15512
rect 14096 15360 14148 15366
rect 14096 15302 14148 15308
rect 14108 15094 14136 15302
rect 15212 15162 15240 16050
rect 15200 15156 15252 15162
rect 15200 15098 15252 15104
rect 14096 15088 14148 15094
rect 14096 15030 14148 15036
rect 16776 15026 16804 16730
rect 16868 16522 16896 16934
rect 16856 16516 16908 16522
rect 16856 16458 16908 16464
rect 17040 16176 17092 16182
rect 17040 16118 17092 16124
rect 17052 15502 17080 16118
rect 17420 15586 17448 24074
rect 17512 23866 17540 24142
rect 17500 23860 17552 23866
rect 17500 23802 17552 23808
rect 17500 16448 17552 16454
rect 17500 16390 17552 16396
rect 17512 16250 17540 16390
rect 17500 16244 17552 16250
rect 17500 16186 17552 16192
rect 17604 16046 17632 24890
rect 17788 22094 17816 37062
rect 17868 35692 17920 35698
rect 17868 35634 17920 35640
rect 17880 34950 17908 35634
rect 17868 34944 17920 34950
rect 17868 34886 17920 34892
rect 17972 33454 18000 37810
rect 18328 36848 18380 36854
rect 18328 36790 18380 36796
rect 18340 36242 18368 36790
rect 18432 36786 18460 38286
rect 19260 38214 19288 41006
rect 19444 40526 19472 41414
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 19996 41138 20024 42298
rect 20180 41750 20208 42502
rect 20364 42362 20392 42570
rect 20352 42356 20404 42362
rect 20352 42298 20404 42304
rect 20168 41744 20220 41750
rect 20168 41686 20220 41692
rect 20076 41676 20128 41682
rect 20076 41618 20128 41624
rect 20088 41206 20116 41618
rect 20180 41274 20208 41686
rect 20364 41682 20392 42298
rect 20640 42090 20668 42638
rect 22100 42220 22152 42226
rect 22100 42162 22152 42168
rect 20628 42084 20680 42090
rect 20628 42026 20680 42032
rect 20352 41676 20404 41682
rect 20352 41618 20404 41624
rect 20260 41608 20312 41614
rect 20260 41550 20312 41556
rect 20536 41608 20588 41614
rect 20536 41550 20588 41556
rect 20168 41268 20220 41274
rect 20168 41210 20220 41216
rect 20076 41200 20128 41206
rect 20076 41142 20128 41148
rect 19984 41132 20036 41138
rect 19984 41074 20036 41080
rect 20076 40928 20128 40934
rect 20076 40870 20128 40876
rect 20088 40594 20116 40870
rect 20076 40588 20128 40594
rect 20076 40530 20128 40536
rect 19432 40520 19484 40526
rect 19432 40462 19484 40468
rect 19432 40384 19484 40390
rect 19432 40326 19484 40332
rect 19984 40384 20036 40390
rect 19984 40326 20036 40332
rect 19444 40050 19472 40326
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 19432 40044 19484 40050
rect 19432 39986 19484 39992
rect 19432 39364 19484 39370
rect 19432 39306 19484 39312
rect 19248 38208 19300 38214
rect 19248 38150 19300 38156
rect 18696 37868 18748 37874
rect 18696 37810 18748 37816
rect 18708 37262 18736 37810
rect 18696 37256 18748 37262
rect 18696 37198 18748 37204
rect 18420 36780 18472 36786
rect 18420 36722 18472 36728
rect 18328 36236 18380 36242
rect 18328 36178 18380 36184
rect 18708 34542 18736 37198
rect 19260 35698 19288 38150
rect 19340 37256 19392 37262
rect 19340 37198 19392 37204
rect 19352 36666 19380 37198
rect 19444 37194 19472 39306
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 19996 39098 20024 40326
rect 19984 39092 20036 39098
rect 19984 39034 20036 39040
rect 19616 38956 19668 38962
rect 19616 38898 19668 38904
rect 19984 38956 20036 38962
rect 19984 38898 20036 38904
rect 19628 38554 19656 38898
rect 19616 38548 19668 38554
rect 19616 38490 19668 38496
rect 19996 38282 20024 38898
rect 19984 38276 20036 38282
rect 19984 38218 20036 38224
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 19996 37466 20024 38218
rect 20272 38010 20300 41550
rect 20548 41206 20576 41550
rect 20536 41200 20588 41206
rect 20536 41142 20588 41148
rect 20352 41132 20404 41138
rect 20352 41074 20404 41080
rect 20364 40186 20392 41074
rect 20444 40928 20496 40934
rect 20444 40870 20496 40876
rect 20456 40526 20484 40870
rect 20640 40526 20668 42026
rect 20996 42016 21048 42022
rect 20996 41958 21048 41964
rect 21008 41682 21036 41958
rect 22112 41682 22140 42162
rect 22572 42158 22600 42706
rect 22836 42696 22888 42702
rect 22836 42638 22888 42644
rect 23112 42696 23164 42702
rect 23112 42638 23164 42644
rect 22848 42362 22876 42638
rect 23020 42628 23072 42634
rect 23020 42570 23072 42576
rect 22836 42356 22888 42362
rect 22836 42298 22888 42304
rect 22560 42152 22612 42158
rect 22560 42094 22612 42100
rect 22572 41818 22600 42094
rect 22560 41812 22612 41818
rect 22560 41754 22612 41760
rect 20996 41676 21048 41682
rect 20996 41618 21048 41624
rect 22100 41676 22152 41682
rect 22100 41618 22152 41624
rect 21008 41414 21036 41618
rect 21824 41608 21876 41614
rect 21824 41550 21876 41556
rect 21008 41386 21128 41414
rect 20444 40520 20496 40526
rect 20444 40462 20496 40468
rect 20628 40520 20680 40526
rect 20628 40462 20680 40468
rect 20352 40180 20404 40186
rect 20352 40122 20404 40128
rect 20456 38894 20484 40462
rect 20536 40452 20588 40458
rect 20536 40394 20588 40400
rect 20548 38962 20576 40394
rect 20640 39506 20668 40462
rect 20628 39500 20680 39506
rect 20628 39442 20680 39448
rect 20536 38956 20588 38962
rect 20536 38898 20588 38904
rect 20444 38888 20496 38894
rect 20444 38830 20496 38836
rect 20260 38004 20312 38010
rect 20260 37946 20312 37952
rect 20168 37868 20220 37874
rect 20168 37810 20220 37816
rect 20076 37800 20128 37806
rect 20076 37742 20128 37748
rect 19984 37460 20036 37466
rect 19984 37402 20036 37408
rect 20088 37262 20116 37742
rect 20076 37256 20128 37262
rect 20076 37198 20128 37204
rect 19432 37188 19484 37194
rect 19432 37130 19484 37136
rect 19444 36825 19472 37130
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 20074 36952 20130 36961
rect 20074 36887 20130 36896
rect 20088 36854 20116 36887
rect 20076 36848 20128 36854
rect 19430 36816 19486 36825
rect 20076 36790 20128 36796
rect 19430 36751 19486 36760
rect 19892 36780 19944 36786
rect 19892 36722 19944 36728
rect 19984 36780 20036 36786
rect 19984 36722 20036 36728
rect 19904 36689 19932 36722
rect 19890 36680 19946 36689
rect 19352 36638 19472 36666
rect 19444 36582 19472 36638
rect 19890 36615 19946 36624
rect 19432 36576 19484 36582
rect 19432 36518 19484 36524
rect 19708 36576 19760 36582
rect 19708 36518 19760 36524
rect 19340 36032 19392 36038
rect 19340 35974 19392 35980
rect 19352 35766 19380 35974
rect 19340 35760 19392 35766
rect 19340 35702 19392 35708
rect 19064 35692 19116 35698
rect 19064 35634 19116 35640
rect 19248 35692 19300 35698
rect 19248 35634 19300 35640
rect 18880 35624 18932 35630
rect 18880 35566 18932 35572
rect 18892 35086 18920 35566
rect 19076 35222 19104 35634
rect 19064 35216 19116 35222
rect 19064 35158 19116 35164
rect 18880 35080 18932 35086
rect 18880 35022 18932 35028
rect 18696 34536 18748 34542
rect 18696 34478 18748 34484
rect 18236 33516 18288 33522
rect 18236 33458 18288 33464
rect 17960 33448 18012 33454
rect 17960 33390 18012 33396
rect 18052 33312 18104 33318
rect 18052 33254 18104 33260
rect 18064 32910 18092 33254
rect 18052 32904 18104 32910
rect 18052 32846 18104 32852
rect 18248 32570 18276 33458
rect 18604 33380 18656 33386
rect 18604 33322 18656 33328
rect 18328 33312 18380 33318
rect 18328 33254 18380 33260
rect 18340 32774 18368 33254
rect 18512 32904 18564 32910
rect 18512 32846 18564 32852
rect 18328 32768 18380 32774
rect 18328 32710 18380 32716
rect 18236 32564 18288 32570
rect 18236 32506 18288 32512
rect 18340 31754 18368 32710
rect 18524 32434 18552 32846
rect 18616 32502 18644 33322
rect 18892 32774 18920 35022
rect 19064 33448 19116 33454
rect 19064 33390 19116 33396
rect 18880 32768 18932 32774
rect 18880 32710 18932 32716
rect 18604 32496 18656 32502
rect 18604 32438 18656 32444
rect 18892 32434 18920 32710
rect 18512 32428 18564 32434
rect 18512 32370 18564 32376
rect 18880 32428 18932 32434
rect 18880 32370 18932 32376
rect 19076 31754 19104 33390
rect 18248 31726 18368 31754
rect 18984 31726 19104 31754
rect 17960 30932 18012 30938
rect 17960 30874 18012 30880
rect 17868 30660 17920 30666
rect 17868 30602 17920 30608
rect 17880 30394 17908 30602
rect 17868 30388 17920 30394
rect 17868 30330 17920 30336
rect 17880 30258 17908 30330
rect 17868 30252 17920 30258
rect 17868 30194 17920 30200
rect 17972 28150 18000 30874
rect 18052 30592 18104 30598
rect 18052 30534 18104 30540
rect 18064 30326 18092 30534
rect 18052 30320 18104 30326
rect 18052 30262 18104 30268
rect 17960 28144 18012 28150
rect 17960 28086 18012 28092
rect 18052 26512 18104 26518
rect 18052 26454 18104 26460
rect 17868 26308 17920 26314
rect 17868 26250 17920 26256
rect 17880 26042 17908 26250
rect 17868 26036 17920 26042
rect 17868 25978 17920 25984
rect 18064 25906 18092 26454
rect 18052 25900 18104 25906
rect 18052 25842 18104 25848
rect 18248 25702 18276 31726
rect 18604 30592 18656 30598
rect 18604 30534 18656 30540
rect 18788 30592 18840 30598
rect 18788 30534 18840 30540
rect 18512 30320 18564 30326
rect 18512 30262 18564 30268
rect 18524 29170 18552 30262
rect 18616 30258 18644 30534
rect 18800 30258 18828 30534
rect 18604 30252 18656 30258
rect 18604 30194 18656 30200
rect 18788 30252 18840 30258
rect 18788 30194 18840 30200
rect 18512 29164 18564 29170
rect 18512 29106 18564 29112
rect 18420 28416 18472 28422
rect 18420 28358 18472 28364
rect 18432 28082 18460 28358
rect 18524 28150 18552 29106
rect 18788 28484 18840 28490
rect 18788 28426 18840 28432
rect 18800 28218 18828 28426
rect 18788 28212 18840 28218
rect 18788 28154 18840 28160
rect 18512 28144 18564 28150
rect 18512 28086 18564 28092
rect 18420 28076 18472 28082
rect 18420 28018 18472 28024
rect 18604 27124 18656 27130
rect 18604 27066 18656 27072
rect 18616 26382 18644 27066
rect 18604 26376 18656 26382
rect 18604 26318 18656 26324
rect 18512 26308 18564 26314
rect 18512 26250 18564 26256
rect 18236 25696 18288 25702
rect 18236 25638 18288 25644
rect 18248 25430 18276 25638
rect 18236 25424 18288 25430
rect 18236 25366 18288 25372
rect 18420 25152 18472 25158
rect 18420 25094 18472 25100
rect 18432 24886 18460 25094
rect 18420 24880 18472 24886
rect 18420 24822 18472 24828
rect 18144 24744 18196 24750
rect 18144 24686 18196 24692
rect 17960 23724 18012 23730
rect 17960 23666 18012 23672
rect 17696 22066 17816 22094
rect 17696 16574 17724 22066
rect 17776 21956 17828 21962
rect 17776 21898 17828 21904
rect 17788 21690 17816 21898
rect 17776 21684 17828 21690
rect 17776 21626 17828 21632
rect 17972 20602 18000 23666
rect 18052 23588 18104 23594
rect 18052 23530 18104 23536
rect 18064 23322 18092 23530
rect 18052 23316 18104 23322
rect 18052 23258 18104 23264
rect 18156 23118 18184 24686
rect 18524 24138 18552 26250
rect 18788 25492 18840 25498
rect 18788 25434 18840 25440
rect 18800 25158 18828 25434
rect 18788 25152 18840 25158
rect 18788 25094 18840 25100
rect 18512 24132 18564 24138
rect 18512 24074 18564 24080
rect 18524 23798 18552 24074
rect 18512 23792 18564 23798
rect 18512 23734 18564 23740
rect 18880 23724 18932 23730
rect 18880 23666 18932 23672
rect 18420 23180 18472 23186
rect 18420 23122 18472 23128
rect 18144 23112 18196 23118
rect 18144 23054 18196 23060
rect 18052 22432 18104 22438
rect 18052 22374 18104 22380
rect 18064 21554 18092 22374
rect 18156 22030 18184 23054
rect 18432 22574 18460 23122
rect 18892 23118 18920 23666
rect 18512 23112 18564 23118
rect 18512 23054 18564 23060
rect 18880 23112 18932 23118
rect 18880 23054 18932 23060
rect 18420 22568 18472 22574
rect 18420 22510 18472 22516
rect 18524 22234 18552 23054
rect 18788 22636 18840 22642
rect 18788 22578 18840 22584
rect 18512 22228 18564 22234
rect 18512 22170 18564 22176
rect 18144 22024 18196 22030
rect 18144 21966 18196 21972
rect 18052 21548 18104 21554
rect 18052 21490 18104 21496
rect 17868 20596 17920 20602
rect 17868 20538 17920 20544
rect 17960 20596 18012 20602
rect 17960 20538 18012 20544
rect 17880 20058 17908 20538
rect 17868 20052 17920 20058
rect 17868 19994 17920 20000
rect 17972 19854 18000 20538
rect 18156 20398 18184 21966
rect 18800 21894 18828 22578
rect 18788 21888 18840 21894
rect 18788 21830 18840 21836
rect 18800 21486 18828 21830
rect 18788 21480 18840 21486
rect 18788 21422 18840 21428
rect 18144 20392 18196 20398
rect 18144 20334 18196 20340
rect 18156 19922 18184 20334
rect 18236 20256 18288 20262
rect 18236 20198 18288 20204
rect 18144 19916 18196 19922
rect 18144 19858 18196 19864
rect 17960 19848 18012 19854
rect 17960 19790 18012 19796
rect 17868 19372 17920 19378
rect 17868 19314 17920 19320
rect 17880 18630 17908 19314
rect 18156 18766 18184 19858
rect 18144 18760 18196 18766
rect 18144 18702 18196 18708
rect 18248 18698 18276 20198
rect 18892 19446 18920 23054
rect 18984 22778 19012 31726
rect 19260 30938 19288 35634
rect 19352 35086 19380 35702
rect 19340 35080 19392 35086
rect 19340 35022 19392 35028
rect 19444 33590 19472 36518
rect 19720 36106 19748 36518
rect 19708 36100 19760 36106
rect 19708 36042 19760 36048
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19996 35834 20024 36722
rect 20088 36258 20116 36790
rect 20180 36378 20208 37810
rect 20352 37120 20404 37126
rect 20352 37062 20404 37068
rect 20168 36372 20220 36378
rect 20168 36314 20220 36320
rect 20088 36230 20300 36258
rect 20168 36168 20220 36174
rect 20168 36110 20220 36116
rect 20076 36100 20128 36106
rect 20076 36042 20128 36048
rect 19984 35828 20036 35834
rect 19984 35770 20036 35776
rect 20088 35698 20116 36042
rect 19616 35692 19668 35698
rect 19616 35634 19668 35640
rect 20076 35692 20128 35698
rect 20076 35634 20128 35640
rect 19524 35488 19576 35494
rect 19524 35430 19576 35436
rect 19536 35222 19564 35430
rect 19628 35290 19656 35634
rect 19800 35556 19852 35562
rect 19800 35498 19852 35504
rect 19616 35284 19668 35290
rect 19616 35226 19668 35232
rect 19812 35222 19840 35498
rect 19524 35216 19576 35222
rect 19524 35158 19576 35164
rect 19800 35216 19852 35222
rect 19800 35158 19852 35164
rect 20088 35018 20116 35634
rect 20180 35630 20208 36110
rect 20168 35624 20220 35630
rect 20168 35566 20220 35572
rect 20076 35012 20128 35018
rect 20076 34954 20128 34960
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 20168 33992 20220 33998
rect 20168 33934 20220 33940
rect 19984 33856 20036 33862
rect 19984 33798 20036 33804
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19996 33590 20024 33798
rect 19432 33584 19484 33590
rect 19432 33526 19484 33532
rect 19984 33584 20036 33590
rect 19984 33526 20036 33532
rect 19444 31890 19472 33526
rect 20180 33114 20208 33934
rect 20168 33108 20220 33114
rect 20168 33050 20220 33056
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 20076 32360 20128 32366
rect 20076 32302 20128 32308
rect 19432 31884 19484 31890
rect 19432 31826 19484 31832
rect 19248 30932 19300 30938
rect 19248 30874 19300 30880
rect 19260 30394 19288 30874
rect 19444 30802 19472 31826
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19432 30796 19484 30802
rect 19432 30738 19484 30744
rect 19340 30660 19392 30666
rect 19340 30602 19392 30608
rect 19248 30388 19300 30394
rect 19248 30330 19300 30336
rect 19064 30252 19116 30258
rect 19064 30194 19116 30200
rect 19076 29306 19104 30194
rect 19352 30122 19380 30602
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19432 30320 19484 30326
rect 19432 30262 19484 30268
rect 19340 30116 19392 30122
rect 19340 30058 19392 30064
rect 19064 29300 19116 29306
rect 19064 29242 19116 29248
rect 19076 28082 19104 29242
rect 19444 28098 19472 30262
rect 19524 30116 19576 30122
rect 19524 30058 19576 30064
rect 19536 29714 19564 30058
rect 19524 29708 19576 29714
rect 19524 29650 19576 29656
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19064 28076 19116 28082
rect 19064 28018 19116 28024
rect 19352 28070 19472 28098
rect 19984 28076 20036 28082
rect 19352 25362 19380 28070
rect 19984 28018 20036 28024
rect 19432 28008 19484 28014
rect 19432 27950 19484 27956
rect 19444 26450 19472 27950
rect 19996 27674 20024 28018
rect 19984 27668 20036 27674
rect 19984 27610 20036 27616
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 20088 27010 20116 32302
rect 20272 30190 20300 36230
rect 20364 36174 20392 37062
rect 20352 36168 20404 36174
rect 20352 36110 20404 36116
rect 20456 31142 20484 38830
rect 20548 36768 20576 38898
rect 20640 38418 20668 39442
rect 21100 39098 21128 41386
rect 21836 41206 21864 41550
rect 21824 41200 21876 41206
rect 21824 41142 21876 41148
rect 21836 40730 21864 41142
rect 22112 41138 22140 41618
rect 22100 41132 22152 41138
rect 22100 41074 22152 41080
rect 22836 41132 22888 41138
rect 22836 41074 22888 41080
rect 22928 41132 22980 41138
rect 22928 41074 22980 41080
rect 22744 40928 22796 40934
rect 22744 40870 22796 40876
rect 21824 40724 21876 40730
rect 21824 40666 21876 40672
rect 21836 40118 21864 40666
rect 22756 40594 22784 40870
rect 22744 40588 22796 40594
rect 22744 40530 22796 40536
rect 21824 40112 21876 40118
rect 21824 40054 21876 40060
rect 22848 40050 22876 41074
rect 22940 40730 22968 41074
rect 23032 40730 23060 42570
rect 22928 40724 22980 40730
rect 22928 40666 22980 40672
rect 23020 40724 23072 40730
rect 23020 40666 23072 40672
rect 23124 40662 23152 42638
rect 24308 42560 24360 42566
rect 24308 42502 24360 42508
rect 24320 42362 24348 42502
rect 24308 42356 24360 42362
rect 24308 42298 24360 42304
rect 23664 42220 23716 42226
rect 23664 42162 23716 42168
rect 24216 42220 24268 42226
rect 24216 42162 24268 42168
rect 24676 42220 24728 42226
rect 24676 42162 24728 42168
rect 23480 42084 23532 42090
rect 23480 42026 23532 42032
rect 23204 42016 23256 42022
rect 23204 41958 23256 41964
rect 23216 41818 23244 41958
rect 23204 41812 23256 41818
rect 23204 41754 23256 41760
rect 23296 41608 23348 41614
rect 23296 41550 23348 41556
rect 23308 41274 23336 41550
rect 23296 41268 23348 41274
rect 23296 41210 23348 41216
rect 23492 41206 23520 42026
rect 23480 41200 23532 41206
rect 23480 41142 23532 41148
rect 23204 40724 23256 40730
rect 23204 40666 23256 40672
rect 23112 40656 23164 40662
rect 22940 40604 23112 40610
rect 22940 40598 23164 40604
rect 22940 40582 23152 40598
rect 22940 40526 22968 40582
rect 22928 40520 22980 40526
rect 22928 40462 22980 40468
rect 22836 40044 22888 40050
rect 22836 39986 22888 39992
rect 21088 39092 21140 39098
rect 21088 39034 21140 39040
rect 22376 39092 22428 39098
rect 22376 39034 22428 39040
rect 20628 38412 20680 38418
rect 20628 38354 20680 38360
rect 21272 38208 21324 38214
rect 21272 38150 21324 38156
rect 21284 37262 21312 38150
rect 22284 37868 22336 37874
rect 22284 37810 22336 37816
rect 21732 37664 21784 37670
rect 21732 37606 21784 37612
rect 21744 37262 21772 37606
rect 21272 37256 21324 37262
rect 21272 37198 21324 37204
rect 21548 37256 21600 37262
rect 21548 37198 21600 37204
rect 21732 37256 21784 37262
rect 21732 37198 21784 37204
rect 20628 36780 20680 36786
rect 20548 36740 20628 36768
rect 20628 36722 20680 36728
rect 20534 36680 20590 36689
rect 20534 36615 20536 36624
rect 20588 36615 20590 36624
rect 20536 36586 20588 36592
rect 21284 36582 21312 37198
rect 21272 36576 21324 36582
rect 21272 36518 21324 36524
rect 20628 36236 20680 36242
rect 20628 36178 20680 36184
rect 20536 36168 20588 36174
rect 20536 36110 20588 36116
rect 20548 34066 20576 36110
rect 20640 36009 20668 36178
rect 20626 36000 20682 36009
rect 20626 35935 20682 35944
rect 20904 35488 20956 35494
rect 20904 35430 20956 35436
rect 20536 34060 20588 34066
rect 20536 34002 20588 34008
rect 20812 34060 20864 34066
rect 20812 34002 20864 34008
rect 20444 31136 20496 31142
rect 20444 31078 20496 31084
rect 20628 30252 20680 30258
rect 20628 30194 20680 30200
rect 20260 30184 20312 30190
rect 20260 30126 20312 30132
rect 20640 29850 20668 30194
rect 20628 29844 20680 29850
rect 20628 29786 20680 29792
rect 20720 29640 20772 29646
rect 20720 29582 20772 29588
rect 20732 29510 20760 29582
rect 20720 29504 20772 29510
rect 20720 29446 20772 29452
rect 20732 29238 20760 29446
rect 20720 29232 20772 29238
rect 20720 29174 20772 29180
rect 20824 28506 20852 34002
rect 20916 33658 20944 35430
rect 21456 35012 21508 35018
rect 21456 34954 21508 34960
rect 21468 34542 21496 34954
rect 21456 34536 21508 34542
rect 21456 34478 21508 34484
rect 21456 33992 21508 33998
rect 21456 33934 21508 33940
rect 20904 33652 20956 33658
rect 20904 33594 20956 33600
rect 20916 32892 20944 33594
rect 20996 32904 21048 32910
rect 20916 32864 20996 32892
rect 20996 32846 21048 32852
rect 21180 32768 21232 32774
rect 21180 32710 21232 32716
rect 20996 31748 21048 31754
rect 20996 31690 21048 31696
rect 21008 31482 21036 31690
rect 20996 31476 21048 31482
rect 20996 31418 21048 31424
rect 21192 31346 21220 32710
rect 21468 31754 21496 33934
rect 21560 32978 21588 37198
rect 21744 36922 21772 37198
rect 21732 36916 21784 36922
rect 21732 36858 21784 36864
rect 21732 36780 21784 36786
rect 21732 36722 21784 36728
rect 21640 35148 21692 35154
rect 21640 35090 21692 35096
rect 21652 33998 21680 35090
rect 21744 35086 21772 36722
rect 22008 36712 22060 36718
rect 22008 36654 22060 36660
rect 22020 35630 22048 36654
rect 22192 36168 22244 36174
rect 22192 36110 22244 36116
rect 22204 35834 22232 36110
rect 22296 36106 22324 37810
rect 22284 36100 22336 36106
rect 22284 36042 22336 36048
rect 22192 35828 22244 35834
rect 22192 35770 22244 35776
rect 22100 35692 22152 35698
rect 22100 35634 22152 35640
rect 22008 35624 22060 35630
rect 22008 35566 22060 35572
rect 21732 35080 21784 35086
rect 21732 35022 21784 35028
rect 21640 33992 21692 33998
rect 21640 33934 21692 33940
rect 21744 33318 21772 35022
rect 21916 35012 21968 35018
rect 21916 34954 21968 34960
rect 21732 33312 21784 33318
rect 21732 33254 21784 33260
rect 21928 33114 21956 34954
rect 21916 33108 21968 33114
rect 21916 33050 21968 33056
rect 21548 32972 21600 32978
rect 21548 32914 21600 32920
rect 21560 32858 21588 32914
rect 21824 32904 21876 32910
rect 21560 32830 21772 32858
rect 21824 32846 21876 32852
rect 21744 32774 21772 32830
rect 21732 32768 21784 32774
rect 21732 32710 21784 32716
rect 21836 31822 21864 32846
rect 21928 32026 21956 33050
rect 22020 33046 22048 35566
rect 22112 34202 22140 35634
rect 22204 34950 22232 35770
rect 22388 35154 22416 39034
rect 22652 38956 22704 38962
rect 22652 38898 22704 38904
rect 22560 38752 22612 38758
rect 22560 38694 22612 38700
rect 22572 38486 22600 38694
rect 22560 38480 22612 38486
rect 22560 38422 22612 38428
rect 22560 38276 22612 38282
rect 22560 38218 22612 38224
rect 22468 38208 22520 38214
rect 22468 38150 22520 38156
rect 22480 37874 22508 38150
rect 22468 37868 22520 37874
rect 22468 37810 22520 37816
rect 22480 37398 22508 37810
rect 22572 37738 22600 38218
rect 22560 37732 22612 37738
rect 22560 37674 22612 37680
rect 22664 37466 22692 38898
rect 22744 38752 22796 38758
rect 22744 38694 22796 38700
rect 22756 37942 22784 38694
rect 22928 38344 22980 38350
rect 22928 38286 22980 38292
rect 22836 38208 22888 38214
rect 22836 38150 22888 38156
rect 22744 37936 22796 37942
rect 22744 37878 22796 37884
rect 22652 37460 22704 37466
rect 22652 37402 22704 37408
rect 22468 37392 22520 37398
rect 22848 37346 22876 38150
rect 22940 37913 22968 38286
rect 22926 37904 22982 37913
rect 22926 37839 22982 37848
rect 22468 37334 22520 37340
rect 22480 36786 22508 37334
rect 22664 37318 22876 37346
rect 22664 37194 22692 37318
rect 22652 37188 22704 37194
rect 22836 37188 22888 37194
rect 22652 37130 22704 37136
rect 22756 37148 22836 37176
rect 22468 36780 22520 36786
rect 22468 36722 22520 36728
rect 22652 36168 22704 36174
rect 22652 36110 22704 36116
rect 22664 35494 22692 36110
rect 22756 36038 22784 37148
rect 22940 37176 22968 37839
rect 22888 37148 22968 37176
rect 22836 37130 22888 37136
rect 23032 36961 23060 40582
rect 23112 40520 23164 40526
rect 23112 40462 23164 40468
rect 23124 40118 23152 40462
rect 23216 40458 23244 40666
rect 23204 40452 23256 40458
rect 23204 40394 23256 40400
rect 23492 40390 23520 41142
rect 23676 40526 23704 42162
rect 24228 42022 24256 42162
rect 24216 42016 24268 42022
rect 24216 41958 24268 41964
rect 24124 41608 24176 41614
rect 24124 41550 24176 41556
rect 24136 41206 24164 41550
rect 24228 41546 24256 41958
rect 24216 41540 24268 41546
rect 24216 41482 24268 41488
rect 24308 41472 24360 41478
rect 24308 41414 24360 41420
rect 24320 41274 24348 41414
rect 24308 41268 24360 41274
rect 24308 41210 24360 41216
rect 24124 41200 24176 41206
rect 24124 41142 24176 41148
rect 24320 41138 24348 41210
rect 24308 41132 24360 41138
rect 24308 41074 24360 41080
rect 23756 41064 23808 41070
rect 23756 41006 23808 41012
rect 23768 40730 23796 41006
rect 24688 40934 24716 42162
rect 24768 41540 24820 41546
rect 24768 41482 24820 41488
rect 24780 41138 24808 41482
rect 25424 41414 25452 46922
rect 25700 46646 25728 46990
rect 25688 46640 25740 46646
rect 25688 46582 25740 46588
rect 25792 46510 25820 49200
rect 25780 46504 25832 46510
rect 25780 46446 25832 46452
rect 27080 43858 27108 49200
rect 29656 46510 29684 49200
rect 29736 47048 29788 47054
rect 29736 46990 29788 46996
rect 29184 46504 29236 46510
rect 29184 46446 29236 46452
rect 29644 46504 29696 46510
rect 29644 46446 29696 46452
rect 29196 46170 29224 46446
rect 29184 46164 29236 46170
rect 29184 46106 29236 46112
rect 29748 45966 29776 46990
rect 29184 45960 29236 45966
rect 29184 45902 29236 45908
rect 29736 45960 29788 45966
rect 29736 45902 29788 45908
rect 29196 45490 29224 45902
rect 30300 45898 30328 49200
rect 31588 47138 31616 49200
rect 32220 47184 32272 47190
rect 31588 47110 31800 47138
rect 32220 47126 32272 47132
rect 31772 47054 31800 47110
rect 31760 47048 31812 47054
rect 31760 46990 31812 46996
rect 29920 45892 29972 45898
rect 29920 45834 29972 45840
rect 30288 45892 30340 45898
rect 30288 45834 30340 45840
rect 29932 45626 29960 45834
rect 29920 45620 29972 45626
rect 29920 45562 29972 45568
rect 29184 45484 29236 45490
rect 29184 45426 29236 45432
rect 29736 45484 29788 45490
rect 29736 45426 29788 45432
rect 27068 43852 27120 43858
rect 27068 43794 27120 43800
rect 27160 43376 27212 43382
rect 27160 43318 27212 43324
rect 25504 43308 25556 43314
rect 25504 43250 25556 43256
rect 26240 43308 26292 43314
rect 26240 43250 26292 43256
rect 25516 42362 25544 43250
rect 26148 43240 26200 43246
rect 26148 43182 26200 43188
rect 26056 43104 26108 43110
rect 26056 43046 26108 43052
rect 26068 42634 26096 43046
rect 26056 42628 26108 42634
rect 26056 42570 26108 42576
rect 26160 42566 26188 43182
rect 26148 42560 26200 42566
rect 26148 42502 26200 42508
rect 25504 42356 25556 42362
rect 25504 42298 25556 42304
rect 26160 42158 26188 42502
rect 26148 42152 26200 42158
rect 26148 42094 26200 42100
rect 26160 41682 26188 42094
rect 26148 41676 26200 41682
rect 26148 41618 26200 41624
rect 25780 41608 25832 41614
rect 25780 41550 25832 41556
rect 25424 41386 25544 41414
rect 24768 41132 24820 41138
rect 24768 41074 24820 41080
rect 24676 40928 24728 40934
rect 24676 40870 24728 40876
rect 23756 40724 23808 40730
rect 23756 40666 23808 40672
rect 24688 40526 24716 40870
rect 23664 40520 23716 40526
rect 23664 40462 23716 40468
rect 24676 40520 24728 40526
rect 24676 40462 24728 40468
rect 23480 40384 23532 40390
rect 23480 40326 23532 40332
rect 23112 40112 23164 40118
rect 23112 40054 23164 40060
rect 23676 39982 23704 40462
rect 23664 39976 23716 39982
rect 23664 39918 23716 39924
rect 25412 39024 25464 39030
rect 25412 38966 25464 38972
rect 24216 38956 24268 38962
rect 24216 38898 24268 38904
rect 25044 38956 25096 38962
rect 25044 38898 25096 38904
rect 25320 38956 25372 38962
rect 25320 38898 25372 38904
rect 23388 38888 23440 38894
rect 23388 38830 23440 38836
rect 23112 38548 23164 38554
rect 23112 38490 23164 38496
rect 23124 37738 23152 38490
rect 23400 37777 23428 38830
rect 23480 38820 23532 38826
rect 23480 38762 23532 38768
rect 23492 38350 23520 38762
rect 23572 38752 23624 38758
rect 23572 38694 23624 38700
rect 23480 38344 23532 38350
rect 23480 38286 23532 38292
rect 23492 37806 23520 38286
rect 23584 38282 23612 38694
rect 24228 38554 24256 38898
rect 24952 38888 25004 38894
rect 24952 38830 25004 38836
rect 24860 38752 24912 38758
rect 24860 38694 24912 38700
rect 24872 38554 24900 38694
rect 24216 38548 24268 38554
rect 24216 38490 24268 38496
rect 24860 38548 24912 38554
rect 24860 38490 24912 38496
rect 23848 38480 23900 38486
rect 23848 38422 23900 38428
rect 23940 38480 23992 38486
rect 23940 38422 23992 38428
rect 23572 38276 23624 38282
rect 23572 38218 23624 38224
rect 23860 37913 23888 38422
rect 23846 37904 23902 37913
rect 23846 37839 23848 37848
rect 23900 37839 23902 37848
rect 23848 37810 23900 37816
rect 23952 37806 23980 38422
rect 24860 38412 24912 38418
rect 24860 38354 24912 38360
rect 24872 38010 24900 38354
rect 24964 38214 24992 38830
rect 25056 38554 25084 38898
rect 25136 38888 25188 38894
rect 25136 38830 25188 38836
rect 25044 38548 25096 38554
rect 25044 38490 25096 38496
rect 25148 38434 25176 38830
rect 25056 38406 25176 38434
rect 24952 38208 25004 38214
rect 24952 38150 25004 38156
rect 24860 38004 24912 38010
rect 24860 37946 24912 37952
rect 23480 37800 23532 37806
rect 23386 37768 23442 37777
rect 23112 37732 23164 37738
rect 23940 37800 23992 37806
rect 23480 37742 23532 37748
rect 23938 37768 23940 37777
rect 23992 37768 23994 37777
rect 23386 37703 23442 37712
rect 23112 37674 23164 37680
rect 23124 37262 23152 37674
rect 23112 37256 23164 37262
rect 23112 37198 23164 37204
rect 23018 36952 23074 36961
rect 23018 36887 23074 36896
rect 22836 36100 22888 36106
rect 22836 36042 22888 36048
rect 22744 36032 22796 36038
rect 22744 35974 22796 35980
rect 22652 35488 22704 35494
rect 22652 35430 22704 35436
rect 22376 35148 22428 35154
rect 22376 35090 22428 35096
rect 22664 35086 22692 35430
rect 22284 35080 22336 35086
rect 22284 35022 22336 35028
rect 22652 35080 22704 35086
rect 22652 35022 22704 35028
rect 22192 34944 22244 34950
rect 22192 34886 22244 34892
rect 22296 34746 22324 35022
rect 22468 34944 22520 34950
rect 22468 34886 22520 34892
rect 22284 34740 22336 34746
rect 22284 34682 22336 34688
rect 22192 34536 22244 34542
rect 22192 34478 22244 34484
rect 22100 34196 22152 34202
rect 22100 34138 22152 34144
rect 22008 33040 22060 33046
rect 22008 32982 22060 32988
rect 22100 33040 22152 33046
rect 22100 32982 22152 32988
rect 22020 32434 22048 32982
rect 22112 32774 22140 32982
rect 22100 32768 22152 32774
rect 22100 32710 22152 32716
rect 22008 32428 22060 32434
rect 22008 32370 22060 32376
rect 22100 32428 22152 32434
rect 22100 32370 22152 32376
rect 21916 32020 21968 32026
rect 21916 31962 21968 31968
rect 21824 31816 21876 31822
rect 21824 31758 21876 31764
rect 21468 31726 21588 31754
rect 21180 31340 21232 31346
rect 21180 31282 21232 31288
rect 21560 31278 21588 31726
rect 22112 31482 22140 32370
rect 22100 31476 22152 31482
rect 22100 31418 22152 31424
rect 21548 31272 21600 31278
rect 21548 31214 21600 31220
rect 21272 29640 21324 29646
rect 21272 29582 21324 29588
rect 21284 29034 21312 29582
rect 21364 29504 21416 29510
rect 21364 29446 21416 29452
rect 21272 29028 21324 29034
rect 21272 28970 21324 28976
rect 20732 28478 20852 28506
rect 20168 28416 20220 28422
rect 20168 28358 20220 28364
rect 20180 27470 20208 28358
rect 20168 27464 20220 27470
rect 20168 27406 20220 27412
rect 19996 26982 20116 27010
rect 20732 26994 20760 28478
rect 20812 28416 20864 28422
rect 20812 28358 20864 28364
rect 20904 28416 20956 28422
rect 20904 28358 20956 28364
rect 20824 28218 20852 28358
rect 20916 28218 20944 28358
rect 20812 28212 20864 28218
rect 20812 28154 20864 28160
rect 20904 28212 20956 28218
rect 20904 28154 20956 28160
rect 20824 27470 20852 28154
rect 21284 27606 21312 28970
rect 21376 28150 21404 29446
rect 21364 28144 21416 28150
rect 21364 28086 21416 28092
rect 21456 28076 21508 28082
rect 21456 28018 21508 28024
rect 21364 28008 21416 28014
rect 21364 27950 21416 27956
rect 21272 27600 21324 27606
rect 21272 27542 21324 27548
rect 20812 27464 20864 27470
rect 20812 27406 20864 27412
rect 21088 27464 21140 27470
rect 21088 27406 21140 27412
rect 20536 26988 20588 26994
rect 19432 26444 19484 26450
rect 19432 26386 19484 26392
rect 19340 25356 19392 25362
rect 19340 25298 19392 25304
rect 19248 25288 19300 25294
rect 19248 25230 19300 25236
rect 19260 24206 19288 25230
rect 19352 24954 19380 25298
rect 19340 24948 19392 24954
rect 19340 24890 19392 24896
rect 19248 24200 19300 24206
rect 19248 24142 19300 24148
rect 19444 23798 19472 26386
rect 19996 26246 20024 26982
rect 20536 26930 20588 26936
rect 20720 26988 20772 26994
rect 20720 26930 20772 26936
rect 20352 26784 20404 26790
rect 20352 26726 20404 26732
rect 20364 26382 20392 26726
rect 20352 26376 20404 26382
rect 20352 26318 20404 26324
rect 19984 26240 20036 26246
rect 19984 26182 20036 26188
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19996 25294 20024 26182
rect 20548 26042 20576 26930
rect 20732 26586 20760 26930
rect 21100 26586 21128 27406
rect 20720 26580 20772 26586
rect 20720 26522 20772 26528
rect 21088 26580 21140 26586
rect 21088 26522 21140 26528
rect 20628 26308 20680 26314
rect 20628 26250 20680 26256
rect 20536 26036 20588 26042
rect 20536 25978 20588 25984
rect 19984 25288 20036 25294
rect 19984 25230 20036 25236
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19996 24818 20024 25230
rect 19984 24812 20036 24818
rect 19984 24754 20036 24760
rect 20260 24812 20312 24818
rect 20260 24754 20312 24760
rect 20272 24138 20300 24754
rect 20640 24206 20668 26250
rect 21100 25906 21128 26522
rect 21088 25900 21140 25906
rect 21088 25842 21140 25848
rect 20812 25492 20864 25498
rect 20812 25434 20864 25440
rect 20824 25226 20852 25434
rect 21376 25294 21404 27950
rect 21468 27470 21496 28018
rect 21456 27464 21508 27470
rect 21456 27406 21508 27412
rect 21364 25288 21416 25294
rect 21364 25230 21416 25236
rect 20812 25220 20864 25226
rect 20812 25162 20864 25168
rect 20628 24200 20680 24206
rect 20628 24142 20680 24148
rect 20260 24132 20312 24138
rect 20260 24074 20312 24080
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19432 23792 19484 23798
rect 19432 23734 19484 23740
rect 20168 23792 20220 23798
rect 20168 23734 20220 23740
rect 19444 23186 19472 23734
rect 19432 23180 19484 23186
rect 19432 23122 19484 23128
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 20180 22778 20208 23734
rect 18972 22772 19024 22778
rect 18972 22714 19024 22720
rect 20168 22772 20220 22778
rect 20168 22714 20220 22720
rect 19340 22568 19392 22574
rect 19340 22510 19392 22516
rect 19064 20460 19116 20466
rect 19064 20402 19116 20408
rect 19076 19514 19104 20402
rect 19352 19922 19380 22510
rect 20272 21962 20300 24074
rect 20536 22976 20588 22982
rect 20536 22918 20588 22924
rect 20548 22778 20576 22918
rect 20536 22772 20588 22778
rect 20536 22714 20588 22720
rect 20260 21956 20312 21962
rect 20260 21898 20312 21904
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19984 20936 20036 20942
rect 19984 20878 20036 20884
rect 19432 20800 19484 20806
rect 19432 20742 19484 20748
rect 19444 20534 19472 20742
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19432 20528 19484 20534
rect 19432 20470 19484 20476
rect 19340 19916 19392 19922
rect 19340 19858 19392 19864
rect 19064 19508 19116 19514
rect 19064 19450 19116 19456
rect 18880 19440 18932 19446
rect 18880 19382 18932 19388
rect 18236 18692 18288 18698
rect 18236 18634 18288 18640
rect 17868 18624 17920 18630
rect 17868 18566 17920 18572
rect 17880 18358 17908 18566
rect 17868 18352 17920 18358
rect 17868 18294 17920 18300
rect 18696 18080 18748 18086
rect 18696 18022 18748 18028
rect 18708 17814 18736 18022
rect 18696 17808 18748 17814
rect 18696 17750 18748 17756
rect 18892 17678 18920 19382
rect 19352 19310 19380 19858
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19996 19514 20024 20878
rect 20076 19712 20128 19718
rect 20076 19654 20128 19660
rect 19984 19508 20036 19514
rect 19984 19450 20036 19456
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 19064 18284 19116 18290
rect 19064 18226 19116 18232
rect 18512 17672 18564 17678
rect 18512 17614 18564 17620
rect 18880 17672 18932 17678
rect 18880 17614 18932 17620
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 17696 16546 17816 16574
rect 17592 16040 17644 16046
rect 17592 15982 17644 15988
rect 17684 16040 17736 16046
rect 17684 15982 17736 15988
rect 17512 15638 17540 15669
rect 17500 15632 17552 15638
rect 17420 15580 17500 15586
rect 17420 15574 17552 15580
rect 17420 15558 17540 15574
rect 17040 15496 17092 15502
rect 17040 15438 17092 15444
rect 17408 15496 17460 15502
rect 17408 15438 17460 15444
rect 17132 15360 17184 15366
rect 17132 15302 17184 15308
rect 13912 15020 13964 15026
rect 13912 14962 13964 14968
rect 16764 15020 16816 15026
rect 16764 14962 16816 14968
rect 16120 14816 16172 14822
rect 16120 14758 16172 14764
rect 16132 14346 16160 14758
rect 16776 14414 16804 14962
rect 17144 14890 17172 15302
rect 17132 14884 17184 14890
rect 17132 14826 17184 14832
rect 17420 14618 17448 15438
rect 17512 15366 17540 15558
rect 17500 15360 17552 15366
rect 17500 15302 17552 15308
rect 17408 14612 17460 14618
rect 17408 14554 17460 14560
rect 16764 14408 16816 14414
rect 16764 14350 16816 14356
rect 16120 14340 16172 14346
rect 16120 14282 16172 14288
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12544 10742 12572 10950
rect 12532 10736 12584 10742
rect 12532 10678 12584 10684
rect 12636 10606 12664 11086
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 13268 4072 13320 4078
rect 13268 4014 13320 4020
rect 10140 4004 10192 4010
rect 10140 3946 10192 3952
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 9864 3664 9916 3670
rect 9864 3606 9916 3612
rect 10704 3602 10732 3878
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 10508 3528 10560 3534
rect 10508 3470 10560 3476
rect 9588 3460 9640 3466
rect 9588 3402 9640 3408
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 7472 3120 7524 3126
rect 7472 3062 7524 3068
rect 10520 3058 10548 3470
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 6828 2848 6880 2854
rect 6828 2790 6880 2796
rect 6840 2514 6868 2790
rect 6828 2508 6880 2514
rect 6828 2450 6880 2456
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 6748 2378 6868 2394
rect 6748 2372 6880 2378
rect 6748 2366 6828 2372
rect 6828 2314 6880 2320
rect 7116 800 7144 2450
rect 7760 800 7788 2926
rect 10980 800 11008 3538
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 11624 800 11652 2382
rect 12912 800 12940 3674
rect 13004 3058 13032 3878
rect 13280 3398 13308 4014
rect 14200 3738 14228 10542
rect 16120 5704 16172 5710
rect 16120 5646 16172 5652
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 16132 3670 16160 5646
rect 17132 4072 17184 4078
rect 17132 4014 17184 4020
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16120 3664 16172 3670
rect 16120 3606 16172 3612
rect 16132 3534 16160 3606
rect 16776 3602 16804 3878
rect 16764 3596 16816 3602
rect 16764 3538 16816 3544
rect 16120 3528 16172 3534
rect 16120 3470 16172 3476
rect 17144 3466 17172 4014
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 17132 3460 17184 3466
rect 17132 3402 17184 3408
rect 13176 3392 13228 3398
rect 13176 3334 13228 3340
rect 13268 3392 13320 3398
rect 13268 3334 13320 3340
rect 13188 3126 13216 3334
rect 13176 3120 13228 3126
rect 13176 3062 13228 3068
rect 17328 3058 17356 3878
rect 17408 3596 17460 3602
rect 17408 3538 17460 3544
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 17316 3052 17368 3058
rect 17316 2994 17368 3000
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 13556 800 13584 2926
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 14200 800 14228 2382
rect 17420 800 17448 3538
rect 17512 2038 17540 15302
rect 17604 2650 17632 15982
rect 17696 15570 17724 15982
rect 17684 15564 17736 15570
rect 17684 15506 17736 15512
rect 17592 2644 17644 2650
rect 17592 2586 17644 2592
rect 17788 2582 17816 16546
rect 18340 16232 18368 17138
rect 18420 17128 18472 17134
rect 18420 17070 18472 17076
rect 18432 16726 18460 17070
rect 18420 16720 18472 16726
rect 18420 16662 18472 16668
rect 18524 16574 18552 17614
rect 19076 17338 19104 18226
rect 19352 18222 19380 19246
rect 20088 19242 20116 19654
rect 20272 19446 20300 21898
rect 20548 20058 20576 22714
rect 20640 21622 20668 24142
rect 21376 24070 21404 25230
rect 21364 24064 21416 24070
rect 21364 24006 21416 24012
rect 21456 23520 21508 23526
rect 21456 23462 21508 23468
rect 21468 23118 21496 23462
rect 21456 23112 21508 23118
rect 21456 23054 21508 23060
rect 21456 21888 21508 21894
rect 21456 21830 21508 21836
rect 21468 21690 21496 21830
rect 21456 21684 21508 21690
rect 21456 21626 21508 21632
rect 20628 21616 20680 21622
rect 20628 21558 20680 21564
rect 20628 20324 20680 20330
rect 20628 20266 20680 20272
rect 20536 20052 20588 20058
rect 20536 19994 20588 20000
rect 20640 19854 20668 20266
rect 20628 19848 20680 19854
rect 20628 19790 20680 19796
rect 20260 19440 20312 19446
rect 20260 19382 20312 19388
rect 20076 19236 20128 19242
rect 20076 19178 20128 19184
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19340 18216 19392 18222
rect 19340 18158 19392 18164
rect 19064 17332 19116 17338
rect 19064 17274 19116 17280
rect 18524 16546 18644 16574
rect 18420 16244 18472 16250
rect 18340 16204 18420 16232
rect 18420 16186 18472 16192
rect 18616 16114 18644 16546
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 18880 16108 18932 16114
rect 18880 16050 18932 16056
rect 18616 15434 18644 16050
rect 18892 15706 18920 16050
rect 19156 15904 19208 15910
rect 19156 15846 19208 15852
rect 18880 15700 18932 15706
rect 18880 15642 18932 15648
rect 18604 15428 18656 15434
rect 18604 15370 18656 15376
rect 18616 15094 18644 15370
rect 19168 15094 19196 15846
rect 19352 15570 19380 18158
rect 19432 17536 19484 17542
rect 19432 17478 19484 17484
rect 19444 17270 19472 17478
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19432 17264 19484 17270
rect 19432 17206 19484 17212
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 19984 15428 20036 15434
rect 19984 15370 20036 15376
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19996 15162 20024 15370
rect 19984 15156 20036 15162
rect 19984 15098 20036 15104
rect 18604 15088 18656 15094
rect 18604 15030 18656 15036
rect 19156 15088 19208 15094
rect 19156 15030 19208 15036
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 20996 13728 21048 13734
rect 20996 13670 21048 13676
rect 21008 13258 21036 13670
rect 21560 13530 21588 31214
rect 21640 30048 21692 30054
rect 21640 29990 21692 29996
rect 21652 29714 21680 29990
rect 22204 29850 22232 34478
rect 22480 33998 22508 34886
rect 22652 34740 22704 34746
rect 22652 34682 22704 34688
rect 22560 34604 22612 34610
rect 22560 34546 22612 34552
rect 22572 34406 22600 34546
rect 22560 34400 22612 34406
rect 22560 34342 22612 34348
rect 22468 33992 22520 33998
rect 22468 33934 22520 33940
rect 22284 33108 22336 33114
rect 22284 33050 22336 33056
rect 22296 32910 22324 33050
rect 22284 32904 22336 32910
rect 22284 32846 22336 32852
rect 22376 32836 22428 32842
rect 22376 32778 22428 32784
rect 22388 31754 22416 32778
rect 22376 31748 22428 31754
rect 22376 31690 22428 31696
rect 22284 31680 22336 31686
rect 22284 31622 22336 31628
rect 22296 31346 22324 31622
rect 22466 31376 22522 31385
rect 22284 31340 22336 31346
rect 22466 31311 22522 31320
rect 22284 31282 22336 31288
rect 22480 31278 22508 31311
rect 22468 31272 22520 31278
rect 22468 31214 22520 31220
rect 22376 31204 22428 31210
rect 22376 31146 22428 31152
rect 22388 30326 22416 31146
rect 22376 30320 22428 30326
rect 22376 30262 22428 30268
rect 22468 30252 22520 30258
rect 22468 30194 22520 30200
rect 22480 30054 22508 30194
rect 22572 30122 22600 34342
rect 22664 34202 22692 34682
rect 22652 34196 22704 34202
rect 22652 34138 22704 34144
rect 22756 33998 22784 35974
rect 22744 33992 22796 33998
rect 22744 33934 22796 33940
rect 22848 33114 22876 36042
rect 23124 35018 23152 37198
rect 23400 36922 23428 37703
rect 23492 37466 23520 37742
rect 23938 37703 23994 37712
rect 24768 37664 24820 37670
rect 24768 37606 24820 37612
rect 23480 37460 23532 37466
rect 23480 37402 23532 37408
rect 24780 37262 24808 37606
rect 23572 37256 23624 37262
rect 23572 37198 23624 37204
rect 24768 37256 24820 37262
rect 24768 37198 24820 37204
rect 23388 36916 23440 36922
rect 23388 36858 23440 36864
rect 23584 36854 23612 37198
rect 23572 36848 23624 36854
rect 23572 36790 23624 36796
rect 24582 36816 24638 36825
rect 24582 36751 24584 36760
rect 24636 36751 24638 36760
rect 24584 36722 24636 36728
rect 24780 36310 24808 37198
rect 25056 37194 25084 38406
rect 25332 38010 25360 38898
rect 25320 38004 25372 38010
rect 25320 37946 25372 37952
rect 25044 37188 25096 37194
rect 25044 37130 25096 37136
rect 24768 36304 24820 36310
rect 24768 36246 24820 36252
rect 25056 36174 25084 37130
rect 25136 37120 25188 37126
rect 25136 37062 25188 37068
rect 25044 36168 25096 36174
rect 25044 36110 25096 36116
rect 23296 35828 23348 35834
rect 23296 35770 23348 35776
rect 23308 35018 23336 35770
rect 24584 35488 24636 35494
rect 24584 35430 24636 35436
rect 23388 35284 23440 35290
rect 23388 35226 23440 35232
rect 23112 35012 23164 35018
rect 23112 34954 23164 34960
rect 23296 35012 23348 35018
rect 23296 34954 23348 34960
rect 23400 34746 23428 35226
rect 24400 35012 24452 35018
rect 24400 34954 24452 34960
rect 23664 34944 23716 34950
rect 23664 34886 23716 34892
rect 23388 34740 23440 34746
rect 23388 34682 23440 34688
rect 23676 34066 23704 34886
rect 24412 34746 24440 34954
rect 24400 34740 24452 34746
rect 24400 34682 24452 34688
rect 24596 34610 24624 35430
rect 25148 34610 25176 37062
rect 25228 36032 25280 36038
rect 25228 35974 25280 35980
rect 25240 35834 25268 35974
rect 25228 35828 25280 35834
rect 25228 35770 25280 35776
rect 25424 35630 25452 38966
rect 25516 38434 25544 41386
rect 25792 41206 25820 41550
rect 25964 41540 26016 41546
rect 25964 41482 26016 41488
rect 25780 41200 25832 41206
rect 25780 41142 25832 41148
rect 25688 40996 25740 41002
rect 25688 40938 25740 40944
rect 25700 40526 25728 40938
rect 25792 40594 25820 41142
rect 25976 41002 26004 41482
rect 25964 40996 26016 41002
rect 25964 40938 26016 40944
rect 25780 40588 25832 40594
rect 25780 40530 25832 40536
rect 25688 40520 25740 40526
rect 25688 40462 25740 40468
rect 25700 40118 25728 40462
rect 25792 40186 25820 40530
rect 25780 40180 25832 40186
rect 25780 40122 25832 40128
rect 25688 40112 25740 40118
rect 25688 40054 25740 40060
rect 26252 39982 26280 43250
rect 27172 42906 27200 43318
rect 29000 43308 29052 43314
rect 29000 43250 29052 43256
rect 27160 42900 27212 42906
rect 27160 42842 27212 42848
rect 27528 42764 27580 42770
rect 27528 42706 27580 42712
rect 27068 42696 27120 42702
rect 27068 42638 27120 42644
rect 27252 42696 27304 42702
rect 27252 42638 27304 42644
rect 27080 42022 27108 42638
rect 27264 42226 27292 42638
rect 27540 42226 27568 42706
rect 29012 42294 29040 43250
rect 29092 43240 29144 43246
rect 29092 43182 29144 43188
rect 29104 42838 29132 43182
rect 29092 42832 29144 42838
rect 29092 42774 29144 42780
rect 29000 42288 29052 42294
rect 29000 42230 29052 42236
rect 27252 42220 27304 42226
rect 27252 42162 27304 42168
rect 27528 42220 27580 42226
rect 27528 42162 27580 42168
rect 27068 42016 27120 42022
rect 27068 41958 27120 41964
rect 27160 42016 27212 42022
rect 27160 41958 27212 41964
rect 26976 41608 27028 41614
rect 26976 41550 27028 41556
rect 26988 41138 27016 41550
rect 27080 41274 27108 41958
rect 27172 41614 27200 41958
rect 27160 41608 27212 41614
rect 27160 41550 27212 41556
rect 27068 41268 27120 41274
rect 27068 41210 27120 41216
rect 26976 41132 27028 41138
rect 26976 41074 27028 41080
rect 26792 41064 26844 41070
rect 26792 41006 26844 41012
rect 26804 40526 26832 41006
rect 26988 40594 27016 41074
rect 26976 40588 27028 40594
rect 26976 40530 27028 40536
rect 26516 40520 26568 40526
rect 26516 40462 26568 40468
rect 26792 40520 26844 40526
rect 26792 40462 26844 40468
rect 27068 40520 27120 40526
rect 27068 40462 27120 40468
rect 26528 40390 26556 40462
rect 26516 40384 26568 40390
rect 26516 40326 26568 40332
rect 26700 40384 26752 40390
rect 26700 40326 26752 40332
rect 26240 39976 26292 39982
rect 26240 39918 26292 39924
rect 25596 39908 25648 39914
rect 25596 39850 25648 39856
rect 25608 38826 25636 39850
rect 26528 39574 26556 40326
rect 26712 40118 26740 40326
rect 26700 40112 26752 40118
rect 26700 40054 26752 40060
rect 26516 39568 26568 39574
rect 26516 39510 26568 39516
rect 26804 39506 26832 40462
rect 26884 40452 26936 40458
rect 26884 40394 26936 40400
rect 26792 39500 26844 39506
rect 26792 39442 26844 39448
rect 26896 39438 26924 40394
rect 26884 39432 26936 39438
rect 26884 39374 26936 39380
rect 27080 38894 27108 40462
rect 27540 40458 27568 42162
rect 27804 41540 27856 41546
rect 27804 41482 27856 41488
rect 27528 40452 27580 40458
rect 27528 40394 27580 40400
rect 27712 40384 27764 40390
rect 27712 40326 27764 40332
rect 27724 40186 27752 40326
rect 27816 40186 27844 41482
rect 28448 41064 28500 41070
rect 28448 41006 28500 41012
rect 28460 40458 28488 41006
rect 28448 40452 28500 40458
rect 28448 40394 28500 40400
rect 27712 40180 27764 40186
rect 27712 40122 27764 40128
rect 27804 40180 27856 40186
rect 27804 40122 27856 40128
rect 27160 40044 27212 40050
rect 27160 39986 27212 39992
rect 27528 40044 27580 40050
rect 27528 39986 27580 39992
rect 27172 39642 27200 39986
rect 27160 39636 27212 39642
rect 27160 39578 27212 39584
rect 26148 38888 26200 38894
rect 26068 38836 26148 38842
rect 26068 38830 26200 38836
rect 27068 38888 27120 38894
rect 27068 38830 27120 38836
rect 25596 38820 25648 38826
rect 25596 38762 25648 38768
rect 26068 38814 26188 38830
rect 25516 38406 25636 38434
rect 25504 38276 25556 38282
rect 25504 38218 25556 38224
rect 25516 36786 25544 38218
rect 25504 36780 25556 36786
rect 25504 36722 25556 36728
rect 25412 35624 25464 35630
rect 25412 35566 25464 35572
rect 25424 34610 25452 35566
rect 24584 34604 24636 34610
rect 24584 34546 24636 34552
rect 25136 34604 25188 34610
rect 25136 34546 25188 34552
rect 25412 34604 25464 34610
rect 25412 34546 25464 34552
rect 23664 34060 23716 34066
rect 23664 34002 23716 34008
rect 23204 33312 23256 33318
rect 23204 33254 23256 33260
rect 22836 33108 22888 33114
rect 22836 33050 22888 33056
rect 23216 32910 23244 33254
rect 24584 32972 24636 32978
rect 24584 32914 24636 32920
rect 23020 32904 23072 32910
rect 23020 32846 23072 32852
rect 23204 32904 23256 32910
rect 23256 32864 23336 32892
rect 23204 32846 23256 32852
rect 23032 30326 23060 32846
rect 23204 31272 23256 31278
rect 23204 31214 23256 31220
rect 23020 30320 23072 30326
rect 23020 30262 23072 30268
rect 22560 30116 22612 30122
rect 22560 30058 22612 30064
rect 22652 30116 22704 30122
rect 22652 30058 22704 30064
rect 22376 30048 22428 30054
rect 22376 29990 22428 29996
rect 22468 30048 22520 30054
rect 22468 29990 22520 29996
rect 22388 29850 22416 29990
rect 22192 29844 22244 29850
rect 22192 29786 22244 29792
rect 22376 29844 22428 29850
rect 22376 29786 22428 29792
rect 21640 29708 21692 29714
rect 21640 29650 21692 29656
rect 22388 29170 22416 29786
rect 22480 29782 22508 29990
rect 22468 29776 22520 29782
rect 22468 29718 22520 29724
rect 22664 29170 22692 30058
rect 22836 29640 22888 29646
rect 22836 29582 22888 29588
rect 22848 29306 22876 29582
rect 23032 29578 23060 30262
rect 23216 29594 23244 31214
rect 23308 30394 23336 32864
rect 23940 32836 23992 32842
rect 23940 32778 23992 32784
rect 23388 32768 23440 32774
rect 23388 32710 23440 32716
rect 23400 32570 23428 32710
rect 23952 32570 23980 32778
rect 23388 32564 23440 32570
rect 23388 32506 23440 32512
rect 23940 32564 23992 32570
rect 23940 32506 23992 32512
rect 24400 32564 24452 32570
rect 24400 32506 24452 32512
rect 23400 31822 23428 32506
rect 24412 32366 24440 32506
rect 24596 32366 24624 32914
rect 24952 32428 25004 32434
rect 24952 32370 25004 32376
rect 24400 32360 24452 32366
rect 24400 32302 24452 32308
rect 24584 32360 24636 32366
rect 24584 32302 24636 32308
rect 24308 32224 24360 32230
rect 24308 32166 24360 32172
rect 24320 32026 24348 32166
rect 23940 32020 23992 32026
rect 23940 31962 23992 31968
rect 24308 32020 24360 32026
rect 24308 31962 24360 31968
rect 23388 31816 23440 31822
rect 23388 31758 23440 31764
rect 23756 31816 23808 31822
rect 23756 31758 23808 31764
rect 23768 31482 23796 31758
rect 23756 31476 23808 31482
rect 23756 31418 23808 31424
rect 23952 31142 23980 31962
rect 24412 31754 24440 32302
rect 24596 31890 24624 32302
rect 24964 32026 24992 32370
rect 24952 32020 25004 32026
rect 24952 31962 25004 31968
rect 24584 31884 24636 31890
rect 24584 31826 24636 31832
rect 24320 31726 24440 31754
rect 23940 31136 23992 31142
rect 23940 31078 23992 31084
rect 23296 30388 23348 30394
rect 23296 30330 23348 30336
rect 23756 30388 23808 30394
rect 23756 30330 23808 30336
rect 23572 30320 23624 30326
rect 23572 30262 23624 30268
rect 23296 30048 23348 30054
rect 23296 29990 23348 29996
rect 23308 29782 23336 29990
rect 23480 29844 23532 29850
rect 23480 29786 23532 29792
rect 23296 29776 23348 29782
rect 23296 29718 23348 29724
rect 23020 29572 23072 29578
rect 23216 29566 23336 29594
rect 23020 29514 23072 29520
rect 23204 29504 23256 29510
rect 23204 29446 23256 29452
rect 22836 29300 22888 29306
rect 22836 29242 22888 29248
rect 23216 29170 23244 29446
rect 22376 29164 22428 29170
rect 22376 29106 22428 29112
rect 22652 29164 22704 29170
rect 22652 29106 22704 29112
rect 23204 29164 23256 29170
rect 23204 29106 23256 29112
rect 22388 29050 22416 29106
rect 22100 29028 22152 29034
rect 22100 28970 22152 28976
rect 22296 29022 22416 29050
rect 22112 28558 22140 28970
rect 22296 28558 22324 29022
rect 22376 28960 22428 28966
rect 22376 28902 22428 28908
rect 22100 28552 22152 28558
rect 22100 28494 22152 28500
rect 22284 28552 22336 28558
rect 22284 28494 22336 28500
rect 22192 28416 22244 28422
rect 22192 28358 22244 28364
rect 22204 28082 22232 28358
rect 22388 28082 22416 28902
rect 22664 28626 22692 29106
rect 22652 28620 22704 28626
rect 22652 28562 22704 28568
rect 22192 28076 22244 28082
rect 22192 28018 22244 28024
rect 22376 28076 22428 28082
rect 22376 28018 22428 28024
rect 22652 28076 22704 28082
rect 22652 28018 22704 28024
rect 22560 28008 22612 28014
rect 22560 27950 22612 27956
rect 22572 27538 22600 27950
rect 22560 27532 22612 27538
rect 22560 27474 22612 27480
rect 22468 26988 22520 26994
rect 22468 26930 22520 26936
rect 22284 26784 22336 26790
rect 22284 26726 22336 26732
rect 22296 26314 22324 26726
rect 22284 26308 22336 26314
rect 22284 26250 22336 26256
rect 22480 26042 22508 26930
rect 22560 26920 22612 26926
rect 22560 26862 22612 26868
rect 22468 26036 22520 26042
rect 22468 25978 22520 25984
rect 21916 25900 21968 25906
rect 21916 25842 21968 25848
rect 21928 25498 21956 25842
rect 22468 25696 22520 25702
rect 22468 25638 22520 25644
rect 21916 25492 21968 25498
rect 21916 25434 21968 25440
rect 21640 25152 21692 25158
rect 21640 25094 21692 25100
rect 21652 24954 21680 25094
rect 21640 24948 21692 24954
rect 21640 24890 21692 24896
rect 21928 23730 21956 25434
rect 22376 25288 22428 25294
rect 22376 25230 22428 25236
rect 22388 24818 22416 25230
rect 22100 24812 22152 24818
rect 22100 24754 22152 24760
rect 22376 24812 22428 24818
rect 22376 24754 22428 24760
rect 22008 24608 22060 24614
rect 22008 24550 22060 24556
rect 22020 24206 22048 24550
rect 22112 24274 22140 24754
rect 22480 24750 22508 25638
rect 22468 24744 22520 24750
rect 22468 24686 22520 24692
rect 22100 24268 22152 24274
rect 22100 24210 22152 24216
rect 22008 24200 22060 24206
rect 22008 24142 22060 24148
rect 21916 23724 21968 23730
rect 21916 23666 21968 23672
rect 22284 23520 22336 23526
rect 22284 23462 22336 23468
rect 21732 22568 21784 22574
rect 21732 22510 21784 22516
rect 21744 22438 21772 22510
rect 21732 22432 21784 22438
rect 21732 22374 21784 22380
rect 21744 22098 21772 22374
rect 21732 22092 21784 22098
rect 21732 22034 21784 22040
rect 21640 21888 21692 21894
rect 21640 21830 21692 21836
rect 21652 21690 21680 21830
rect 21640 21684 21692 21690
rect 21640 21626 21692 21632
rect 22100 20868 22152 20874
rect 22100 20810 22152 20816
rect 22112 20602 22140 20810
rect 22100 20596 22152 20602
rect 22100 20538 22152 20544
rect 22112 17678 22140 20538
rect 22192 19712 22244 19718
rect 22192 19654 22244 19660
rect 22204 18698 22232 19654
rect 22192 18692 22244 18698
rect 22192 18634 22244 18640
rect 22296 18290 22324 23462
rect 22376 21888 22428 21894
rect 22376 21830 22428 21836
rect 22388 21554 22416 21830
rect 22376 21548 22428 21554
rect 22376 21490 22428 21496
rect 22376 19848 22428 19854
rect 22376 19790 22428 19796
rect 22388 18426 22416 19790
rect 22468 19168 22520 19174
rect 22468 19110 22520 19116
rect 22376 18420 22428 18426
rect 22376 18362 22428 18368
rect 22284 18284 22336 18290
rect 22284 18226 22336 18232
rect 22100 17672 22152 17678
rect 22100 17614 22152 17620
rect 22192 17196 22244 17202
rect 22192 17138 22244 17144
rect 22100 17060 22152 17066
rect 22100 17002 22152 17008
rect 22008 16992 22060 16998
rect 22008 16934 22060 16940
rect 22020 16590 22048 16934
rect 22112 16794 22140 17002
rect 22100 16788 22152 16794
rect 22100 16730 22152 16736
rect 22008 16584 22060 16590
rect 22008 16526 22060 16532
rect 22112 15570 22140 16730
rect 22204 16250 22232 17138
rect 22192 16244 22244 16250
rect 22192 16186 22244 16192
rect 22296 16130 22324 18226
rect 22376 18216 22428 18222
rect 22480 18170 22508 19110
rect 22428 18164 22508 18170
rect 22376 18158 22508 18164
rect 22388 18142 22508 18158
rect 22204 16114 22324 16130
rect 22480 16114 22508 18142
rect 22572 17202 22600 26862
rect 22664 26586 22692 28018
rect 22652 26580 22704 26586
rect 22652 26522 22704 26528
rect 23112 26580 23164 26586
rect 23112 26522 23164 26528
rect 23124 25906 23152 26522
rect 23112 25900 23164 25906
rect 23112 25842 23164 25848
rect 23112 24812 23164 24818
rect 23112 24754 23164 24760
rect 23204 24812 23256 24818
rect 23204 24754 23256 24760
rect 22650 24440 22706 24449
rect 22650 24375 22706 24384
rect 23020 24404 23072 24410
rect 22664 23050 22692 24375
rect 23020 24346 23072 24352
rect 23032 23594 23060 24346
rect 23124 24206 23152 24754
rect 23216 24449 23244 24754
rect 23202 24440 23258 24449
rect 23202 24375 23204 24384
rect 23256 24375 23258 24384
rect 23204 24346 23256 24352
rect 23112 24200 23164 24206
rect 23112 24142 23164 24148
rect 23020 23588 23072 23594
rect 23020 23530 23072 23536
rect 22652 23044 22704 23050
rect 22652 22986 22704 22992
rect 22664 22574 22692 22986
rect 22928 22976 22980 22982
rect 22928 22918 22980 22924
rect 22940 22710 22968 22918
rect 22928 22704 22980 22710
rect 22928 22646 22980 22652
rect 22652 22568 22704 22574
rect 22652 22510 22704 22516
rect 23204 22568 23256 22574
rect 23204 22510 23256 22516
rect 23112 22160 23164 22166
rect 23112 22102 23164 22108
rect 22928 22092 22980 22098
rect 22928 22034 22980 22040
rect 22652 19848 22704 19854
rect 22652 19790 22704 19796
rect 22664 19310 22692 19790
rect 22940 19378 22968 22034
rect 23124 22030 23152 22102
rect 23216 22030 23244 22510
rect 23112 22024 23164 22030
rect 23112 21966 23164 21972
rect 23204 22024 23256 22030
rect 23204 21966 23256 21972
rect 23112 21344 23164 21350
rect 23112 21286 23164 21292
rect 23124 20754 23152 21286
rect 23204 20800 23256 20806
rect 23124 20748 23204 20754
rect 23124 20742 23256 20748
rect 23124 20726 23244 20742
rect 23124 19378 23152 20726
rect 22928 19372 22980 19378
rect 23112 19372 23164 19378
rect 22980 19332 23060 19360
rect 22928 19314 22980 19320
rect 22652 19304 22704 19310
rect 22652 19246 22704 19252
rect 22664 18154 22692 19246
rect 22928 18964 22980 18970
rect 22928 18906 22980 18912
rect 22744 18692 22796 18698
rect 22744 18634 22796 18640
rect 22756 18154 22784 18634
rect 22940 18290 22968 18906
rect 22928 18284 22980 18290
rect 22928 18226 22980 18232
rect 22652 18148 22704 18154
rect 22652 18090 22704 18096
rect 22744 18148 22796 18154
rect 22744 18090 22796 18096
rect 22652 17672 22704 17678
rect 22652 17614 22704 17620
rect 22560 17196 22612 17202
rect 22560 17138 22612 17144
rect 22560 16992 22612 16998
rect 22664 16980 22692 17614
rect 22756 17610 22784 18090
rect 22744 17604 22796 17610
rect 22744 17546 22796 17552
rect 22756 17066 22784 17546
rect 22744 17060 22796 17066
rect 22744 17002 22796 17008
rect 22612 16952 22692 16980
rect 22560 16934 22612 16940
rect 22192 16108 22324 16114
rect 22244 16102 22324 16108
rect 22468 16108 22520 16114
rect 22192 16050 22244 16056
rect 22468 16050 22520 16056
rect 22100 15564 22152 15570
rect 22100 15506 22152 15512
rect 21548 13524 21600 13530
rect 21548 13466 21600 13472
rect 20996 13252 21048 13258
rect 20996 13194 21048 13200
rect 22112 13190 22140 15506
rect 22204 13938 22232 16050
rect 22480 13938 22508 16050
rect 22572 14550 22600 16934
rect 22652 16448 22704 16454
rect 22652 16390 22704 16396
rect 22664 16114 22692 16390
rect 22652 16108 22704 16114
rect 22652 16050 22704 16056
rect 23032 15026 23060 19332
rect 23112 19314 23164 19320
rect 23020 15020 23072 15026
rect 23020 14962 23072 14968
rect 23032 14634 23060 14962
rect 23124 14958 23152 19314
rect 23204 15428 23256 15434
rect 23204 15370 23256 15376
rect 23112 14952 23164 14958
rect 23112 14894 23164 14900
rect 22940 14606 23060 14634
rect 22560 14544 22612 14550
rect 22560 14486 22612 14492
rect 22572 14006 22600 14486
rect 22560 14000 22612 14006
rect 22560 13942 22612 13948
rect 22192 13932 22244 13938
rect 22192 13874 22244 13880
rect 22468 13932 22520 13938
rect 22468 13874 22520 13880
rect 22652 13932 22704 13938
rect 22652 13874 22704 13880
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 22100 13184 22152 13190
rect 22100 13126 22152 13132
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 20732 12306 20760 13126
rect 22204 12850 22232 13874
rect 22480 13462 22508 13874
rect 22664 13530 22692 13874
rect 22652 13524 22704 13530
rect 22652 13466 22704 13472
rect 22468 13456 22520 13462
rect 22468 13398 22520 13404
rect 22940 13410 22968 14606
rect 23020 14544 23072 14550
rect 23020 14486 23072 14492
rect 23032 13530 23060 14486
rect 23020 13524 23072 13530
rect 23020 13466 23072 13472
rect 22480 12850 22508 13398
rect 22940 13382 23060 13410
rect 22836 13320 22888 13326
rect 22836 13262 22888 13268
rect 22928 13320 22980 13326
rect 22928 13262 22980 13268
rect 22652 13184 22704 13190
rect 22652 13126 22704 13132
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 22468 12844 22520 12850
rect 22468 12786 22520 12792
rect 20720 12300 20772 12306
rect 20720 12242 20772 12248
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 20732 11218 20760 12242
rect 22664 12238 22692 13126
rect 22848 12986 22876 13262
rect 22836 12980 22888 12986
rect 22836 12922 22888 12928
rect 22744 12844 22796 12850
rect 22744 12786 22796 12792
rect 22652 12232 22704 12238
rect 22652 12174 22704 12180
rect 22468 12164 22520 12170
rect 22468 12106 22520 12112
rect 22100 12096 22152 12102
rect 22100 12038 22152 12044
rect 22112 11898 22140 12038
rect 22100 11892 22152 11898
rect 22100 11834 22152 11840
rect 22480 11762 22508 12106
rect 22560 12096 22612 12102
rect 22560 12038 22612 12044
rect 22468 11756 22520 11762
rect 22468 11698 22520 11704
rect 20720 11212 20772 11218
rect 20720 11154 20772 11160
rect 21824 11212 21876 11218
rect 21824 11154 21876 11160
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 21836 10606 21864 11154
rect 22468 11076 22520 11082
rect 22468 11018 22520 11024
rect 22480 10810 22508 11018
rect 22468 10804 22520 10810
rect 22468 10746 22520 10752
rect 21824 10600 21876 10606
rect 21824 10542 21876 10548
rect 21836 10130 21864 10542
rect 21824 10124 21876 10130
rect 21824 10066 21876 10072
rect 22376 9988 22428 9994
rect 22376 9930 22428 9936
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 22388 9722 22416 9930
rect 22376 9716 22428 9722
rect 22376 9658 22428 9664
rect 22572 9586 22600 12038
rect 22756 11898 22784 12786
rect 22744 11892 22796 11898
rect 22744 11834 22796 11840
rect 22940 11762 22968 13262
rect 23032 12374 23060 13382
rect 23020 12368 23072 12374
rect 23020 12310 23072 12316
rect 23020 12232 23072 12238
rect 23124 12220 23152 14894
rect 23216 14618 23244 15370
rect 23204 14612 23256 14618
rect 23204 14554 23256 14560
rect 23308 13870 23336 29566
rect 23388 29572 23440 29578
rect 23388 29514 23440 29520
rect 23400 29170 23428 29514
rect 23492 29170 23520 29786
rect 23388 29164 23440 29170
rect 23388 29106 23440 29112
rect 23480 29164 23532 29170
rect 23480 29106 23532 29112
rect 23584 28762 23612 30262
rect 23664 29708 23716 29714
rect 23664 29650 23716 29656
rect 23676 29510 23704 29650
rect 23768 29646 23796 30330
rect 23756 29640 23808 29646
rect 23756 29582 23808 29588
rect 23664 29504 23716 29510
rect 23664 29446 23716 29452
rect 23676 29034 23704 29446
rect 23768 29170 23796 29582
rect 23756 29164 23808 29170
rect 23756 29106 23808 29112
rect 23664 29028 23716 29034
rect 23664 28970 23716 28976
rect 23572 28756 23624 28762
rect 23572 28698 23624 28704
rect 23676 28558 23704 28970
rect 23664 28552 23716 28558
rect 23664 28494 23716 28500
rect 23664 26852 23716 26858
rect 23664 26794 23716 26800
rect 23676 25838 23704 26794
rect 23756 25968 23808 25974
rect 23756 25910 23808 25916
rect 23664 25832 23716 25838
rect 23664 25774 23716 25780
rect 23676 25362 23704 25774
rect 23664 25356 23716 25362
rect 23664 25298 23716 25304
rect 23664 25220 23716 25226
rect 23664 25162 23716 25168
rect 23388 24608 23440 24614
rect 23388 24550 23440 24556
rect 23400 24342 23428 24550
rect 23676 24410 23704 25162
rect 23768 24818 23796 25910
rect 23756 24812 23808 24818
rect 23756 24754 23808 24760
rect 24216 24812 24268 24818
rect 24216 24754 24268 24760
rect 23664 24404 23716 24410
rect 23664 24346 23716 24352
rect 23388 24336 23440 24342
rect 23388 24278 23440 24284
rect 23400 24206 23428 24278
rect 23388 24200 23440 24206
rect 23388 24142 23440 24148
rect 23400 23526 23428 24142
rect 23480 24132 23532 24138
rect 23480 24074 23532 24080
rect 23388 23520 23440 23526
rect 23388 23462 23440 23468
rect 23400 23050 23428 23462
rect 23492 23322 23520 24074
rect 24228 23730 24256 24754
rect 24216 23724 24268 23730
rect 24216 23666 24268 23672
rect 23480 23316 23532 23322
rect 23480 23258 23532 23264
rect 23388 23044 23440 23050
rect 23388 22986 23440 22992
rect 23400 20942 23428 22986
rect 23492 22642 23520 23258
rect 23480 22636 23532 22642
rect 23480 22578 23532 22584
rect 23492 22250 23520 22578
rect 24228 22506 24256 23666
rect 24216 22500 24268 22506
rect 24216 22442 24268 22448
rect 23664 22432 23716 22438
rect 23664 22374 23716 22380
rect 23492 22222 23612 22250
rect 23584 22166 23612 22222
rect 23572 22160 23624 22166
rect 23572 22102 23624 22108
rect 23480 21888 23532 21894
rect 23480 21830 23532 21836
rect 23492 21078 23520 21830
rect 23480 21072 23532 21078
rect 23480 21014 23532 21020
rect 23388 20936 23440 20942
rect 23388 20878 23440 20884
rect 23400 20602 23428 20878
rect 23388 20596 23440 20602
rect 23388 20538 23440 20544
rect 23400 20466 23428 20538
rect 23492 20466 23520 21014
rect 23388 20460 23440 20466
rect 23388 20402 23440 20408
rect 23480 20460 23532 20466
rect 23480 20402 23532 20408
rect 23400 19990 23428 20402
rect 23388 19984 23440 19990
rect 23388 19926 23440 19932
rect 23492 19854 23520 20402
rect 23584 20262 23612 22102
rect 23676 21554 23704 22374
rect 23664 21548 23716 21554
rect 23664 21490 23716 21496
rect 23848 21548 23900 21554
rect 23848 21490 23900 21496
rect 23860 21010 23888 21490
rect 23848 21004 23900 21010
rect 23848 20946 23900 20952
rect 23756 20392 23808 20398
rect 23756 20334 23808 20340
rect 23572 20256 23624 20262
rect 23572 20198 23624 20204
rect 23572 20052 23624 20058
rect 23572 19994 23624 20000
rect 23480 19848 23532 19854
rect 23480 19790 23532 19796
rect 23584 18086 23612 19994
rect 23768 19174 23796 20334
rect 23756 19168 23808 19174
rect 23756 19110 23808 19116
rect 23572 18080 23624 18086
rect 23572 18022 23624 18028
rect 23584 17882 23612 18022
rect 23572 17876 23624 17882
rect 23572 17818 23624 17824
rect 23480 17264 23532 17270
rect 23480 17206 23532 17212
rect 23492 16794 23520 17206
rect 23848 17196 23900 17202
rect 23848 17138 23900 17144
rect 23480 16788 23532 16794
rect 23480 16730 23532 16736
rect 23664 15360 23716 15366
rect 23664 15302 23716 15308
rect 23388 14816 23440 14822
rect 23388 14758 23440 14764
rect 23400 14414 23428 14758
rect 23676 14482 23704 15302
rect 23860 15026 23888 17138
rect 23848 15020 23900 15026
rect 23848 14962 23900 14968
rect 23664 14476 23716 14482
rect 23664 14418 23716 14424
rect 23388 14408 23440 14414
rect 23388 14350 23440 14356
rect 23296 13864 23348 13870
rect 23296 13806 23348 13812
rect 23204 13388 23256 13394
rect 23204 13330 23256 13336
rect 23216 12918 23244 13330
rect 23204 12912 23256 12918
rect 23204 12854 23256 12860
rect 23308 12238 23336 13806
rect 23072 12192 23152 12220
rect 23296 12232 23348 12238
rect 23020 12174 23072 12180
rect 23296 12174 23348 12180
rect 23032 11830 23060 12174
rect 23020 11824 23072 11830
rect 23020 11766 23072 11772
rect 22928 11756 22980 11762
rect 22928 11698 22980 11704
rect 22652 11552 22704 11558
rect 22652 11494 22704 11500
rect 22664 10674 22692 11494
rect 23296 11348 23348 11354
rect 23296 11290 23348 11296
rect 23308 11014 23336 11290
rect 23296 11008 23348 11014
rect 23296 10950 23348 10956
rect 22652 10668 22704 10674
rect 22652 10610 22704 10616
rect 23308 10606 23336 10950
rect 23296 10600 23348 10606
rect 23296 10542 23348 10548
rect 22744 10464 22796 10470
rect 22744 10406 22796 10412
rect 22756 10180 22784 10406
rect 22836 10192 22888 10198
rect 22756 10152 22836 10180
rect 22756 9586 22784 10152
rect 22836 10134 22888 10140
rect 23204 9920 23256 9926
rect 23204 9862 23256 9868
rect 23216 9722 23244 9862
rect 23204 9716 23256 9722
rect 23204 9658 23256 9664
rect 23216 9586 23244 9658
rect 22560 9580 22612 9586
rect 22560 9522 22612 9528
rect 22744 9580 22796 9586
rect 22744 9522 22796 9528
rect 23204 9580 23256 9586
rect 23204 9522 23256 9528
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 18420 3392 18472 3398
rect 18420 3334 18472 3340
rect 17776 2576 17828 2582
rect 17776 2518 17828 2524
rect 18432 2446 18460 3334
rect 19444 3194 19472 4082
rect 19708 4072 19760 4078
rect 19708 4014 19760 4020
rect 22192 4072 22244 4078
rect 22192 4014 22244 4020
rect 22560 4072 22612 4078
rect 22560 4014 22612 4020
rect 19720 3602 19748 4014
rect 19892 3936 19944 3942
rect 19892 3878 19944 3884
rect 20168 3936 20220 3942
rect 20168 3878 20220 3884
rect 19904 3602 19932 3878
rect 19708 3596 19760 3602
rect 19708 3538 19760 3544
rect 19892 3596 19944 3602
rect 19892 3538 19944 3544
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19432 3188 19484 3194
rect 19432 3130 19484 3136
rect 18512 2984 18564 2990
rect 18512 2926 18564 2932
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 18524 2650 18552 2926
rect 18512 2644 18564 2650
rect 18512 2586 18564 2592
rect 18420 2440 18472 2446
rect 18420 2382 18472 2388
rect 17500 2032 17552 2038
rect 17500 1974 17552 1980
rect 19352 800 19380 2926
rect 19444 2446 19472 3130
rect 20180 3126 20208 3878
rect 22204 3738 22232 4014
rect 22008 3732 22060 3738
rect 22008 3674 22060 3680
rect 22192 3732 22244 3738
rect 22192 3674 22244 3680
rect 22284 3732 22336 3738
rect 22284 3674 22336 3680
rect 22020 3618 22048 3674
rect 22296 3618 22324 3674
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 22020 3590 22324 3618
rect 20168 3120 20220 3126
rect 20168 3062 20220 3068
rect 19800 2984 19852 2990
rect 19800 2926 19852 2932
rect 19812 2650 19840 2926
rect 19800 2644 19852 2650
rect 19800 2586 19852 2592
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19996 800 20024 2382
rect 20640 800 20668 3538
rect 22020 3534 22048 3590
rect 22008 3528 22060 3534
rect 22008 3470 22060 3476
rect 22572 800 22600 4014
rect 23860 2310 23888 14962
rect 24320 12306 24348 31726
rect 24596 29714 24624 31826
rect 24860 31340 24912 31346
rect 24964 31328 24992 31962
rect 24912 31300 24992 31328
rect 24860 31282 24912 31288
rect 24768 31136 24820 31142
rect 24768 31078 24820 31084
rect 24584 29708 24636 29714
rect 24412 29668 24584 29696
rect 24412 29238 24440 29668
rect 24584 29650 24636 29656
rect 24676 29572 24728 29578
rect 24676 29514 24728 29520
rect 24688 29306 24716 29514
rect 24676 29300 24728 29306
rect 24676 29242 24728 29248
rect 24400 29232 24452 29238
rect 24400 29174 24452 29180
rect 24584 28076 24636 28082
rect 24584 28018 24636 28024
rect 24596 27130 24624 28018
rect 24780 27878 24808 31078
rect 24872 28098 24900 31282
rect 25148 30326 25176 34546
rect 25228 32428 25280 32434
rect 25228 32370 25280 32376
rect 25240 31686 25268 32370
rect 25320 32020 25372 32026
rect 25320 31962 25372 31968
rect 25228 31680 25280 31686
rect 25228 31622 25280 31628
rect 25240 31278 25268 31622
rect 25332 31346 25360 31962
rect 25320 31340 25372 31346
rect 25320 31282 25372 31288
rect 25228 31272 25280 31278
rect 25228 31214 25280 31220
rect 25136 30320 25188 30326
rect 25136 30262 25188 30268
rect 24952 29504 25004 29510
rect 24952 29446 25004 29452
rect 24964 28626 24992 29446
rect 25044 29232 25096 29238
rect 25044 29174 25096 29180
rect 24952 28620 25004 28626
rect 24952 28562 25004 28568
rect 24872 28070 24992 28098
rect 24768 27872 24820 27878
rect 24768 27814 24820 27820
rect 24860 27872 24912 27878
rect 24860 27814 24912 27820
rect 24584 27124 24636 27130
rect 24584 27066 24636 27072
rect 24676 26988 24728 26994
rect 24676 26930 24728 26936
rect 24584 26784 24636 26790
rect 24584 26726 24636 26732
rect 24596 25226 24624 26726
rect 24688 26382 24716 26930
rect 24780 26790 24808 27814
rect 24872 27402 24900 27814
rect 24860 27396 24912 27402
rect 24860 27338 24912 27344
rect 24964 26926 24992 28070
rect 25056 27334 25084 29174
rect 25044 27328 25096 27334
rect 25044 27270 25096 27276
rect 25056 26994 25084 27270
rect 25240 27062 25268 31214
rect 25412 28960 25464 28966
rect 25412 28902 25464 28908
rect 25424 28014 25452 28902
rect 25412 28008 25464 28014
rect 25412 27950 25464 27956
rect 25228 27056 25280 27062
rect 25228 26998 25280 27004
rect 25044 26988 25096 26994
rect 25044 26930 25096 26936
rect 24952 26920 25004 26926
rect 24952 26862 25004 26868
rect 24768 26784 24820 26790
rect 24768 26726 24820 26732
rect 24676 26376 24728 26382
rect 24676 26318 24728 26324
rect 24688 25974 24716 26318
rect 24676 25968 24728 25974
rect 24676 25910 24728 25916
rect 24964 25498 24992 26862
rect 25136 26784 25188 26790
rect 25136 26726 25188 26732
rect 25148 26586 25176 26726
rect 25136 26580 25188 26586
rect 25136 26522 25188 26528
rect 25148 26314 25176 26522
rect 25136 26308 25188 26314
rect 25136 26250 25188 26256
rect 25044 26240 25096 26246
rect 25044 26182 25096 26188
rect 25056 25770 25084 26182
rect 25044 25764 25096 25770
rect 25044 25706 25096 25712
rect 24952 25492 25004 25498
rect 24952 25434 25004 25440
rect 24584 25220 24636 25226
rect 24584 25162 24636 25168
rect 24400 24744 24452 24750
rect 24400 24686 24452 24692
rect 24412 24070 24440 24686
rect 24596 24290 24624 25162
rect 24768 24676 24820 24682
rect 24768 24618 24820 24624
rect 24676 24608 24728 24614
rect 24676 24550 24728 24556
rect 24504 24274 24624 24290
rect 24492 24268 24624 24274
rect 24544 24262 24624 24268
rect 24492 24210 24544 24216
rect 24400 24064 24452 24070
rect 24400 24006 24452 24012
rect 24412 23798 24440 24006
rect 24400 23792 24452 23798
rect 24400 23734 24452 23740
rect 24412 22438 24440 23734
rect 24596 23322 24624 24262
rect 24584 23316 24636 23322
rect 24584 23258 24636 23264
rect 24688 23118 24716 24550
rect 24780 24138 24808 24618
rect 24768 24132 24820 24138
rect 24768 24074 24820 24080
rect 24780 23526 24808 24074
rect 25056 23866 25084 25706
rect 25044 23860 25096 23866
rect 25044 23802 25096 23808
rect 24768 23520 24820 23526
rect 24768 23462 24820 23468
rect 24676 23112 24728 23118
rect 24676 23054 24728 23060
rect 24400 22432 24452 22438
rect 24400 22374 24452 22380
rect 24412 20942 24440 22374
rect 24492 22024 24544 22030
rect 24492 21966 24544 21972
rect 25044 22024 25096 22030
rect 25044 21966 25096 21972
rect 24400 20936 24452 20942
rect 24400 20878 24452 20884
rect 24412 20534 24440 20878
rect 24400 20528 24452 20534
rect 24400 20470 24452 20476
rect 24400 17196 24452 17202
rect 24400 17138 24452 17144
rect 24412 16998 24440 17138
rect 24400 16992 24452 16998
rect 24400 16934 24452 16940
rect 24412 16114 24440 16934
rect 24504 16658 24532 21966
rect 24584 21888 24636 21894
rect 24584 21830 24636 21836
rect 24596 21622 24624 21830
rect 24584 21616 24636 21622
rect 24584 21558 24636 21564
rect 25056 21146 25084 21966
rect 25228 21480 25280 21486
rect 25228 21422 25280 21428
rect 25044 21140 25096 21146
rect 25044 21082 25096 21088
rect 24860 20256 24912 20262
rect 24860 20198 24912 20204
rect 24768 19440 24820 19446
rect 24768 19382 24820 19388
rect 24676 19168 24728 19174
rect 24676 19110 24728 19116
rect 24688 18902 24716 19110
rect 24676 18896 24728 18902
rect 24676 18838 24728 18844
rect 24780 18766 24808 19382
rect 24872 19378 24900 20198
rect 25136 19780 25188 19786
rect 25136 19722 25188 19728
rect 24860 19372 24912 19378
rect 24912 19332 25084 19360
rect 24860 19314 24912 19320
rect 24768 18760 24820 18766
rect 24768 18702 24820 18708
rect 24584 18624 24636 18630
rect 24584 18566 24636 18572
rect 24596 18358 24624 18566
rect 24584 18352 24636 18358
rect 24584 18294 24636 18300
rect 24860 16992 24912 16998
rect 24860 16934 24912 16940
rect 24492 16652 24544 16658
rect 24492 16594 24544 16600
rect 24872 16590 24900 16934
rect 24860 16584 24912 16590
rect 24860 16526 24912 16532
rect 24952 16448 25004 16454
rect 24952 16390 25004 16396
rect 24964 16182 24992 16390
rect 24952 16176 25004 16182
rect 24952 16118 25004 16124
rect 24400 16108 24452 16114
rect 24400 16050 24452 16056
rect 24584 16108 24636 16114
rect 24584 16050 24636 16056
rect 24768 16108 24820 16114
rect 24768 16050 24820 16056
rect 24596 15502 24624 16050
rect 24780 15978 24808 16050
rect 24768 15972 24820 15978
rect 24768 15914 24820 15920
rect 24780 15570 24808 15914
rect 24768 15564 24820 15570
rect 24768 15506 24820 15512
rect 24584 15496 24636 15502
rect 24584 15438 24636 15444
rect 24596 15366 24624 15438
rect 24584 15360 24636 15366
rect 24584 15302 24636 15308
rect 25056 14618 25084 19332
rect 25148 17678 25176 19722
rect 25136 17672 25188 17678
rect 25136 17614 25188 17620
rect 25240 16658 25268 21422
rect 25320 17128 25372 17134
rect 25320 17070 25372 17076
rect 25228 16652 25280 16658
rect 25228 16594 25280 16600
rect 25332 16522 25360 17070
rect 25320 16516 25372 16522
rect 25320 16458 25372 16464
rect 25044 14612 25096 14618
rect 25044 14554 25096 14560
rect 24860 14408 24912 14414
rect 24860 14350 24912 14356
rect 24584 14272 24636 14278
rect 24584 14214 24636 14220
rect 24596 13938 24624 14214
rect 24584 13932 24636 13938
rect 24584 13874 24636 13880
rect 24872 13530 24900 14350
rect 24860 13524 24912 13530
rect 24860 13466 24912 13472
rect 24952 13320 25004 13326
rect 24952 13262 25004 13268
rect 24860 13252 24912 13258
rect 24860 13194 24912 13200
rect 24308 12300 24360 12306
rect 24308 12242 24360 12248
rect 24872 12170 24900 13194
rect 24964 12238 24992 13262
rect 24952 12232 25004 12238
rect 24952 12174 25004 12180
rect 24860 12164 24912 12170
rect 24860 12106 24912 12112
rect 24872 11830 24900 12106
rect 24860 11824 24912 11830
rect 24860 11766 24912 11772
rect 24860 11688 24912 11694
rect 24964 11676 24992 12174
rect 24912 11648 24992 11676
rect 24860 11630 24912 11636
rect 25056 11626 25084 14554
rect 25424 13326 25452 27950
rect 25516 26586 25544 36722
rect 25608 32978 25636 38406
rect 25964 38344 26016 38350
rect 25964 38286 26016 38292
rect 25780 37868 25832 37874
rect 25780 37810 25832 37816
rect 25792 37330 25820 37810
rect 25780 37324 25832 37330
rect 25780 37266 25832 37272
rect 25792 36786 25820 37266
rect 25872 37256 25924 37262
rect 25872 37198 25924 37204
rect 25780 36780 25832 36786
rect 25780 36722 25832 36728
rect 25792 36378 25820 36722
rect 25884 36718 25912 37198
rect 25872 36712 25924 36718
rect 25872 36654 25924 36660
rect 25780 36372 25832 36378
rect 25780 36314 25832 36320
rect 25884 36242 25912 36654
rect 25872 36236 25924 36242
rect 25872 36178 25924 36184
rect 25688 36168 25740 36174
rect 25688 36110 25740 36116
rect 25700 34746 25728 36110
rect 25688 34740 25740 34746
rect 25688 34682 25740 34688
rect 25976 34626 26004 38286
rect 26068 37942 26096 38814
rect 26148 38752 26200 38758
rect 26148 38694 26200 38700
rect 26160 38486 26188 38694
rect 26148 38480 26200 38486
rect 26148 38422 26200 38428
rect 26056 37936 26108 37942
rect 26056 37878 26108 37884
rect 26160 37874 26188 38422
rect 27080 38214 27108 38830
rect 27540 38418 27568 39986
rect 27816 39438 27844 40122
rect 28460 39846 28488 40394
rect 28540 40384 28592 40390
rect 28540 40326 28592 40332
rect 28552 40118 28580 40326
rect 28540 40112 28592 40118
rect 28540 40054 28592 40060
rect 28448 39840 28500 39846
rect 28448 39782 28500 39788
rect 27804 39432 27856 39438
rect 27804 39374 27856 39380
rect 27528 38412 27580 38418
rect 27528 38354 27580 38360
rect 28264 38344 28316 38350
rect 28264 38286 28316 38292
rect 27252 38276 27304 38282
rect 27252 38218 27304 38224
rect 27712 38276 27764 38282
rect 27712 38218 27764 38224
rect 27068 38208 27120 38214
rect 27068 38150 27120 38156
rect 26148 37868 26200 37874
rect 26148 37810 26200 37816
rect 27080 37806 27108 38150
rect 27068 37800 27120 37806
rect 27068 37742 27120 37748
rect 26424 37664 26476 37670
rect 26424 37606 26476 37612
rect 26436 37330 26464 37606
rect 26424 37324 26476 37330
rect 26424 37266 26476 37272
rect 26436 36854 26464 37266
rect 26884 37188 26936 37194
rect 26884 37130 26936 37136
rect 26896 36922 26924 37130
rect 26884 36916 26936 36922
rect 26884 36858 26936 36864
rect 26424 36848 26476 36854
rect 26424 36790 26476 36796
rect 27080 36786 27108 37742
rect 27264 37466 27292 38218
rect 27620 38208 27672 38214
rect 27620 38150 27672 38156
rect 27632 37942 27660 38150
rect 27620 37936 27672 37942
rect 27620 37878 27672 37884
rect 27252 37460 27304 37466
rect 27252 37402 27304 37408
rect 27724 37262 27752 38218
rect 27896 37868 27948 37874
rect 27896 37810 27948 37816
rect 27908 37466 27936 37810
rect 27896 37460 27948 37466
rect 27896 37402 27948 37408
rect 28276 37330 28304 38286
rect 28264 37324 28316 37330
rect 28264 37266 28316 37272
rect 27712 37256 27764 37262
rect 27712 37198 27764 37204
rect 27068 36780 27120 36786
rect 27068 36722 27120 36728
rect 26332 36168 26384 36174
rect 26332 36110 26384 36116
rect 26424 36168 26476 36174
rect 26424 36110 26476 36116
rect 26884 36168 26936 36174
rect 26884 36110 26936 36116
rect 26344 35766 26372 36110
rect 26332 35760 26384 35766
rect 26332 35702 26384 35708
rect 26344 35290 26372 35702
rect 26436 35698 26464 36110
rect 26700 36100 26752 36106
rect 26700 36042 26752 36048
rect 26424 35692 26476 35698
rect 26424 35634 26476 35640
rect 26332 35284 26384 35290
rect 26332 35226 26384 35232
rect 26424 35012 26476 35018
rect 26424 34954 26476 34960
rect 25884 34598 26004 34626
rect 25884 34474 25912 34598
rect 25964 34536 26016 34542
rect 25964 34478 26016 34484
rect 26332 34536 26384 34542
rect 26332 34478 26384 34484
rect 25872 34468 25924 34474
rect 25872 34410 25924 34416
rect 25596 32972 25648 32978
rect 25596 32914 25648 32920
rect 25976 32026 26004 34478
rect 26344 33114 26372 34478
rect 26332 33108 26384 33114
rect 26332 33050 26384 33056
rect 26240 32496 26292 32502
rect 26240 32438 26292 32444
rect 25964 32020 26016 32026
rect 25964 31962 26016 31968
rect 26252 30258 26280 32438
rect 26344 32434 26372 33050
rect 26436 32570 26464 34954
rect 26712 34610 26740 36042
rect 26896 35834 26924 36110
rect 26884 35828 26936 35834
rect 26884 35770 26936 35776
rect 27080 35086 27108 36722
rect 28276 36258 28304 37266
rect 28276 36230 28396 36258
rect 28264 36168 28316 36174
rect 28264 36110 28316 36116
rect 27620 36100 27672 36106
rect 27620 36042 27672 36048
rect 27436 35692 27488 35698
rect 27436 35634 27488 35640
rect 27068 35080 27120 35086
rect 27068 35022 27120 35028
rect 27160 35080 27212 35086
rect 27160 35022 27212 35028
rect 26976 34944 27028 34950
rect 26976 34886 27028 34892
rect 26988 34678 27016 34886
rect 26976 34672 27028 34678
rect 26976 34614 27028 34620
rect 27080 34610 27108 35022
rect 26700 34604 26752 34610
rect 26700 34546 26752 34552
rect 27068 34604 27120 34610
rect 27068 34546 27120 34552
rect 26424 32564 26476 32570
rect 26424 32506 26476 32512
rect 26332 32428 26384 32434
rect 26332 32370 26384 32376
rect 26608 30320 26660 30326
rect 26608 30262 26660 30268
rect 25688 30252 25740 30258
rect 25688 30194 25740 30200
rect 26240 30252 26292 30258
rect 26240 30194 26292 30200
rect 26516 30252 26568 30258
rect 26516 30194 26568 30200
rect 25596 26920 25648 26926
rect 25596 26862 25648 26868
rect 25504 26580 25556 26586
rect 25504 26522 25556 26528
rect 25608 26382 25636 26862
rect 25700 26518 25728 30194
rect 26148 29572 26200 29578
rect 26148 29514 26200 29520
rect 26160 29306 26188 29514
rect 26148 29300 26200 29306
rect 26148 29242 26200 29248
rect 26252 27554 26280 30194
rect 26332 30048 26384 30054
rect 26332 29990 26384 29996
rect 26344 29170 26372 29990
rect 26528 29510 26556 30194
rect 26516 29504 26568 29510
rect 26516 29446 26568 29452
rect 26332 29164 26384 29170
rect 26332 29106 26384 29112
rect 26620 27606 26648 30262
rect 26712 28966 26740 34546
rect 27172 34202 27200 35022
rect 27160 34196 27212 34202
rect 27160 34138 27212 34144
rect 26884 33992 26936 33998
rect 26884 33934 26936 33940
rect 26896 31822 26924 33934
rect 27068 33924 27120 33930
rect 27068 33866 27120 33872
rect 27080 33046 27108 33866
rect 27068 33040 27120 33046
rect 27068 32982 27120 32988
rect 27080 31890 27108 32982
rect 27252 32428 27304 32434
rect 27252 32370 27304 32376
rect 27068 31884 27120 31890
rect 27068 31826 27120 31832
rect 26884 31816 26936 31822
rect 26884 31758 26936 31764
rect 26792 31680 26844 31686
rect 26792 31622 26844 31628
rect 26804 31346 26832 31622
rect 26792 31340 26844 31346
rect 26792 31282 26844 31288
rect 26700 28960 26752 28966
rect 26700 28902 26752 28908
rect 26712 28082 26740 28902
rect 26700 28076 26752 28082
rect 26700 28018 26752 28024
rect 26608 27600 26660 27606
rect 26252 27526 26372 27554
rect 26608 27542 26660 27548
rect 26240 27396 26292 27402
rect 26240 27338 26292 27344
rect 25872 26988 25924 26994
rect 25872 26930 25924 26936
rect 25780 26784 25832 26790
rect 25780 26726 25832 26732
rect 25688 26512 25740 26518
rect 25688 26454 25740 26460
rect 25700 26382 25728 26454
rect 25596 26376 25648 26382
rect 25596 26318 25648 26324
rect 25688 26376 25740 26382
rect 25688 26318 25740 26324
rect 25608 25888 25636 26318
rect 25700 26042 25728 26318
rect 25688 26036 25740 26042
rect 25688 25978 25740 25984
rect 25688 25900 25740 25906
rect 25608 25860 25688 25888
rect 25688 25842 25740 25848
rect 25700 25294 25728 25842
rect 25688 25288 25740 25294
rect 25688 25230 25740 25236
rect 25688 24812 25740 24818
rect 25688 24754 25740 24760
rect 25596 24336 25648 24342
rect 25596 24278 25648 24284
rect 25608 23730 25636 24278
rect 25700 23866 25728 24754
rect 25792 24138 25820 26726
rect 25884 25974 25912 26930
rect 26252 26450 26280 27338
rect 26344 26518 26372 27526
rect 26424 27464 26476 27470
rect 26424 27406 26476 27412
rect 26332 26512 26384 26518
rect 26332 26454 26384 26460
rect 26240 26444 26292 26450
rect 26240 26386 26292 26392
rect 25872 25968 25924 25974
rect 25872 25910 25924 25916
rect 25884 24818 25912 25910
rect 25872 24812 25924 24818
rect 25872 24754 25924 24760
rect 25884 24138 25912 24754
rect 26252 24614 26280 26386
rect 26436 26042 26464 27406
rect 26712 27062 26740 28018
rect 26700 27056 26752 27062
rect 26700 26998 26752 27004
rect 27080 26314 27108 31826
rect 27264 31482 27292 32370
rect 27448 32230 27476 35634
rect 27528 35148 27580 35154
rect 27632 35136 27660 36042
rect 27896 35216 27948 35222
rect 27896 35158 27948 35164
rect 27580 35108 27660 35136
rect 27528 35090 27580 35096
rect 27436 32224 27488 32230
rect 27436 32166 27488 32172
rect 27448 31822 27476 32166
rect 27436 31816 27488 31822
rect 27436 31758 27488 31764
rect 27252 31476 27304 31482
rect 27252 31418 27304 31424
rect 27540 31142 27568 35090
rect 27804 32020 27856 32026
rect 27804 31962 27856 31968
rect 27816 31278 27844 31962
rect 27804 31272 27856 31278
rect 27804 31214 27856 31220
rect 27528 31136 27580 31142
rect 27528 31078 27580 31084
rect 27540 29170 27568 31078
rect 27620 29572 27672 29578
rect 27620 29514 27672 29520
rect 27528 29164 27580 29170
rect 27528 29106 27580 29112
rect 27632 28762 27660 29514
rect 27712 28960 27764 28966
rect 27712 28902 27764 28908
rect 27620 28756 27672 28762
rect 27620 28698 27672 28704
rect 27160 28620 27212 28626
rect 27160 28562 27212 28568
rect 27172 27402 27200 28562
rect 27724 28558 27752 28902
rect 27712 28552 27764 28558
rect 27712 28494 27764 28500
rect 27160 27396 27212 27402
rect 27160 27338 27212 27344
rect 27172 26994 27200 27338
rect 27160 26988 27212 26994
rect 27160 26930 27212 26936
rect 27252 26988 27304 26994
rect 27252 26930 27304 26936
rect 27068 26308 27120 26314
rect 27068 26250 27120 26256
rect 27264 26042 27292 26930
rect 27344 26240 27396 26246
rect 27344 26182 27396 26188
rect 26424 26036 26476 26042
rect 26424 25978 26476 25984
rect 27252 26036 27304 26042
rect 27252 25978 27304 25984
rect 27356 25906 27384 26182
rect 27344 25900 27396 25906
rect 27344 25842 27396 25848
rect 27528 25696 27580 25702
rect 27528 25638 27580 25644
rect 27540 25430 27568 25638
rect 27528 25424 27580 25430
rect 27528 25366 27580 25372
rect 27712 25288 27764 25294
rect 27712 25230 27764 25236
rect 27528 24812 27580 24818
rect 27528 24754 27580 24760
rect 27620 24812 27672 24818
rect 27620 24754 27672 24760
rect 26240 24608 26292 24614
rect 26240 24550 26292 24556
rect 27160 24608 27212 24614
rect 27160 24550 27212 24556
rect 26252 24274 26280 24550
rect 26240 24268 26292 24274
rect 26240 24210 26292 24216
rect 27172 24206 27200 24550
rect 27160 24200 27212 24206
rect 27160 24142 27212 24148
rect 25780 24132 25832 24138
rect 25780 24074 25832 24080
rect 25872 24132 25924 24138
rect 25872 24074 25924 24080
rect 27540 23866 27568 24754
rect 25688 23860 25740 23866
rect 25688 23802 25740 23808
rect 27528 23860 27580 23866
rect 27528 23802 27580 23808
rect 25596 23724 25648 23730
rect 25596 23666 25648 23672
rect 25780 23724 25832 23730
rect 25780 23666 25832 23672
rect 25792 23526 25820 23666
rect 26700 23656 26752 23662
rect 26700 23598 26752 23604
rect 25780 23520 25832 23526
rect 25780 23462 25832 23468
rect 25792 22094 25820 23462
rect 26240 23112 26292 23118
rect 26240 23054 26292 23060
rect 25608 22066 25820 22094
rect 25608 21962 25636 22066
rect 26252 21962 26280 23054
rect 26712 22030 26740 23598
rect 27632 22030 27660 24754
rect 27724 23118 27752 25230
rect 27712 23112 27764 23118
rect 27712 23054 27764 23060
rect 27712 22976 27764 22982
rect 27712 22918 27764 22924
rect 27724 22778 27752 22918
rect 27712 22772 27764 22778
rect 27712 22714 27764 22720
rect 26700 22024 26752 22030
rect 26700 21966 26752 21972
rect 27620 22024 27672 22030
rect 27620 21966 27672 21972
rect 25596 21956 25648 21962
rect 25596 21898 25648 21904
rect 25872 21956 25924 21962
rect 25872 21898 25924 21904
rect 26240 21956 26292 21962
rect 26240 21898 26292 21904
rect 27160 21956 27212 21962
rect 27160 21898 27212 21904
rect 25884 21690 25912 21898
rect 26148 21888 26200 21894
rect 26148 21830 26200 21836
rect 25872 21684 25924 21690
rect 25872 21626 25924 21632
rect 25884 21554 25912 21626
rect 25872 21548 25924 21554
rect 25872 21490 25924 21496
rect 25884 20942 25912 21490
rect 26160 20942 26188 21830
rect 26252 21554 26280 21898
rect 26240 21548 26292 21554
rect 26240 21490 26292 21496
rect 27172 21146 27200 21898
rect 27344 21888 27396 21894
rect 27344 21830 27396 21836
rect 27252 21548 27304 21554
rect 27252 21490 27304 21496
rect 27160 21140 27212 21146
rect 27160 21082 27212 21088
rect 25872 20936 25924 20942
rect 25872 20878 25924 20884
rect 26148 20936 26200 20942
rect 26148 20878 26200 20884
rect 26700 20800 26752 20806
rect 26700 20742 26752 20748
rect 26240 20256 26292 20262
rect 26240 20198 26292 20204
rect 26252 18986 26280 20198
rect 26424 19508 26476 19514
rect 26424 19450 26476 19456
rect 26332 19236 26384 19242
rect 26332 19178 26384 19184
rect 25976 18958 26280 18986
rect 25976 18902 26004 18958
rect 25964 18896 26016 18902
rect 25964 18838 26016 18844
rect 26344 18834 26372 19178
rect 26436 18902 26464 19450
rect 26424 18896 26476 18902
rect 26424 18838 26476 18844
rect 26332 18828 26384 18834
rect 26332 18770 26384 18776
rect 26240 18760 26292 18766
rect 26240 18702 26292 18708
rect 26252 17338 26280 18702
rect 26344 18290 26372 18770
rect 26608 18624 26660 18630
rect 26608 18566 26660 18572
rect 26620 18290 26648 18566
rect 26332 18284 26384 18290
rect 26332 18226 26384 18232
rect 26608 18284 26660 18290
rect 26608 18226 26660 18232
rect 26240 17332 26292 17338
rect 26240 17274 26292 17280
rect 26148 17196 26200 17202
rect 26148 17138 26200 17144
rect 26160 16794 26188 17138
rect 26252 17066 26280 17274
rect 26240 17060 26292 17066
rect 26240 17002 26292 17008
rect 26148 16788 26200 16794
rect 26148 16730 26200 16736
rect 26332 16720 26384 16726
rect 26332 16662 26384 16668
rect 25780 16652 25832 16658
rect 25780 16594 25832 16600
rect 25964 16652 26016 16658
rect 25964 16594 26016 16600
rect 25688 14408 25740 14414
rect 25688 14350 25740 14356
rect 25700 14074 25728 14350
rect 25688 14068 25740 14074
rect 25688 14010 25740 14016
rect 25792 13938 25820 16594
rect 25976 16046 26004 16594
rect 26056 16516 26108 16522
rect 26056 16458 26108 16464
rect 25964 16040 26016 16046
rect 25964 15982 26016 15988
rect 25780 13932 25832 13938
rect 25780 13874 25832 13880
rect 25412 13320 25464 13326
rect 25412 13262 25464 13268
rect 25596 12096 25648 12102
rect 25596 12038 25648 12044
rect 25608 11762 25636 12038
rect 25872 11824 25924 11830
rect 25872 11766 25924 11772
rect 25136 11756 25188 11762
rect 25136 11698 25188 11704
rect 25596 11756 25648 11762
rect 25596 11698 25648 11704
rect 25044 11620 25096 11626
rect 25044 11562 25096 11568
rect 24768 11552 24820 11558
rect 24768 11494 24820 11500
rect 24584 10668 24636 10674
rect 24584 10610 24636 10616
rect 24596 10266 24624 10610
rect 24584 10260 24636 10266
rect 24584 10202 24636 10208
rect 24780 10062 24808 11494
rect 25044 10736 25096 10742
rect 25044 10678 25096 10684
rect 25056 10130 25084 10678
rect 25044 10124 25096 10130
rect 25044 10066 25096 10072
rect 24768 10056 24820 10062
rect 24768 9998 24820 10004
rect 24768 3936 24820 3942
rect 24768 3878 24820 3884
rect 24780 3058 24808 3878
rect 24952 3392 25004 3398
rect 24952 3334 25004 3340
rect 24964 3126 24992 3334
rect 24952 3120 25004 3126
rect 24952 3062 25004 3068
rect 24768 3052 24820 3058
rect 24768 2994 24820 3000
rect 25148 2774 25176 11698
rect 25884 11558 25912 11766
rect 25964 11620 26016 11626
rect 25964 11562 26016 11568
rect 25412 11552 25464 11558
rect 25412 11494 25464 11500
rect 25780 11552 25832 11558
rect 25780 11494 25832 11500
rect 25872 11552 25924 11558
rect 25872 11494 25924 11500
rect 25424 11082 25452 11494
rect 25412 11076 25464 11082
rect 25412 11018 25464 11024
rect 25792 10198 25820 11494
rect 25976 11286 26004 11562
rect 25964 11280 26016 11286
rect 25964 11222 26016 11228
rect 25780 10192 25832 10198
rect 25780 10134 25832 10140
rect 25964 3936 26016 3942
rect 25964 3878 26016 3884
rect 25976 3602 26004 3878
rect 25964 3596 26016 3602
rect 25964 3538 26016 3544
rect 25320 3528 25372 3534
rect 25320 3470 25372 3476
rect 25056 2746 25176 2774
rect 25056 2582 25084 2746
rect 25044 2576 25096 2582
rect 25044 2518 25096 2524
rect 25332 2378 25360 3470
rect 25780 2984 25832 2990
rect 25780 2926 25832 2932
rect 25320 2372 25372 2378
rect 25320 2314 25372 2320
rect 23848 2304 23900 2310
rect 23848 2246 23900 2252
rect 25792 800 25820 2926
rect 26068 2514 26096 16458
rect 26344 16250 26372 16662
rect 26712 16590 26740 20742
rect 27264 20602 27292 21490
rect 27252 20596 27304 20602
rect 27252 20538 27304 20544
rect 27356 20466 27384 21830
rect 27344 20460 27396 20466
rect 27344 20402 27396 20408
rect 26792 19372 26844 19378
rect 26792 19314 26844 19320
rect 27344 19372 27396 19378
rect 27344 19314 27396 19320
rect 26804 18970 26832 19314
rect 27068 19168 27120 19174
rect 27068 19110 27120 19116
rect 26792 18964 26844 18970
rect 26792 18906 26844 18912
rect 27080 18902 27108 19110
rect 27068 18896 27120 18902
rect 27068 18838 27120 18844
rect 27252 18692 27304 18698
rect 27252 18634 27304 18640
rect 27264 18358 27292 18634
rect 27252 18352 27304 18358
rect 27252 18294 27304 18300
rect 27356 18290 27384 19314
rect 27712 19236 27764 19242
rect 27712 19178 27764 19184
rect 27528 19168 27580 19174
rect 27528 19110 27580 19116
rect 27540 18970 27568 19110
rect 27528 18964 27580 18970
rect 27528 18906 27580 18912
rect 27540 18766 27568 18906
rect 27528 18760 27580 18766
rect 27528 18702 27580 18708
rect 27436 18624 27488 18630
rect 27436 18566 27488 18572
rect 27344 18284 27396 18290
rect 27344 18226 27396 18232
rect 27448 18170 27476 18566
rect 27540 18358 27568 18702
rect 27528 18352 27580 18358
rect 27528 18294 27580 18300
rect 27724 18290 27752 19178
rect 27712 18284 27764 18290
rect 27712 18226 27764 18232
rect 27528 18216 27580 18222
rect 27448 18164 27528 18170
rect 27448 18158 27580 18164
rect 27448 18142 27568 18158
rect 27252 18080 27304 18086
rect 27252 18022 27304 18028
rect 27264 16590 27292 18022
rect 27436 17060 27488 17066
rect 27436 17002 27488 17008
rect 26700 16584 26752 16590
rect 26700 16526 26752 16532
rect 27068 16584 27120 16590
rect 27068 16526 27120 16532
rect 27252 16584 27304 16590
rect 27252 16526 27304 16532
rect 27344 16584 27396 16590
rect 27344 16526 27396 16532
rect 26424 16516 26476 16522
rect 26424 16458 26476 16464
rect 26516 16516 26568 16522
rect 26516 16458 26568 16464
rect 26436 16250 26464 16458
rect 26332 16244 26384 16250
rect 26332 16186 26384 16192
rect 26424 16244 26476 16250
rect 26424 16186 26476 16192
rect 26240 16108 26292 16114
rect 26240 16050 26292 16056
rect 26252 15706 26280 16050
rect 26424 15904 26476 15910
rect 26424 15846 26476 15852
rect 26240 15700 26292 15706
rect 26240 15642 26292 15648
rect 26436 15502 26464 15846
rect 26528 15570 26556 16458
rect 26516 15564 26568 15570
rect 26516 15506 26568 15512
rect 26424 15496 26476 15502
rect 26424 15438 26476 15444
rect 26712 15366 26740 16526
rect 27080 15978 27108 16526
rect 27068 15972 27120 15978
rect 27068 15914 27120 15920
rect 26792 15904 26844 15910
rect 26792 15846 26844 15852
rect 26804 15434 26832 15846
rect 27080 15638 27108 15914
rect 27068 15632 27120 15638
rect 27120 15580 27200 15586
rect 27068 15574 27200 15580
rect 27080 15558 27200 15574
rect 27264 15570 27292 16526
rect 27068 15496 27120 15502
rect 27068 15438 27120 15444
rect 26792 15428 26844 15434
rect 26792 15370 26844 15376
rect 26700 15360 26752 15366
rect 26700 15302 26752 15308
rect 26332 14952 26384 14958
rect 26332 14894 26384 14900
rect 26344 14346 26372 14894
rect 27080 14618 27108 15438
rect 27172 15162 27200 15558
rect 27252 15564 27304 15570
rect 27252 15506 27304 15512
rect 27356 15434 27384 16526
rect 27344 15428 27396 15434
rect 27344 15370 27396 15376
rect 27160 15156 27212 15162
rect 27160 15098 27212 15104
rect 27252 15020 27304 15026
rect 27448 15008 27476 17002
rect 27540 16114 27568 18142
rect 27724 17678 27752 18226
rect 27712 17672 27764 17678
rect 27712 17614 27764 17620
rect 27620 16788 27672 16794
rect 27620 16730 27672 16736
rect 27528 16108 27580 16114
rect 27528 16050 27580 16056
rect 27632 16046 27660 16730
rect 27620 16040 27672 16046
rect 27620 15982 27672 15988
rect 27252 14962 27304 14968
rect 27356 14980 27476 15008
rect 27068 14612 27120 14618
rect 27068 14554 27120 14560
rect 27264 14414 27292 14962
rect 27252 14408 27304 14414
rect 27252 14350 27304 14356
rect 26332 14340 26384 14346
rect 26332 14282 26384 14288
rect 27252 14272 27304 14278
rect 27252 14214 27304 14220
rect 27264 13938 27292 14214
rect 27252 13932 27304 13938
rect 27252 13874 27304 13880
rect 26516 13864 26568 13870
rect 26516 13806 26568 13812
rect 26148 12232 26200 12238
rect 26148 12174 26200 12180
rect 26160 11150 26188 12174
rect 26148 11144 26200 11150
rect 26148 11086 26200 11092
rect 26160 10130 26188 11086
rect 26528 10674 26556 13806
rect 27158 11792 27214 11801
rect 27158 11727 27160 11736
rect 27212 11727 27214 11736
rect 27252 11756 27304 11762
rect 27160 11698 27212 11704
rect 27356 11744 27384 14980
rect 27816 14550 27844 31214
rect 27908 30326 27936 35158
rect 28172 34604 28224 34610
rect 28172 34546 28224 34552
rect 28080 30796 28132 30802
rect 28080 30738 28132 30744
rect 27896 30320 27948 30326
rect 27896 30262 27948 30268
rect 28092 30258 28120 30738
rect 28080 30252 28132 30258
rect 28080 30194 28132 30200
rect 27988 29504 28040 29510
rect 27988 29446 28040 29452
rect 28000 29306 28028 29446
rect 27988 29300 28040 29306
rect 27988 29242 28040 29248
rect 27896 29164 27948 29170
rect 27896 29106 27948 29112
rect 27908 25906 27936 29106
rect 28000 28558 28028 29242
rect 28092 28762 28120 30194
rect 28184 29102 28212 34546
rect 28172 29096 28224 29102
rect 28172 29038 28224 29044
rect 28080 28756 28132 28762
rect 28080 28698 28132 28704
rect 27988 28552 28040 28558
rect 27988 28494 28040 28500
rect 27896 25900 27948 25906
rect 27896 25842 27948 25848
rect 27988 25832 28040 25838
rect 27988 25774 28040 25780
rect 27896 25152 27948 25158
rect 27896 25094 27948 25100
rect 27908 23594 27936 25094
rect 27896 23588 27948 23594
rect 27896 23530 27948 23536
rect 28000 19854 28028 25774
rect 28172 24064 28224 24070
rect 28172 24006 28224 24012
rect 28184 23730 28212 24006
rect 28172 23724 28224 23730
rect 28172 23666 28224 23672
rect 28184 21554 28212 23666
rect 28276 23526 28304 36110
rect 28368 34746 28396 36230
rect 28460 36038 28488 39782
rect 29196 38758 29224 45426
rect 29748 44402 29776 45426
rect 29736 44396 29788 44402
rect 29736 44338 29788 44344
rect 29748 44010 29776 44338
rect 29748 43982 29868 44010
rect 29736 43920 29788 43926
rect 29736 43862 29788 43868
rect 29748 42770 29776 43862
rect 29840 43858 29868 43982
rect 29828 43852 29880 43858
rect 29828 43794 29880 43800
rect 30104 43784 30156 43790
rect 30104 43726 30156 43732
rect 30472 43784 30524 43790
rect 30472 43726 30524 43732
rect 30656 43784 30708 43790
rect 30656 43726 30708 43732
rect 29828 43716 29880 43722
rect 29828 43658 29880 43664
rect 29840 43296 29868 43658
rect 30116 43314 30144 43726
rect 30484 43382 30512 43726
rect 30668 43450 30696 43726
rect 31116 43648 31168 43654
rect 31116 43590 31168 43596
rect 30656 43444 30708 43450
rect 30656 43386 30708 43392
rect 30472 43376 30524 43382
rect 30472 43318 30524 43324
rect 29920 43308 29972 43314
rect 29840 43268 29920 43296
rect 29920 43250 29972 43256
rect 30104 43308 30156 43314
rect 30104 43250 30156 43256
rect 29932 43178 29960 43250
rect 30288 43240 30340 43246
rect 30288 43182 30340 43188
rect 29920 43172 29972 43178
rect 29920 43114 29972 43120
rect 29932 42906 29960 43114
rect 30012 43104 30064 43110
rect 30012 43046 30064 43052
rect 29920 42900 29972 42906
rect 29920 42842 29972 42848
rect 29736 42764 29788 42770
rect 29736 42706 29788 42712
rect 30024 42702 30052 43046
rect 30300 42922 30328 43182
rect 30116 42894 30328 42922
rect 30012 42696 30064 42702
rect 30012 42638 30064 42644
rect 30116 41818 30144 42894
rect 30288 42764 30340 42770
rect 30288 42706 30340 42712
rect 30196 42628 30248 42634
rect 30196 42570 30248 42576
rect 30104 41812 30156 41818
rect 30104 41754 30156 41760
rect 29460 41676 29512 41682
rect 29460 41618 29512 41624
rect 29472 40934 29500 41618
rect 30104 41268 30156 41274
rect 30104 41210 30156 41216
rect 29460 40928 29512 40934
rect 29460 40870 29512 40876
rect 29472 39506 29500 40870
rect 29460 39500 29512 39506
rect 29460 39442 29512 39448
rect 30116 39302 30144 41210
rect 30208 40934 30236 42570
rect 30300 41818 30328 42706
rect 30484 42362 30512 43318
rect 30668 43314 30696 43386
rect 30564 43308 30616 43314
rect 30564 43250 30616 43256
rect 30656 43308 30708 43314
rect 30656 43250 30708 43256
rect 31024 43308 31076 43314
rect 31024 43250 31076 43256
rect 30576 42634 30604 43250
rect 30564 42628 30616 42634
rect 30564 42570 30616 42576
rect 30840 42560 30892 42566
rect 30840 42502 30892 42508
rect 30472 42356 30524 42362
rect 30472 42298 30524 42304
rect 30852 42294 30880 42502
rect 30840 42288 30892 42294
rect 30840 42230 30892 42236
rect 30380 42084 30432 42090
rect 30380 42026 30432 42032
rect 30288 41812 30340 41818
rect 30288 41754 30340 41760
rect 30196 40928 30248 40934
rect 30196 40870 30248 40876
rect 30208 39982 30236 40870
rect 30288 40724 30340 40730
rect 30392 40712 30420 42026
rect 31036 42022 31064 43250
rect 31128 43178 31156 43590
rect 31484 43376 31536 43382
rect 31484 43318 31536 43324
rect 31116 43172 31168 43178
rect 31116 43114 31168 43120
rect 31128 42226 31156 43114
rect 31300 43104 31352 43110
rect 31300 43046 31352 43052
rect 31208 42628 31260 42634
rect 31208 42570 31260 42576
rect 31116 42220 31168 42226
rect 31116 42162 31168 42168
rect 31220 42158 31248 42570
rect 31312 42226 31340 43046
rect 31496 42702 31524 43318
rect 31944 43308 31996 43314
rect 31944 43250 31996 43256
rect 31956 42702 31984 43250
rect 31484 42696 31536 42702
rect 31484 42638 31536 42644
rect 31944 42696 31996 42702
rect 31944 42638 31996 42644
rect 31392 42628 31444 42634
rect 31392 42570 31444 42576
rect 31300 42220 31352 42226
rect 31300 42162 31352 42168
rect 31208 42152 31260 42158
rect 31208 42094 31260 42100
rect 31024 42016 31076 42022
rect 31024 41958 31076 41964
rect 31036 41614 31064 41958
rect 30748 41608 30800 41614
rect 30748 41550 30800 41556
rect 31024 41608 31076 41614
rect 31024 41550 31076 41556
rect 30340 40684 30420 40712
rect 30288 40666 30340 40672
rect 30472 40656 30524 40662
rect 30472 40598 30524 40604
rect 30484 40118 30512 40598
rect 30472 40112 30524 40118
rect 30472 40054 30524 40060
rect 30196 39976 30248 39982
rect 30196 39918 30248 39924
rect 30380 39840 30432 39846
rect 30380 39782 30432 39788
rect 30104 39296 30156 39302
rect 30104 39238 30156 39244
rect 29736 38956 29788 38962
rect 29736 38898 29788 38904
rect 29184 38752 29236 38758
rect 29184 38694 29236 38700
rect 29748 38554 29776 38898
rect 29736 38548 29788 38554
rect 29736 38490 29788 38496
rect 30116 38282 30144 39238
rect 28540 38276 28592 38282
rect 28540 38218 28592 38224
rect 30104 38276 30156 38282
rect 30104 38218 30156 38224
rect 28552 38010 28580 38218
rect 28540 38004 28592 38010
rect 28540 37946 28592 37952
rect 28632 36780 28684 36786
rect 28632 36722 28684 36728
rect 28644 36378 28672 36722
rect 28724 36576 28776 36582
rect 28724 36518 28776 36524
rect 28632 36372 28684 36378
rect 28632 36314 28684 36320
rect 28448 36032 28500 36038
rect 28448 35974 28500 35980
rect 28736 35086 28764 36518
rect 30116 35834 30144 38218
rect 30392 38214 30420 39782
rect 30484 39642 30512 40054
rect 30760 39982 30788 41550
rect 30932 41472 30984 41478
rect 30932 41414 30984 41420
rect 30944 41138 30972 41414
rect 31220 41274 31248 42094
rect 31404 42090 31432 42570
rect 31392 42084 31444 42090
rect 31392 42026 31444 42032
rect 31496 41818 31524 42638
rect 31956 42294 31984 42638
rect 31944 42288 31996 42294
rect 31944 42230 31996 42236
rect 32128 42220 32180 42226
rect 32128 42162 32180 42168
rect 32036 42016 32088 42022
rect 32036 41958 32088 41964
rect 31484 41812 31536 41818
rect 31484 41754 31536 41760
rect 32048 41750 32076 41958
rect 32140 41750 32168 42162
rect 32036 41744 32088 41750
rect 32036 41686 32088 41692
rect 32128 41744 32180 41750
rect 32128 41686 32180 41692
rect 31208 41268 31260 41274
rect 31208 41210 31260 41216
rect 30932 41132 30984 41138
rect 30932 41074 30984 41080
rect 30944 40526 30972 41074
rect 30932 40520 30984 40526
rect 30932 40462 30984 40468
rect 31116 40384 31168 40390
rect 31116 40326 31168 40332
rect 30932 40044 30984 40050
rect 30932 39986 30984 39992
rect 30748 39976 30800 39982
rect 30748 39918 30800 39924
rect 30472 39636 30524 39642
rect 30472 39578 30524 39584
rect 30484 39494 30788 39522
rect 30484 39438 30512 39494
rect 30472 39432 30524 39438
rect 30472 39374 30524 39380
rect 30656 39432 30708 39438
rect 30656 39374 30708 39380
rect 30564 39364 30616 39370
rect 30564 39306 30616 39312
rect 30472 39296 30524 39302
rect 30472 39238 30524 39244
rect 30484 38894 30512 39238
rect 30576 39098 30604 39306
rect 30564 39092 30616 39098
rect 30564 39034 30616 39040
rect 30472 38888 30524 38894
rect 30472 38830 30524 38836
rect 30576 38486 30604 39034
rect 30564 38480 30616 38486
rect 30564 38422 30616 38428
rect 30576 38350 30604 38422
rect 30564 38344 30616 38350
rect 30564 38286 30616 38292
rect 30472 38276 30524 38282
rect 30472 38218 30524 38224
rect 30380 38208 30432 38214
rect 30380 38150 30432 38156
rect 30288 36168 30340 36174
rect 30288 36110 30340 36116
rect 30104 35828 30156 35834
rect 30104 35770 30156 35776
rect 30300 35766 30328 36110
rect 30484 35766 30512 38218
rect 30564 38208 30616 38214
rect 30564 38150 30616 38156
rect 30576 37874 30604 38150
rect 30668 37942 30696 39374
rect 30760 39250 30788 39494
rect 30944 39438 30972 39986
rect 31024 39976 31076 39982
rect 31024 39918 31076 39924
rect 30932 39432 30984 39438
rect 30932 39374 30984 39380
rect 30760 39222 30972 39250
rect 30944 38962 30972 39222
rect 31036 39098 31064 39918
rect 31128 39914 31156 40326
rect 31116 39908 31168 39914
rect 31116 39850 31168 39856
rect 32036 39432 32088 39438
rect 32036 39374 32088 39380
rect 31668 39364 31720 39370
rect 31668 39306 31720 39312
rect 31484 39296 31536 39302
rect 31484 39238 31536 39244
rect 31576 39296 31628 39302
rect 31576 39238 31628 39244
rect 31024 39092 31076 39098
rect 31024 39034 31076 39040
rect 30932 38956 30984 38962
rect 30932 38898 30984 38904
rect 30944 38282 30972 38898
rect 31496 38418 31524 39238
rect 31588 38962 31616 39238
rect 31576 38956 31628 38962
rect 31576 38898 31628 38904
rect 31484 38412 31536 38418
rect 31484 38354 31536 38360
rect 31680 38350 31708 39306
rect 32048 38554 32076 39374
rect 32036 38548 32088 38554
rect 32036 38490 32088 38496
rect 31208 38344 31260 38350
rect 31208 38286 31260 38292
rect 31668 38344 31720 38350
rect 31668 38286 31720 38292
rect 30932 38276 30984 38282
rect 30932 38218 30984 38224
rect 31220 38010 31248 38286
rect 31668 38208 31720 38214
rect 31668 38150 31720 38156
rect 31208 38004 31260 38010
rect 31208 37946 31260 37952
rect 30656 37936 30708 37942
rect 30656 37878 30708 37884
rect 30564 37868 30616 37874
rect 30564 37810 30616 37816
rect 31680 37262 31708 38150
rect 31668 37256 31720 37262
rect 31668 37198 31720 37204
rect 31680 36922 31708 37198
rect 31668 36916 31720 36922
rect 31668 36858 31720 36864
rect 30932 35828 30984 35834
rect 30932 35770 30984 35776
rect 30288 35760 30340 35766
rect 30288 35702 30340 35708
rect 30472 35760 30524 35766
rect 30472 35702 30524 35708
rect 29000 35692 29052 35698
rect 29000 35634 29052 35640
rect 30104 35692 30156 35698
rect 30104 35634 30156 35640
rect 28724 35080 28776 35086
rect 28724 35022 28776 35028
rect 28356 34740 28408 34746
rect 28356 34682 28408 34688
rect 28368 33998 28396 34682
rect 28356 33992 28408 33998
rect 28356 33934 28408 33940
rect 28540 32904 28592 32910
rect 28540 32846 28592 32852
rect 28552 32026 28580 32846
rect 28540 32020 28592 32026
rect 28540 31962 28592 31968
rect 28736 31822 28764 35022
rect 29012 34746 29040 35634
rect 29092 35080 29144 35086
rect 29092 35022 29144 35028
rect 29000 34740 29052 34746
rect 29000 34682 29052 34688
rect 29104 32858 29132 35022
rect 29184 34944 29236 34950
rect 29184 34886 29236 34892
rect 29196 34610 29224 34886
rect 30116 34678 30144 35634
rect 30196 35488 30248 35494
rect 30196 35430 30248 35436
rect 30208 35086 30236 35430
rect 30196 35080 30248 35086
rect 30196 35022 30248 35028
rect 30104 34672 30156 34678
rect 30104 34614 30156 34620
rect 29184 34604 29236 34610
rect 29184 34546 29236 34552
rect 29368 34536 29420 34542
rect 29368 34478 29420 34484
rect 29380 33114 29408 34478
rect 30116 33930 30144 34614
rect 30208 33998 30236 35022
rect 30300 34610 30328 35702
rect 30484 35562 30512 35702
rect 30472 35556 30524 35562
rect 30472 35498 30524 35504
rect 30748 35080 30800 35086
rect 30748 35022 30800 35028
rect 30564 34944 30616 34950
rect 30564 34886 30616 34892
rect 30576 34678 30604 34886
rect 30564 34672 30616 34678
rect 30564 34614 30616 34620
rect 30288 34604 30340 34610
rect 30288 34546 30340 34552
rect 30196 33992 30248 33998
rect 30196 33934 30248 33940
rect 30104 33924 30156 33930
rect 30104 33866 30156 33872
rect 29368 33108 29420 33114
rect 29368 33050 29420 33056
rect 29104 32830 29224 32858
rect 29092 32768 29144 32774
rect 29092 32710 29144 32716
rect 29104 32434 29132 32710
rect 29000 32428 29052 32434
rect 29000 32370 29052 32376
rect 29092 32428 29144 32434
rect 29092 32370 29144 32376
rect 28724 31816 28776 31822
rect 28724 31758 28776 31764
rect 28540 29640 28592 29646
rect 28540 29582 28592 29588
rect 28552 28558 28580 29582
rect 28540 28552 28592 28558
rect 28540 28494 28592 28500
rect 28552 27554 28580 28494
rect 28552 27526 28672 27554
rect 28540 27464 28592 27470
rect 28540 27406 28592 27412
rect 28552 26518 28580 27406
rect 28644 27130 28672 27526
rect 28736 27418 28764 31758
rect 29012 31346 29040 32370
rect 29092 31816 29144 31822
rect 29196 31804 29224 32830
rect 29144 31776 29224 31804
rect 29092 31758 29144 31764
rect 29000 31340 29052 31346
rect 29000 31282 29052 31288
rect 28816 30592 28868 30598
rect 28816 30534 28868 30540
rect 28828 30258 28856 30534
rect 28816 30252 28868 30258
rect 28816 30194 28868 30200
rect 28736 27390 28856 27418
rect 28724 27328 28776 27334
rect 28724 27270 28776 27276
rect 28632 27124 28684 27130
rect 28632 27066 28684 27072
rect 28540 26512 28592 26518
rect 28540 26454 28592 26460
rect 28644 26382 28672 27066
rect 28736 27062 28764 27270
rect 28724 27056 28776 27062
rect 28724 26998 28776 27004
rect 28632 26376 28684 26382
rect 28632 26318 28684 26324
rect 28724 26376 28776 26382
rect 28828 26364 28856 27390
rect 29104 27010 29132 31758
rect 29276 30048 29328 30054
rect 29276 29990 29328 29996
rect 29288 29306 29316 29990
rect 29276 29300 29328 29306
rect 29276 29242 29328 29248
rect 29184 29164 29236 29170
rect 29184 29106 29236 29112
rect 28920 26982 29132 27010
rect 28920 26790 28948 26982
rect 29196 26790 29224 29106
rect 29380 27606 29408 33050
rect 30300 32502 30328 34546
rect 30760 34202 30788 35022
rect 30944 35018 30972 35770
rect 31680 35698 31708 36858
rect 31668 35692 31720 35698
rect 31668 35634 31720 35640
rect 31668 35556 31720 35562
rect 31668 35498 31720 35504
rect 31024 35080 31076 35086
rect 31024 35022 31076 35028
rect 30932 35012 30984 35018
rect 30932 34954 30984 34960
rect 30840 34604 30892 34610
rect 30840 34546 30892 34552
rect 30748 34196 30800 34202
rect 30748 34138 30800 34144
rect 30656 32972 30708 32978
rect 30656 32914 30708 32920
rect 30288 32496 30340 32502
rect 30288 32438 30340 32444
rect 30380 32224 30432 32230
rect 30380 32166 30432 32172
rect 30392 31822 30420 32166
rect 30472 31952 30524 31958
rect 30472 31894 30524 31900
rect 30380 31816 30432 31822
rect 30380 31758 30432 31764
rect 30196 31340 30248 31346
rect 30196 31282 30248 31288
rect 30104 30660 30156 30666
rect 30104 30602 30156 30608
rect 30116 29850 30144 30602
rect 30208 30394 30236 31282
rect 30380 30592 30432 30598
rect 30380 30534 30432 30540
rect 30196 30388 30248 30394
rect 30196 30330 30248 30336
rect 30392 30258 30420 30534
rect 30380 30252 30432 30258
rect 30380 30194 30432 30200
rect 30484 30190 30512 31894
rect 30564 30728 30616 30734
rect 30564 30670 30616 30676
rect 30472 30184 30524 30190
rect 30472 30126 30524 30132
rect 30104 29844 30156 29850
rect 30104 29786 30156 29792
rect 30472 28076 30524 28082
rect 30576 28064 30604 30670
rect 30668 29102 30696 32914
rect 30748 30728 30800 30734
rect 30748 30670 30800 30676
rect 30656 29096 30708 29102
rect 30656 29038 30708 29044
rect 30656 28960 30708 28966
rect 30656 28902 30708 28908
rect 30668 28558 30696 28902
rect 30656 28552 30708 28558
rect 30656 28494 30708 28500
rect 30760 28150 30788 30670
rect 30852 30258 30880 34546
rect 31036 34202 31064 35022
rect 31392 34400 31444 34406
rect 31392 34342 31444 34348
rect 31024 34196 31076 34202
rect 31024 34138 31076 34144
rect 31404 34066 31432 34342
rect 31392 34060 31444 34066
rect 31392 34002 31444 34008
rect 31300 33992 31352 33998
rect 31300 33934 31352 33940
rect 31312 33114 31340 33934
rect 31404 33538 31432 34002
rect 31576 33924 31628 33930
rect 31576 33866 31628 33872
rect 31404 33522 31524 33538
rect 31392 33516 31524 33522
rect 31444 33510 31524 33516
rect 31392 33458 31444 33464
rect 31392 33380 31444 33386
rect 31392 33322 31444 33328
rect 31300 33108 31352 33114
rect 31300 33050 31352 33056
rect 31404 32910 31432 33322
rect 31496 32978 31524 33510
rect 31484 32972 31536 32978
rect 31484 32914 31536 32920
rect 31392 32904 31444 32910
rect 31392 32846 31444 32852
rect 31116 32428 31168 32434
rect 31116 32370 31168 32376
rect 31128 32026 31156 32370
rect 31116 32020 31168 32026
rect 31116 31962 31168 31968
rect 31404 31482 31432 32846
rect 31588 32842 31616 33866
rect 31576 32836 31628 32842
rect 31576 32778 31628 32784
rect 31588 32434 31616 32778
rect 31680 32502 31708 35498
rect 32232 34610 32260 47126
rect 33232 47048 33284 47054
rect 33232 46990 33284 46996
rect 33244 46646 33272 46990
rect 33232 46640 33284 46646
rect 33232 46582 33284 46588
rect 33520 46510 33548 49200
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 33140 46504 33192 46510
rect 33140 46446 33192 46452
rect 33508 46504 33560 46510
rect 33508 46446 33560 46452
rect 33152 46170 33180 46446
rect 35440 46368 35492 46374
rect 35440 46310 35492 46316
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 33140 46164 33192 46170
rect 33140 46106 33192 46112
rect 35452 46034 35480 46310
rect 36096 46034 36124 49200
rect 36740 46442 36768 49200
rect 37648 46504 37700 46510
rect 37648 46446 37700 46452
rect 36728 46436 36780 46442
rect 36728 46378 36780 46384
rect 35440 46028 35492 46034
rect 35440 45970 35492 45976
rect 36084 46028 36136 46034
rect 36084 45970 36136 45976
rect 32956 45960 33008 45966
rect 32956 45902 33008 45908
rect 32968 45626 32996 45902
rect 35624 45892 35676 45898
rect 35624 45834 35676 45840
rect 34520 45824 34572 45830
rect 34520 45766 34572 45772
rect 32956 45620 33008 45626
rect 32956 45562 33008 45568
rect 32312 43444 32364 43450
rect 32312 43386 32364 43392
rect 32324 42702 32352 43386
rect 32496 43308 32548 43314
rect 32496 43250 32548 43256
rect 32312 42696 32364 42702
rect 32312 42638 32364 42644
rect 32324 41818 32352 42638
rect 32508 42634 32536 43250
rect 32772 43104 32824 43110
rect 32772 43046 32824 43052
rect 32784 42770 32812 43046
rect 32772 42764 32824 42770
rect 32772 42706 32824 42712
rect 32496 42628 32548 42634
rect 32496 42570 32548 42576
rect 32680 42560 32732 42566
rect 32680 42502 32732 42508
rect 32692 42362 32720 42502
rect 32680 42356 32732 42362
rect 32680 42298 32732 42304
rect 32496 42220 32548 42226
rect 32496 42162 32548 42168
rect 32680 42220 32732 42226
rect 32680 42162 32732 42168
rect 32312 41812 32364 41818
rect 32312 41754 32364 41760
rect 32508 41614 32536 42162
rect 32692 42022 32720 42162
rect 32680 42016 32732 42022
rect 32680 41958 32732 41964
rect 32864 42016 32916 42022
rect 32864 41958 32916 41964
rect 32496 41608 32548 41614
rect 32496 41550 32548 41556
rect 32876 40594 32904 41958
rect 32864 40588 32916 40594
rect 32864 40530 32916 40536
rect 32772 40520 32824 40526
rect 32772 40462 32824 40468
rect 32312 40384 32364 40390
rect 32312 40326 32364 40332
rect 32324 40118 32352 40326
rect 32312 40112 32364 40118
rect 32312 40054 32364 40060
rect 32680 40044 32732 40050
rect 32680 39986 32732 39992
rect 32404 39296 32456 39302
rect 32404 39238 32456 39244
rect 32312 38276 32364 38282
rect 32312 38218 32364 38224
rect 32324 36786 32352 38218
rect 32416 38010 32444 39238
rect 32692 39098 32720 39986
rect 32680 39092 32732 39098
rect 32680 39034 32732 39040
rect 32680 38752 32732 38758
rect 32680 38694 32732 38700
rect 32404 38004 32456 38010
rect 32404 37946 32456 37952
rect 32312 36780 32364 36786
rect 32312 36722 32364 36728
rect 32692 36378 32720 38694
rect 32784 38554 32812 40462
rect 32876 40118 32904 40530
rect 32864 40112 32916 40118
rect 32864 40054 32916 40060
rect 32864 39024 32916 39030
rect 32864 38966 32916 38972
rect 32876 38554 32904 38966
rect 32772 38548 32824 38554
rect 32772 38490 32824 38496
rect 32864 38548 32916 38554
rect 32864 38490 32916 38496
rect 32968 38400 32996 45562
rect 34532 45490 34560 45766
rect 35636 45626 35664 45834
rect 35624 45620 35676 45626
rect 35624 45562 35676 45568
rect 37660 45558 37688 46446
rect 38672 46442 38700 49200
rect 39764 47048 39816 47054
rect 39764 46990 39816 46996
rect 40224 47048 40276 47054
rect 40224 46990 40276 46996
rect 39776 46578 39804 46990
rect 39764 46572 39816 46578
rect 39764 46514 39816 46520
rect 39948 46504 40000 46510
rect 39948 46446 40000 46452
rect 38660 46436 38712 46442
rect 38660 46378 38712 46384
rect 39960 46170 39988 46446
rect 39948 46164 40000 46170
rect 39948 46106 40000 46112
rect 40236 46034 40264 46990
rect 40604 46034 40632 49200
rect 41420 47048 41472 47054
rect 41420 46990 41472 46996
rect 41432 46578 41460 46990
rect 41420 46572 41472 46578
rect 41420 46514 41472 46520
rect 41892 46442 41920 49200
rect 42536 47054 42564 49200
rect 42892 47184 42944 47190
rect 42892 47126 42944 47132
rect 42524 47048 42576 47054
rect 42524 46990 42576 46996
rect 42800 46504 42852 46510
rect 42800 46446 42852 46452
rect 41880 46436 41932 46442
rect 41880 46378 41932 46384
rect 41328 46096 41380 46102
rect 41328 46038 41380 46044
rect 40224 46028 40276 46034
rect 40224 45970 40276 45976
rect 40592 46028 40644 46034
rect 40592 45970 40644 45976
rect 38660 45960 38712 45966
rect 38660 45902 38712 45908
rect 39948 45960 40000 45966
rect 39948 45902 40000 45908
rect 37648 45552 37700 45558
rect 37648 45494 37700 45500
rect 38672 45490 38700 45902
rect 39960 45490 39988 45902
rect 40224 45892 40276 45898
rect 40224 45834 40276 45840
rect 40236 45626 40264 45834
rect 40224 45620 40276 45626
rect 40224 45562 40276 45568
rect 41340 45490 41368 46038
rect 42812 45558 42840 46446
rect 42800 45552 42852 45558
rect 42800 45494 42852 45500
rect 34520 45484 34572 45490
rect 34520 45426 34572 45432
rect 35624 45484 35676 45490
rect 35624 45426 35676 45432
rect 38660 45484 38712 45490
rect 38660 45426 38712 45432
rect 39948 45484 40000 45490
rect 39948 45426 40000 45432
rect 40592 45484 40644 45490
rect 40592 45426 40644 45432
rect 41328 45484 41380 45490
rect 41328 45426 41380 45432
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 33692 43308 33744 43314
rect 33692 43250 33744 43256
rect 34520 43308 34572 43314
rect 34520 43250 34572 43256
rect 33324 43240 33376 43246
rect 33324 43182 33376 43188
rect 33336 42838 33364 43182
rect 33508 43172 33560 43178
rect 33508 43114 33560 43120
rect 33324 42832 33376 42838
rect 33324 42774 33376 42780
rect 33336 42226 33364 42774
rect 33416 42696 33468 42702
rect 33416 42638 33468 42644
rect 33428 42226 33456 42638
rect 33324 42220 33376 42226
rect 33324 42162 33376 42168
rect 33416 42220 33468 42226
rect 33416 42162 33468 42168
rect 33428 41682 33456 42162
rect 33416 41676 33468 41682
rect 33416 41618 33468 41624
rect 33048 41064 33100 41070
rect 33048 41006 33100 41012
rect 33060 40526 33088 41006
rect 33048 40520 33100 40526
rect 33048 40462 33100 40468
rect 33060 39982 33088 40462
rect 33048 39976 33100 39982
rect 33048 39918 33100 39924
rect 33140 39092 33192 39098
rect 33140 39034 33192 39040
rect 32876 38372 32996 38400
rect 32680 36372 32732 36378
rect 32680 36314 32732 36320
rect 32692 36242 32720 36314
rect 32680 36236 32732 36242
rect 32680 36178 32732 36184
rect 32692 35630 32720 36178
rect 32680 35624 32732 35630
rect 32680 35566 32732 35572
rect 32220 34604 32272 34610
rect 32220 34546 32272 34552
rect 31760 33992 31812 33998
rect 31760 33934 31812 33940
rect 31772 33318 31800 33934
rect 31760 33312 31812 33318
rect 31760 33254 31812 33260
rect 32220 33312 32272 33318
rect 32220 33254 32272 33260
rect 31852 33040 31904 33046
rect 31852 32982 31904 32988
rect 31668 32496 31720 32502
rect 31668 32438 31720 32444
rect 31576 32428 31628 32434
rect 31576 32370 31628 32376
rect 31392 31476 31444 31482
rect 31392 31418 31444 31424
rect 31404 30734 31432 31418
rect 31392 30728 31444 30734
rect 31392 30670 31444 30676
rect 30840 30252 30892 30258
rect 30840 30194 30892 30200
rect 31024 30048 31076 30054
rect 31024 29990 31076 29996
rect 30840 29164 30892 29170
rect 30840 29106 30892 29112
rect 30852 28218 30880 29106
rect 31036 29034 31064 29990
rect 31680 29782 31708 32438
rect 31864 31822 31892 32982
rect 32232 32910 32260 33254
rect 32220 32904 32272 32910
rect 32220 32846 32272 32852
rect 32128 32768 32180 32774
rect 32128 32710 32180 32716
rect 32140 31890 32168 32710
rect 32232 32026 32260 32846
rect 32680 32564 32732 32570
rect 32680 32506 32732 32512
rect 32692 32230 32720 32506
rect 32680 32224 32732 32230
rect 32680 32166 32732 32172
rect 32220 32020 32272 32026
rect 32220 31962 32272 31968
rect 32128 31884 32180 31890
rect 32128 31826 32180 31832
rect 31852 31816 31904 31822
rect 31852 31758 31904 31764
rect 32588 31748 32640 31754
rect 32588 31690 32640 31696
rect 32128 31340 32180 31346
rect 32128 31282 32180 31288
rect 32140 30734 32168 31282
rect 32600 30938 32628 31690
rect 32692 31278 32720 32166
rect 32772 31816 32824 31822
rect 32772 31758 32824 31764
rect 32784 31278 32812 31758
rect 32680 31272 32732 31278
rect 32680 31214 32732 31220
rect 32772 31272 32824 31278
rect 32772 31214 32824 31220
rect 32588 30932 32640 30938
rect 32588 30874 32640 30880
rect 32692 30734 32720 31214
rect 32128 30728 32180 30734
rect 32128 30670 32180 30676
rect 32680 30728 32732 30734
rect 32680 30670 32732 30676
rect 31852 30184 31904 30190
rect 31852 30126 31904 30132
rect 31668 29776 31720 29782
rect 31668 29718 31720 29724
rect 31864 29034 31892 30126
rect 31024 29028 31076 29034
rect 31024 28970 31076 28976
rect 31852 29028 31904 29034
rect 31852 28970 31904 28976
rect 30840 28212 30892 28218
rect 30840 28154 30892 28160
rect 30748 28144 30800 28150
rect 30748 28086 30800 28092
rect 30524 28036 30604 28064
rect 30472 28018 30524 28024
rect 29368 27600 29420 27606
rect 29368 27542 29420 27548
rect 29276 27464 29328 27470
rect 29276 27406 29328 27412
rect 28908 26784 28960 26790
rect 28908 26726 28960 26732
rect 29184 26784 29236 26790
rect 29184 26726 29236 26732
rect 28920 26382 28948 26726
rect 29196 26382 29224 26726
rect 28776 26336 28856 26364
rect 28908 26376 28960 26382
rect 28724 26318 28776 26324
rect 28908 26318 28960 26324
rect 29184 26376 29236 26382
rect 29184 26318 29236 26324
rect 28356 25900 28408 25906
rect 28356 25842 28408 25848
rect 28368 25294 28396 25842
rect 28356 25288 28408 25294
rect 28356 25230 28408 25236
rect 28736 25158 28764 26318
rect 29288 25838 29316 27406
rect 29276 25832 29328 25838
rect 29276 25774 29328 25780
rect 29380 25362 29408 27542
rect 29460 27056 29512 27062
rect 29460 26998 29512 27004
rect 29368 25356 29420 25362
rect 29368 25298 29420 25304
rect 28724 25152 28776 25158
rect 28724 25094 28776 25100
rect 29472 24750 29500 26998
rect 30380 26580 30432 26586
rect 30380 26522 30432 26528
rect 29736 26308 29788 26314
rect 29736 26250 29788 26256
rect 29644 24948 29696 24954
rect 29644 24890 29696 24896
rect 29460 24744 29512 24750
rect 29380 24704 29460 24732
rect 28264 23520 28316 23526
rect 28264 23462 28316 23468
rect 29380 22710 29408 24704
rect 29460 24686 29512 24692
rect 29656 24614 29684 24890
rect 29748 24614 29776 26250
rect 30196 25764 30248 25770
rect 30196 25706 30248 25712
rect 30208 25294 30236 25706
rect 30104 25288 30156 25294
rect 30104 25230 30156 25236
rect 30196 25288 30248 25294
rect 30196 25230 30248 25236
rect 29920 25152 29972 25158
rect 29920 25094 29972 25100
rect 29932 24886 29960 25094
rect 29920 24880 29972 24886
rect 29920 24822 29972 24828
rect 29644 24608 29696 24614
rect 29644 24550 29696 24556
rect 29736 24608 29788 24614
rect 29736 24550 29788 24556
rect 29656 23730 29684 24550
rect 30116 24410 30144 25230
rect 30104 24404 30156 24410
rect 30104 24346 30156 24352
rect 29828 24064 29880 24070
rect 29828 24006 29880 24012
rect 29552 23724 29604 23730
rect 29552 23666 29604 23672
rect 29644 23724 29696 23730
rect 29644 23666 29696 23672
rect 29460 23520 29512 23526
rect 29460 23462 29512 23468
rect 29368 22704 29420 22710
rect 29368 22646 29420 22652
rect 29472 22642 29500 23462
rect 29564 23322 29592 23666
rect 29840 23662 29868 24006
rect 29920 23792 29972 23798
rect 29920 23734 29972 23740
rect 29828 23656 29880 23662
rect 29828 23598 29880 23604
rect 29552 23316 29604 23322
rect 29552 23258 29604 23264
rect 29000 22636 29052 22642
rect 29000 22578 29052 22584
rect 29460 22636 29512 22642
rect 29460 22578 29512 22584
rect 29012 21554 29040 22578
rect 29840 22234 29868 23598
rect 29932 23118 29960 23734
rect 30104 23588 30156 23594
rect 30104 23530 30156 23536
rect 30116 23118 30144 23530
rect 29920 23112 29972 23118
rect 29920 23054 29972 23060
rect 30104 23112 30156 23118
rect 30104 23054 30156 23060
rect 29828 22228 29880 22234
rect 29828 22170 29880 22176
rect 28172 21548 28224 21554
rect 28172 21490 28224 21496
rect 28724 21548 28776 21554
rect 28724 21490 28776 21496
rect 29000 21548 29052 21554
rect 29000 21490 29052 21496
rect 29276 21548 29328 21554
rect 29276 21490 29328 21496
rect 28540 21344 28592 21350
rect 28540 21286 28592 21292
rect 28356 21072 28408 21078
rect 28356 21014 28408 21020
rect 28368 20942 28396 21014
rect 28172 20936 28224 20942
rect 28172 20878 28224 20884
rect 28356 20936 28408 20942
rect 28356 20878 28408 20884
rect 28184 20058 28212 20878
rect 28448 20800 28500 20806
rect 28448 20742 28500 20748
rect 28460 20466 28488 20742
rect 28552 20534 28580 21286
rect 28736 20942 28764 21490
rect 29000 21412 29052 21418
rect 29000 21354 29052 21360
rect 28908 21344 28960 21350
rect 29012 21321 29040 21354
rect 28908 21286 28960 21292
rect 28998 21312 29054 21321
rect 28632 20936 28684 20942
rect 28632 20878 28684 20884
rect 28724 20936 28776 20942
rect 28724 20878 28776 20884
rect 28644 20806 28672 20878
rect 28632 20800 28684 20806
rect 28632 20742 28684 20748
rect 28540 20528 28592 20534
rect 28540 20470 28592 20476
rect 28448 20460 28500 20466
rect 28448 20402 28500 20408
rect 28644 20346 28672 20742
rect 28920 20466 28948 21286
rect 28998 21247 29054 21256
rect 29288 21146 29316 21490
rect 29276 21140 29328 21146
rect 29276 21082 29328 21088
rect 29184 20596 29236 20602
rect 29184 20538 29236 20544
rect 28908 20460 28960 20466
rect 28908 20402 28960 20408
rect 28552 20318 28672 20346
rect 28172 20052 28224 20058
rect 28172 19994 28224 20000
rect 27988 19848 28040 19854
rect 27988 19790 28040 19796
rect 28448 19848 28500 19854
rect 28448 19790 28500 19796
rect 28264 19372 28316 19378
rect 28264 19314 28316 19320
rect 28080 19304 28132 19310
rect 28080 19246 28132 19252
rect 27988 18148 28040 18154
rect 27988 18090 28040 18096
rect 28000 17746 28028 18090
rect 28092 17882 28120 19246
rect 28172 18284 28224 18290
rect 28172 18226 28224 18232
rect 28080 17876 28132 17882
rect 28080 17818 28132 17824
rect 27988 17740 28040 17746
rect 27988 17682 28040 17688
rect 28184 16454 28212 18226
rect 28276 17814 28304 19314
rect 28264 17808 28316 17814
rect 28264 17750 28316 17756
rect 28276 17542 28304 17750
rect 28460 17610 28488 19790
rect 28552 18834 28580 20318
rect 29000 20256 29052 20262
rect 29000 20198 29052 20204
rect 29012 20058 29040 20198
rect 29000 20052 29052 20058
rect 29000 19994 29052 20000
rect 28724 19848 28776 19854
rect 28724 19790 28776 19796
rect 28736 19514 28764 19790
rect 28724 19508 28776 19514
rect 28724 19450 28776 19456
rect 28724 19372 28776 19378
rect 28724 19314 28776 19320
rect 28632 19304 28684 19310
rect 28632 19246 28684 19252
rect 28540 18828 28592 18834
rect 28540 18770 28592 18776
rect 28540 18692 28592 18698
rect 28540 18634 28592 18640
rect 28552 18086 28580 18634
rect 28644 18290 28672 19246
rect 28736 19242 28764 19314
rect 28724 19236 28776 19242
rect 28724 19178 28776 19184
rect 29000 19168 29052 19174
rect 29000 19110 29052 19116
rect 29012 18970 29040 19110
rect 29000 18964 29052 18970
rect 29000 18906 29052 18912
rect 28632 18284 28684 18290
rect 28632 18226 28684 18232
rect 29012 18086 29040 18906
rect 29196 18630 29224 20538
rect 29368 20256 29420 20262
rect 29368 20198 29420 20204
rect 29380 19378 29408 20198
rect 29460 19712 29512 19718
rect 29460 19654 29512 19660
rect 29472 19514 29500 19654
rect 29460 19508 29512 19514
rect 29460 19450 29512 19456
rect 29932 19378 29960 23054
rect 30208 22094 30236 25230
rect 30288 24200 30340 24206
rect 30288 24142 30340 24148
rect 30116 22066 30236 22094
rect 30116 20058 30144 22066
rect 30300 21962 30328 24142
rect 30288 21956 30340 21962
rect 30288 21898 30340 21904
rect 30300 20754 30328 21898
rect 30392 21010 30420 26522
rect 30484 25702 30512 28018
rect 30760 26382 30788 28086
rect 30748 26376 30800 26382
rect 30748 26318 30800 26324
rect 30472 25696 30524 25702
rect 30472 25638 30524 25644
rect 30484 22098 30512 25638
rect 31036 25430 31064 28970
rect 31208 27464 31260 27470
rect 31208 27406 31260 27412
rect 31220 26994 31248 27406
rect 31300 27396 31352 27402
rect 31300 27338 31352 27344
rect 31208 26988 31260 26994
rect 31208 26930 31260 26936
rect 31312 26042 31340 27338
rect 31576 26988 31628 26994
rect 31576 26930 31628 26936
rect 31760 26988 31812 26994
rect 31760 26930 31812 26936
rect 31484 26784 31536 26790
rect 31484 26726 31536 26732
rect 31300 26036 31352 26042
rect 31300 25978 31352 25984
rect 31496 25906 31524 26726
rect 31484 25900 31536 25906
rect 31484 25842 31536 25848
rect 31024 25424 31076 25430
rect 31024 25366 31076 25372
rect 30840 25288 30892 25294
rect 30840 25230 30892 25236
rect 30656 24812 30708 24818
rect 30656 24754 30708 24760
rect 30564 23112 30616 23118
rect 30564 23054 30616 23060
rect 30576 22438 30604 23054
rect 30564 22432 30616 22438
rect 30564 22374 30616 22380
rect 30472 22092 30524 22098
rect 30668 22094 30696 24754
rect 30852 24614 30880 25230
rect 31392 25220 31444 25226
rect 31392 25162 31444 25168
rect 31404 24954 31432 25162
rect 31392 24948 31444 24954
rect 31392 24890 31444 24896
rect 30840 24608 30892 24614
rect 30840 24550 30892 24556
rect 30748 24132 30800 24138
rect 30748 24074 30800 24080
rect 30760 23866 30788 24074
rect 30748 23860 30800 23866
rect 30748 23802 30800 23808
rect 30472 22034 30524 22040
rect 30576 22066 30696 22094
rect 30380 21004 30432 21010
rect 30380 20946 30432 20952
rect 30208 20726 30328 20754
rect 30104 20052 30156 20058
rect 30104 19994 30156 20000
rect 29368 19372 29420 19378
rect 29368 19314 29420 19320
rect 29920 19372 29972 19378
rect 29920 19314 29972 19320
rect 29184 18624 29236 18630
rect 29184 18566 29236 18572
rect 30104 18624 30156 18630
rect 30104 18566 30156 18572
rect 28540 18080 28592 18086
rect 28540 18022 28592 18028
rect 29000 18080 29052 18086
rect 29000 18022 29052 18028
rect 29012 17678 29040 18022
rect 29196 17746 29224 18566
rect 30116 18358 30144 18566
rect 30104 18352 30156 18358
rect 30104 18294 30156 18300
rect 29184 17740 29236 17746
rect 29184 17682 29236 17688
rect 29000 17672 29052 17678
rect 29000 17614 29052 17620
rect 28448 17604 28500 17610
rect 28448 17546 28500 17552
rect 28632 17604 28684 17610
rect 28632 17546 28684 17552
rect 28264 17536 28316 17542
rect 28264 17478 28316 17484
rect 28264 16516 28316 16522
rect 28264 16458 28316 16464
rect 28172 16448 28224 16454
rect 28172 16390 28224 16396
rect 28184 16182 28212 16390
rect 28172 16176 28224 16182
rect 28172 16118 28224 16124
rect 27988 16040 28040 16046
rect 27988 15982 28040 15988
rect 27804 14544 27856 14550
rect 27804 14486 27856 14492
rect 27712 14408 27764 14414
rect 27712 14350 27764 14356
rect 27620 14272 27672 14278
rect 27620 14214 27672 14220
rect 27632 13530 27660 14214
rect 27620 13524 27672 13530
rect 27620 13466 27672 13472
rect 27724 13326 27752 14350
rect 27712 13320 27764 13326
rect 27712 13262 27764 13268
rect 27816 12434 27844 14486
rect 27724 12406 27844 12434
rect 27528 12096 27580 12102
rect 27528 12038 27580 12044
rect 27540 11830 27568 12038
rect 27528 11824 27580 11830
rect 27528 11766 27580 11772
rect 27304 11716 27384 11744
rect 27252 11698 27304 11704
rect 26516 10668 26568 10674
rect 27356 10656 27384 11716
rect 27540 11150 27568 11766
rect 27724 11558 27752 12406
rect 27804 12164 27856 12170
rect 27804 12106 27856 12112
rect 27816 11762 27844 12106
rect 28000 11898 28028 15982
rect 28276 15638 28304 16458
rect 28264 15632 28316 15638
rect 28264 15574 28316 15580
rect 28644 15502 28672 17546
rect 30208 17270 30236 20726
rect 30288 19440 30340 19446
rect 30288 19382 30340 19388
rect 30300 18290 30328 19382
rect 30576 18766 30604 22066
rect 30656 22024 30708 22030
rect 30656 21966 30708 21972
rect 30668 21622 30696 21966
rect 30656 21616 30708 21622
rect 30656 21558 30708 21564
rect 30668 19922 30696 21558
rect 30656 19916 30708 19922
rect 30656 19858 30708 19864
rect 30380 18760 30432 18766
rect 30564 18760 30616 18766
rect 30380 18702 30432 18708
rect 30484 18708 30564 18714
rect 30484 18702 30616 18708
rect 30288 18284 30340 18290
rect 30288 18226 30340 18232
rect 30196 17264 30248 17270
rect 30196 17206 30248 17212
rect 30300 16794 30328 18226
rect 30392 17882 30420 18702
rect 30484 18686 30604 18702
rect 30380 17876 30432 17882
rect 30380 17818 30432 17824
rect 30288 16788 30340 16794
rect 30288 16730 30340 16736
rect 30300 16658 30328 16730
rect 30288 16652 30340 16658
rect 30288 16594 30340 16600
rect 28632 15496 28684 15502
rect 28632 15438 28684 15444
rect 28540 15360 28592 15366
rect 28540 15302 28592 15308
rect 28552 14414 28580 15302
rect 28540 14408 28592 14414
rect 28540 14350 28592 14356
rect 28264 14068 28316 14074
rect 28264 14010 28316 14016
rect 28276 13326 28304 14010
rect 28264 13320 28316 13326
rect 28264 13262 28316 13268
rect 28356 13252 28408 13258
rect 28356 13194 28408 13200
rect 27988 11892 28040 11898
rect 27988 11834 28040 11840
rect 27804 11756 27856 11762
rect 27804 11698 27856 11704
rect 27712 11552 27764 11558
rect 27712 11494 27764 11500
rect 27528 11144 27580 11150
rect 27528 11086 27580 11092
rect 27528 10668 27580 10674
rect 27356 10628 27528 10656
rect 26516 10610 26568 10616
rect 27528 10610 27580 10616
rect 27712 10668 27764 10674
rect 27712 10610 27764 10616
rect 27724 10266 27752 10610
rect 27896 10464 27948 10470
rect 27896 10406 27948 10412
rect 27712 10260 27764 10266
rect 27712 10202 27764 10208
rect 26148 10124 26200 10130
rect 26148 10066 26200 10072
rect 27724 9586 27752 10202
rect 27908 10062 27936 10406
rect 27896 10056 27948 10062
rect 27896 9998 27948 10004
rect 28172 10056 28224 10062
rect 28172 9998 28224 10004
rect 28184 9722 28212 9998
rect 28172 9716 28224 9722
rect 28172 9658 28224 9664
rect 27712 9580 27764 9586
rect 27712 9522 27764 9528
rect 27160 3936 27212 3942
rect 27160 3878 27212 3884
rect 26424 3596 26476 3602
rect 26424 3538 26476 3544
rect 26056 2508 26108 2514
rect 26056 2450 26108 2456
rect 26436 800 26464 3538
rect 27172 3058 27200 3878
rect 27344 3392 27396 3398
rect 27344 3334 27396 3340
rect 27356 3126 27384 3334
rect 27344 3120 27396 3126
rect 27344 3062 27396 3068
rect 27160 3052 27212 3058
rect 27160 2994 27212 3000
rect 27712 2984 27764 2990
rect 27712 2926 27764 2932
rect 27724 800 27752 2926
rect 28368 2854 28396 13194
rect 28644 12434 28672 15438
rect 29276 15428 29328 15434
rect 29276 15370 29328 15376
rect 29092 15088 29144 15094
rect 29092 15030 29144 15036
rect 29000 15020 29052 15026
rect 29000 14962 29052 14968
rect 28724 14816 28776 14822
rect 28724 14758 28776 14764
rect 28736 14414 28764 14758
rect 29012 14618 29040 14962
rect 29000 14612 29052 14618
rect 29000 14554 29052 14560
rect 28724 14408 28776 14414
rect 28724 14350 28776 14356
rect 28908 14340 28960 14346
rect 28908 14282 28960 14288
rect 28920 14074 28948 14282
rect 28908 14068 28960 14074
rect 28908 14010 28960 14016
rect 29104 14006 29132 15030
rect 29288 14618 29316 15370
rect 30300 15094 30328 16594
rect 30484 15978 30512 18686
rect 30760 17202 30788 23802
rect 30852 22710 30880 24550
rect 31588 24274 31616 26930
rect 31772 24750 31800 26930
rect 31668 24744 31720 24750
rect 31668 24686 31720 24692
rect 31760 24744 31812 24750
rect 31760 24686 31812 24692
rect 31576 24268 31628 24274
rect 31576 24210 31628 24216
rect 31680 23594 31708 24686
rect 31668 23588 31720 23594
rect 31668 23530 31720 23536
rect 31484 23520 31536 23526
rect 31484 23462 31536 23468
rect 31496 23050 31524 23462
rect 31484 23044 31536 23050
rect 31484 22986 31536 22992
rect 30840 22704 30892 22710
rect 30840 22646 30892 22652
rect 31392 22432 31444 22438
rect 31392 22374 31444 22380
rect 31208 22024 31260 22030
rect 31208 21966 31260 21972
rect 31116 21888 31168 21894
rect 31116 21830 31168 21836
rect 31128 21554 31156 21830
rect 31220 21690 31248 21966
rect 31208 21684 31260 21690
rect 31208 21626 31260 21632
rect 31404 21554 31432 22374
rect 31024 21548 31076 21554
rect 31024 21490 31076 21496
rect 31116 21548 31168 21554
rect 31116 21490 31168 21496
rect 31392 21548 31444 21554
rect 31392 21490 31444 21496
rect 31036 21078 31064 21490
rect 31208 21480 31260 21486
rect 31208 21422 31260 21428
rect 31024 21072 31076 21078
rect 31024 21014 31076 21020
rect 31220 20806 31248 21422
rect 31392 21004 31444 21010
rect 31392 20946 31444 20952
rect 31208 20800 31260 20806
rect 31208 20742 31260 20748
rect 31024 20460 31076 20466
rect 31024 20402 31076 20408
rect 31208 20460 31260 20466
rect 31208 20402 31260 20408
rect 30932 20256 30984 20262
rect 30932 20198 30984 20204
rect 30944 19854 30972 20198
rect 30932 19848 30984 19854
rect 30932 19790 30984 19796
rect 31036 19514 31064 20402
rect 31024 19508 31076 19514
rect 31024 19450 31076 19456
rect 31024 19372 31076 19378
rect 31024 19314 31076 19320
rect 30840 18828 30892 18834
rect 30840 18770 30892 18776
rect 30748 17196 30800 17202
rect 30748 17138 30800 17144
rect 30564 16516 30616 16522
rect 30564 16458 30616 16464
rect 30472 15972 30524 15978
rect 30472 15914 30524 15920
rect 30576 15706 30604 16458
rect 30656 15904 30708 15910
rect 30656 15846 30708 15852
rect 30564 15700 30616 15706
rect 30564 15642 30616 15648
rect 30668 15502 30696 15846
rect 30656 15496 30708 15502
rect 30656 15438 30708 15444
rect 30288 15088 30340 15094
rect 30288 15030 30340 15036
rect 30380 15088 30432 15094
rect 30380 15030 30432 15036
rect 30300 14890 30328 15030
rect 30288 14884 30340 14890
rect 30288 14826 30340 14832
rect 29276 14612 29328 14618
rect 29276 14554 29328 14560
rect 29288 14414 29316 14554
rect 30392 14550 30420 15030
rect 30104 14544 30156 14550
rect 30024 14504 30104 14532
rect 29828 14476 29880 14482
rect 30024 14464 30052 14504
rect 30104 14486 30156 14492
rect 30380 14544 30432 14550
rect 30380 14486 30432 14492
rect 29880 14436 30052 14464
rect 29828 14418 29880 14424
rect 29276 14408 29328 14414
rect 29276 14350 29328 14356
rect 29932 14346 30328 14362
rect 29828 14340 29880 14346
rect 29932 14340 30340 14346
rect 29932 14334 30288 14340
rect 29932 14328 29960 14334
rect 29880 14300 29960 14328
rect 29828 14282 29880 14288
rect 30288 14282 30340 14288
rect 30012 14272 30064 14278
rect 30012 14214 30064 14220
rect 30380 14272 30432 14278
rect 30380 14214 30432 14220
rect 30024 14006 30052 14214
rect 29092 14000 29144 14006
rect 29092 13942 29144 13948
rect 30012 14000 30064 14006
rect 30012 13942 30064 13948
rect 30392 13530 30420 14214
rect 30380 13524 30432 13530
rect 30380 13466 30432 13472
rect 30760 13326 30788 17138
rect 30852 15706 30880 18770
rect 31036 17678 31064 19314
rect 31220 18834 31248 20402
rect 31300 20392 31352 20398
rect 31404 20380 31432 20946
rect 31352 20352 31432 20380
rect 31300 20334 31352 20340
rect 31312 18902 31340 20334
rect 31496 19378 31524 22986
rect 31576 21956 31628 21962
rect 31576 21898 31628 21904
rect 31588 21690 31616 21898
rect 31576 21684 31628 21690
rect 31576 21626 31628 21632
rect 31680 20466 31708 23530
rect 31772 22778 31800 24686
rect 31864 23662 31892 28970
rect 32140 28762 32168 30670
rect 32876 30258 32904 38372
rect 32956 38276 33008 38282
rect 32956 38218 33008 38224
rect 32968 37874 32996 38218
rect 33048 38208 33100 38214
rect 33048 38150 33100 38156
rect 33060 38010 33088 38150
rect 33048 38004 33100 38010
rect 33048 37946 33100 37952
rect 32956 37868 33008 37874
rect 32956 37810 33008 37816
rect 32956 37664 33008 37670
rect 32956 37606 33008 37612
rect 32968 36786 32996 37606
rect 33152 37126 33180 39034
rect 33416 38412 33468 38418
rect 33416 38354 33468 38360
rect 33428 37942 33456 38354
rect 33520 38350 33548 43114
rect 33704 42158 33732 43250
rect 34532 42906 34560 43250
rect 34796 43240 34848 43246
rect 34796 43182 34848 43188
rect 34704 43104 34756 43110
rect 34624 43064 34704 43092
rect 34520 42900 34572 42906
rect 34520 42842 34572 42848
rect 34244 42764 34296 42770
rect 34244 42706 34296 42712
rect 33692 42152 33744 42158
rect 33744 42100 33824 42106
rect 33692 42094 33824 42100
rect 33704 42078 33824 42094
rect 33796 41614 33824 42078
rect 34152 42016 34204 42022
rect 34152 41958 34204 41964
rect 34060 41812 34112 41818
rect 34060 41754 34112 41760
rect 33784 41608 33836 41614
rect 33784 41550 33836 41556
rect 34072 41546 34100 41754
rect 34060 41540 34112 41546
rect 34060 41482 34112 41488
rect 33876 41132 33928 41138
rect 33876 41074 33928 41080
rect 33888 40730 33916 41074
rect 34072 41070 34100 41482
rect 34060 41064 34112 41070
rect 34060 41006 34112 41012
rect 34164 41002 34192 41958
rect 34152 40996 34204 41002
rect 34152 40938 34204 40944
rect 33876 40724 33928 40730
rect 33876 40666 33928 40672
rect 34164 40662 34192 40938
rect 34152 40656 34204 40662
rect 34152 40598 34204 40604
rect 34256 40458 34284 42706
rect 34428 42628 34480 42634
rect 34428 42570 34480 42576
rect 34440 42362 34468 42570
rect 34428 42356 34480 42362
rect 34428 42298 34480 42304
rect 34532 42294 34560 42842
rect 34520 42288 34572 42294
rect 34520 42230 34572 42236
rect 34624 42226 34652 43064
rect 34704 43046 34756 43052
rect 34808 42786 34836 43182
rect 35440 43172 35492 43178
rect 35440 43114 35492 43120
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 35348 42900 35400 42906
rect 35348 42842 35400 42848
rect 34716 42758 34836 42786
rect 34612 42220 34664 42226
rect 34612 42162 34664 42168
rect 34428 42152 34480 42158
rect 34428 42094 34480 42100
rect 34440 41750 34468 42094
rect 34520 42084 34572 42090
rect 34520 42026 34572 42032
rect 34612 42084 34664 42090
rect 34612 42026 34664 42032
rect 34428 41744 34480 41750
rect 34428 41686 34480 41692
rect 34336 40928 34388 40934
rect 34336 40870 34388 40876
rect 34244 40452 34296 40458
rect 34244 40394 34296 40400
rect 34060 39568 34112 39574
rect 34060 39510 34112 39516
rect 34072 38962 34100 39510
rect 34152 39500 34204 39506
rect 34152 39442 34204 39448
rect 34060 38956 34112 38962
rect 34060 38898 34112 38904
rect 34164 38758 34192 39442
rect 34152 38752 34204 38758
rect 34152 38694 34204 38700
rect 34164 38486 34192 38694
rect 34152 38480 34204 38486
rect 34152 38422 34204 38428
rect 34256 38418 34284 40394
rect 34244 38412 34296 38418
rect 34244 38354 34296 38360
rect 33508 38344 33560 38350
rect 33508 38286 33560 38292
rect 33416 37936 33468 37942
rect 33416 37878 33468 37884
rect 33428 37466 33456 37878
rect 33416 37460 33468 37466
rect 33416 37402 33468 37408
rect 33140 37120 33192 37126
rect 33140 37062 33192 37068
rect 33416 37120 33468 37126
rect 33416 37062 33468 37068
rect 33428 36786 33456 37062
rect 32956 36780 33008 36786
rect 32956 36722 33008 36728
rect 33416 36780 33468 36786
rect 33416 36722 33468 36728
rect 32968 35766 32996 36722
rect 33324 36712 33376 36718
rect 33324 36654 33376 36660
rect 33048 36576 33100 36582
rect 33048 36518 33100 36524
rect 33060 36174 33088 36518
rect 33336 36378 33364 36654
rect 33324 36372 33376 36378
rect 33324 36314 33376 36320
rect 33140 36304 33192 36310
rect 33140 36246 33192 36252
rect 33048 36168 33100 36174
rect 33048 36110 33100 36116
rect 33152 36106 33180 36246
rect 33140 36100 33192 36106
rect 33140 36042 33192 36048
rect 33232 36100 33284 36106
rect 33232 36042 33284 36048
rect 33152 35834 33180 36042
rect 33140 35828 33192 35834
rect 33140 35770 33192 35776
rect 32956 35760 33008 35766
rect 32956 35702 33008 35708
rect 33244 35562 33272 36042
rect 33336 35698 33364 36314
rect 33416 36032 33468 36038
rect 33416 35974 33468 35980
rect 33428 35834 33456 35974
rect 33416 35828 33468 35834
rect 33416 35770 33468 35776
rect 33324 35692 33376 35698
rect 33324 35634 33376 35640
rect 33232 35556 33284 35562
rect 33232 35498 33284 35504
rect 33520 32842 33548 38286
rect 33876 38208 33928 38214
rect 33876 38150 33928 38156
rect 34244 38208 34296 38214
rect 34348 38162 34376 40870
rect 34440 40594 34468 41686
rect 34532 41070 34560 42026
rect 34624 41138 34652 42026
rect 34716 41614 34744 42758
rect 34796 42696 34848 42702
rect 34796 42638 34848 42644
rect 34704 41608 34756 41614
rect 34704 41550 34756 41556
rect 34612 41132 34664 41138
rect 34612 41074 34664 41080
rect 34808 41070 34836 42638
rect 35072 42560 35124 42566
rect 35072 42502 35124 42508
rect 35084 42226 35112 42502
rect 35360 42226 35388 42842
rect 35072 42220 35124 42226
rect 35072 42162 35124 42168
rect 35348 42220 35400 42226
rect 35348 42162 35400 42168
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 35360 41614 35388 42162
rect 35452 41818 35480 43114
rect 35532 42356 35584 42362
rect 35532 42298 35584 42304
rect 35440 41812 35492 41818
rect 35440 41754 35492 41760
rect 35544 41750 35572 42298
rect 35532 41744 35584 41750
rect 35532 41686 35584 41692
rect 35348 41608 35400 41614
rect 35348 41550 35400 41556
rect 34520 41064 34572 41070
rect 34520 41006 34572 41012
rect 34796 41064 34848 41070
rect 34796 41006 34848 41012
rect 34428 40588 34480 40594
rect 34428 40530 34480 40536
rect 34808 38894 34836 41006
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 35348 38956 35400 38962
rect 35348 38898 35400 38904
rect 34796 38888 34848 38894
rect 34796 38830 34848 38836
rect 34704 38752 34756 38758
rect 34704 38694 34756 38700
rect 34716 38350 34744 38694
rect 34704 38344 34756 38350
rect 34704 38286 34756 38292
rect 34428 38276 34480 38282
rect 34428 38218 34480 38224
rect 34296 38156 34376 38162
rect 34244 38150 34376 38156
rect 33888 37874 33916 38150
rect 34256 38134 34376 38150
rect 34152 37936 34204 37942
rect 34152 37878 34204 37884
rect 33876 37868 33928 37874
rect 33876 37810 33928 37816
rect 33876 37256 33928 37262
rect 33876 37198 33928 37204
rect 33600 37188 33652 37194
rect 33600 37130 33652 37136
rect 33612 36786 33640 37130
rect 33888 36922 33916 37198
rect 34164 37126 34192 37878
rect 34348 37874 34376 38134
rect 34336 37868 34388 37874
rect 34336 37810 34388 37816
rect 34152 37120 34204 37126
rect 34152 37062 34204 37068
rect 33692 36916 33744 36922
rect 33692 36858 33744 36864
rect 33876 36916 33928 36922
rect 33876 36858 33928 36864
rect 33600 36780 33652 36786
rect 33600 36722 33652 36728
rect 33704 35698 33732 36858
rect 34440 36310 34468 38218
rect 34704 37664 34756 37670
rect 34704 37606 34756 37612
rect 34716 37194 34744 37606
rect 34808 37262 34836 38830
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 35360 38554 35388 38898
rect 35440 38752 35492 38758
rect 35440 38694 35492 38700
rect 35348 38548 35400 38554
rect 35348 38490 35400 38496
rect 35452 38418 35480 38694
rect 35440 38412 35492 38418
rect 35440 38354 35492 38360
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34796 37256 34848 37262
rect 34796 37198 34848 37204
rect 34704 37188 34756 37194
rect 34704 37130 34756 37136
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34428 36304 34480 36310
rect 34428 36246 34480 36252
rect 33876 36168 33928 36174
rect 33876 36110 33928 36116
rect 33692 35692 33744 35698
rect 33692 35634 33744 35640
rect 33888 35630 33916 36110
rect 33876 35624 33928 35630
rect 33876 35566 33928 35572
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 33508 32836 33560 32842
rect 33508 32778 33560 32784
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 32864 30252 32916 30258
rect 32864 30194 32916 30200
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 33416 29164 33468 29170
rect 33416 29106 33468 29112
rect 32128 28756 32180 28762
rect 32128 28698 32180 28704
rect 32140 28082 32168 28698
rect 32128 28076 32180 28082
rect 32128 28018 32180 28024
rect 32772 27464 32824 27470
rect 32772 27406 32824 27412
rect 32128 27328 32180 27334
rect 32128 27270 32180 27276
rect 32140 27130 32168 27270
rect 32128 27124 32180 27130
rect 32128 27066 32180 27072
rect 31944 26512 31996 26518
rect 31944 26454 31996 26460
rect 31956 26382 31984 26454
rect 31944 26376 31996 26382
rect 31944 26318 31996 26324
rect 32140 25906 32168 27066
rect 32784 26926 32812 27406
rect 32404 26920 32456 26926
rect 32404 26862 32456 26868
rect 32772 26920 32824 26926
rect 32772 26862 32824 26868
rect 32128 25900 32180 25906
rect 32128 25842 32180 25848
rect 32220 25900 32272 25906
rect 32220 25842 32272 25848
rect 31852 23656 31904 23662
rect 31852 23598 31904 23604
rect 31864 22982 31892 23598
rect 31852 22976 31904 22982
rect 31852 22918 31904 22924
rect 31760 22772 31812 22778
rect 31760 22714 31812 22720
rect 31852 22568 31904 22574
rect 31852 22510 31904 22516
rect 31864 21894 31892 22510
rect 31852 21888 31904 21894
rect 31852 21830 31904 21836
rect 31944 20868 31996 20874
rect 31944 20810 31996 20816
rect 31668 20460 31720 20466
rect 31668 20402 31720 20408
rect 31484 19372 31536 19378
rect 31484 19314 31536 19320
rect 31496 18970 31524 19314
rect 31576 19304 31628 19310
rect 31576 19246 31628 19252
rect 31588 18970 31616 19246
rect 31484 18964 31536 18970
rect 31484 18906 31536 18912
rect 31576 18964 31628 18970
rect 31576 18906 31628 18912
rect 31300 18896 31352 18902
rect 31300 18838 31352 18844
rect 31208 18828 31260 18834
rect 31208 18770 31260 18776
rect 31116 18692 31168 18698
rect 31116 18634 31168 18640
rect 31024 17672 31076 17678
rect 31024 17614 31076 17620
rect 30932 17128 30984 17134
rect 30932 17070 30984 17076
rect 30840 15700 30892 15706
rect 30840 15642 30892 15648
rect 30944 15570 30972 17070
rect 31036 16114 31064 17614
rect 31024 16108 31076 16114
rect 31024 16050 31076 16056
rect 30932 15564 30984 15570
rect 30932 15506 30984 15512
rect 31024 14068 31076 14074
rect 31024 14010 31076 14016
rect 31036 13326 31064 14010
rect 30748 13320 30800 13326
rect 30748 13262 30800 13268
rect 31024 13320 31076 13326
rect 31024 13262 31076 13268
rect 31128 13258 31156 18634
rect 31392 17672 31444 17678
rect 31496 17660 31524 18906
rect 31760 18148 31812 18154
rect 31760 18090 31812 18096
rect 31772 17678 31800 18090
rect 31852 18080 31904 18086
rect 31852 18022 31904 18028
rect 31444 17632 31524 17660
rect 31760 17672 31812 17678
rect 31392 17614 31444 17620
rect 31760 17614 31812 17620
rect 31404 16182 31432 17614
rect 31484 16448 31536 16454
rect 31484 16390 31536 16396
rect 31392 16176 31444 16182
rect 31392 16118 31444 16124
rect 31496 16114 31524 16390
rect 31484 16108 31536 16114
rect 31484 16050 31536 16056
rect 31484 14408 31536 14414
rect 31484 14350 31536 14356
rect 31576 14408 31628 14414
rect 31576 14350 31628 14356
rect 31116 13252 31168 13258
rect 31116 13194 31168 13200
rect 28644 12406 28856 12434
rect 28630 11792 28686 11801
rect 28828 11762 28856 12406
rect 30012 11892 30064 11898
rect 30012 11834 30064 11840
rect 28630 11727 28632 11736
rect 28684 11727 28686 11736
rect 28816 11756 28868 11762
rect 28632 11698 28684 11704
rect 28816 11698 28868 11704
rect 29000 11756 29052 11762
rect 29000 11698 29052 11704
rect 29092 11756 29144 11762
rect 29092 11698 29144 11704
rect 29736 11756 29788 11762
rect 29736 11698 29788 11704
rect 29920 11756 29972 11762
rect 29920 11698 29972 11704
rect 28724 11212 28776 11218
rect 28724 11154 28776 11160
rect 28736 9994 28764 11154
rect 28828 10606 28856 11698
rect 29012 11354 29040 11698
rect 29000 11348 29052 11354
rect 29000 11290 29052 11296
rect 29000 10668 29052 10674
rect 29104 10656 29132 11698
rect 29748 11150 29776 11698
rect 29184 11144 29236 11150
rect 29184 11086 29236 11092
rect 29736 11144 29788 11150
rect 29736 11086 29788 11092
rect 29196 10674 29224 11086
rect 29052 10628 29132 10656
rect 29000 10610 29052 10616
rect 28816 10600 28868 10606
rect 28816 10542 28868 10548
rect 28908 10532 28960 10538
rect 28908 10474 28960 10480
rect 28724 9988 28776 9994
rect 28724 9930 28776 9936
rect 28920 9382 28948 10474
rect 29000 10464 29052 10470
rect 29000 10406 29052 10412
rect 29012 9586 29040 10406
rect 29104 10266 29132 10628
rect 29184 10668 29236 10674
rect 29184 10610 29236 10616
rect 29748 10606 29776 11086
rect 29932 11082 29960 11698
rect 30024 11150 30052 11834
rect 30656 11756 30708 11762
rect 30656 11698 30708 11704
rect 30012 11144 30064 11150
rect 30012 11086 30064 11092
rect 29920 11076 29972 11082
rect 29920 11018 29972 11024
rect 30564 11008 30616 11014
rect 30564 10950 30616 10956
rect 30576 10674 30604 10950
rect 30668 10810 30696 11698
rect 31496 11336 31524 14350
rect 31588 14074 31616 14350
rect 31864 14226 31892 18022
rect 31956 14414 31984 20810
rect 32036 19712 32088 19718
rect 32036 19654 32088 19660
rect 32048 19378 32076 19654
rect 32036 19372 32088 19378
rect 32036 19314 32088 19320
rect 31944 14408 31996 14414
rect 31944 14350 31996 14356
rect 32036 14272 32088 14278
rect 31864 14198 31984 14226
rect 32036 14214 32088 14220
rect 31576 14068 31628 14074
rect 31576 14010 31628 14016
rect 31760 12232 31812 12238
rect 31760 12174 31812 12180
rect 31668 11348 31720 11354
rect 31496 11308 31668 11336
rect 30656 10804 30708 10810
rect 30656 10746 30708 10752
rect 30932 10804 30984 10810
rect 30932 10746 30984 10752
rect 30944 10674 30972 10746
rect 31496 10742 31524 11308
rect 31668 11290 31720 11296
rect 31772 11150 31800 12174
rect 31956 11898 31984 14198
rect 31944 11892 31996 11898
rect 31944 11834 31996 11840
rect 32048 11762 32076 14214
rect 32036 11756 32088 11762
rect 32036 11698 32088 11704
rect 31852 11688 31904 11694
rect 31852 11630 31904 11636
rect 31760 11144 31812 11150
rect 31760 11086 31812 11092
rect 31484 10736 31536 10742
rect 31484 10678 31536 10684
rect 30564 10668 30616 10674
rect 30564 10610 30616 10616
rect 30932 10668 30984 10674
rect 30932 10610 30984 10616
rect 29736 10600 29788 10606
rect 29736 10542 29788 10548
rect 29920 10600 29972 10606
rect 29920 10542 29972 10548
rect 29828 10464 29880 10470
rect 29828 10406 29880 10412
rect 29092 10260 29144 10266
rect 29092 10202 29144 10208
rect 29736 10124 29788 10130
rect 29736 10066 29788 10072
rect 29184 9988 29236 9994
rect 29184 9930 29236 9936
rect 29196 9738 29224 9930
rect 29104 9710 29224 9738
rect 29104 9654 29132 9710
rect 29092 9648 29144 9654
rect 29092 9590 29144 9596
rect 29000 9580 29052 9586
rect 29000 9522 29052 9528
rect 29748 9382 29776 10066
rect 29840 9722 29868 10406
rect 29932 10266 29960 10542
rect 29920 10260 29972 10266
rect 29920 10202 29972 10208
rect 30840 10192 30892 10198
rect 30840 10134 30892 10140
rect 30196 10056 30248 10062
rect 30196 9998 30248 10004
rect 29828 9716 29880 9722
rect 29828 9658 29880 9664
rect 29840 9518 29868 9658
rect 30208 9654 30236 9998
rect 30852 9994 30880 10134
rect 30840 9988 30892 9994
rect 30840 9930 30892 9936
rect 31392 9988 31444 9994
rect 31392 9930 31444 9936
rect 30196 9648 30248 9654
rect 30196 9590 30248 9596
rect 29828 9512 29880 9518
rect 29828 9454 29880 9460
rect 31404 9382 31432 9930
rect 31864 9450 31892 11630
rect 32128 11552 32180 11558
rect 32128 11494 32180 11500
rect 32140 11286 32168 11494
rect 32128 11280 32180 11286
rect 32128 11222 32180 11228
rect 31944 10532 31996 10538
rect 31944 10474 31996 10480
rect 31956 10062 31984 10474
rect 32128 10464 32180 10470
rect 32128 10406 32180 10412
rect 32036 10192 32088 10198
rect 32036 10134 32088 10140
rect 31944 10056 31996 10062
rect 31944 9998 31996 10004
rect 31852 9444 31904 9450
rect 31852 9386 31904 9392
rect 28908 9376 28960 9382
rect 28908 9318 28960 9324
rect 29736 9376 29788 9382
rect 29736 9318 29788 9324
rect 31392 9376 31444 9382
rect 31392 9318 31444 9324
rect 31956 8974 31984 9998
rect 32048 9586 32076 10134
rect 32036 9580 32088 9586
rect 32036 9522 32088 9528
rect 32048 9382 32076 9522
rect 32036 9376 32088 9382
rect 32036 9318 32088 9324
rect 32048 9178 32076 9318
rect 32036 9172 32088 9178
rect 32036 9114 32088 9120
rect 32140 8974 32168 10406
rect 31944 8968 31996 8974
rect 31944 8910 31996 8916
rect 32128 8968 32180 8974
rect 32128 8910 32180 8916
rect 32232 8430 32260 25842
rect 32416 25702 32444 26862
rect 32784 26450 32812 26862
rect 32772 26444 32824 26450
rect 32772 26386 32824 26392
rect 32496 25968 32548 25974
rect 32496 25910 32548 25916
rect 32404 25696 32456 25702
rect 32404 25638 32456 25644
rect 32416 23866 32444 25638
rect 32508 25498 32536 25910
rect 32496 25492 32548 25498
rect 32496 25434 32548 25440
rect 32508 24954 32536 25434
rect 32496 24948 32548 24954
rect 32496 24890 32548 24896
rect 32784 24818 33180 24834
rect 32772 24812 33192 24818
rect 32824 24806 33140 24812
rect 32772 24754 32824 24760
rect 33140 24754 33192 24760
rect 32772 24608 32824 24614
rect 32772 24550 32824 24556
rect 32588 24132 32640 24138
rect 32588 24074 32640 24080
rect 32600 23866 32628 24074
rect 32404 23860 32456 23866
rect 32404 23802 32456 23808
rect 32588 23860 32640 23866
rect 32588 23802 32640 23808
rect 32784 23730 32812 24550
rect 32772 23724 32824 23730
rect 32772 23666 32824 23672
rect 33140 23588 33192 23594
rect 33140 23530 33192 23536
rect 33152 22574 33180 23530
rect 33140 22568 33192 22574
rect 33140 22510 33192 22516
rect 32864 22500 32916 22506
rect 32864 22442 32916 22448
rect 32680 22432 32732 22438
rect 32680 22374 32732 22380
rect 32494 21312 32550 21321
rect 32494 21247 32550 21256
rect 32508 19854 32536 21247
rect 32692 20942 32720 22374
rect 32876 20942 32904 22442
rect 33152 22166 33180 22510
rect 33140 22160 33192 22166
rect 33140 22102 33192 22108
rect 33428 22030 33456 29106
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 33600 27464 33652 27470
rect 33600 27406 33652 27412
rect 34888 27464 34940 27470
rect 34888 27406 34940 27412
rect 35072 27464 35124 27470
rect 35072 27406 35124 27412
rect 33508 27328 33560 27334
rect 33508 27270 33560 27276
rect 33520 26994 33548 27270
rect 33508 26988 33560 26994
rect 33508 26930 33560 26936
rect 33612 26042 33640 27406
rect 34900 27130 34928 27406
rect 34888 27124 34940 27130
rect 34888 27066 34940 27072
rect 35084 26994 35112 27406
rect 34612 26988 34664 26994
rect 34612 26930 34664 26936
rect 35072 26988 35124 26994
rect 35072 26930 35124 26936
rect 34624 26790 34652 26930
rect 34612 26784 34664 26790
rect 34612 26726 34664 26732
rect 33784 26308 33836 26314
rect 33784 26250 33836 26256
rect 33600 26036 33652 26042
rect 33600 25978 33652 25984
rect 33508 25764 33560 25770
rect 33508 25706 33560 25712
rect 33520 22710 33548 25706
rect 33796 25294 33824 26250
rect 34624 25906 34652 26726
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35440 26240 35492 26246
rect 35440 26182 35492 26188
rect 35452 26042 35480 26182
rect 35440 26036 35492 26042
rect 35440 25978 35492 25984
rect 34612 25900 34664 25906
rect 34612 25842 34664 25848
rect 34244 25832 34296 25838
rect 34244 25774 34296 25780
rect 35440 25832 35492 25838
rect 35440 25774 35492 25780
rect 33784 25288 33836 25294
rect 33784 25230 33836 25236
rect 33796 24206 33824 25230
rect 34152 25152 34204 25158
rect 34152 25094 34204 25100
rect 33876 24812 33928 24818
rect 33876 24754 33928 24760
rect 34060 24812 34112 24818
rect 34060 24754 34112 24760
rect 33888 24206 33916 24754
rect 33968 24744 34020 24750
rect 33968 24686 34020 24692
rect 33784 24200 33836 24206
rect 33784 24142 33836 24148
rect 33876 24200 33928 24206
rect 33876 24142 33928 24148
rect 33796 23730 33824 24142
rect 33784 23724 33836 23730
rect 33784 23666 33836 23672
rect 33876 23724 33928 23730
rect 33876 23666 33928 23672
rect 33692 22976 33744 22982
rect 33692 22918 33744 22924
rect 33508 22704 33560 22710
rect 33508 22646 33560 22652
rect 33704 22642 33732 22918
rect 33692 22636 33744 22642
rect 33692 22578 33744 22584
rect 33416 22024 33468 22030
rect 33416 21966 33468 21972
rect 33796 21622 33824 23666
rect 33888 22778 33916 23666
rect 33980 23118 34008 24686
rect 34072 24342 34100 24754
rect 34060 24336 34112 24342
rect 34060 24278 34112 24284
rect 34060 24200 34112 24206
rect 34060 24142 34112 24148
rect 34072 23526 34100 24142
rect 34060 23520 34112 23526
rect 34060 23462 34112 23468
rect 34072 23118 34100 23462
rect 33968 23112 34020 23118
rect 33968 23054 34020 23060
rect 34060 23112 34112 23118
rect 34060 23054 34112 23060
rect 33876 22772 33928 22778
rect 33876 22714 33928 22720
rect 33980 22658 34008 23054
rect 33888 22630 34008 22658
rect 33888 22030 33916 22630
rect 33968 22228 34020 22234
rect 33968 22170 34020 22176
rect 33876 22024 33928 22030
rect 33876 21966 33928 21972
rect 33980 21622 34008 22170
rect 34072 22030 34100 23054
rect 34060 22024 34112 22030
rect 34060 21966 34112 21972
rect 33784 21616 33836 21622
rect 33784 21558 33836 21564
rect 33968 21616 34020 21622
rect 33968 21558 34020 21564
rect 32956 21548 33008 21554
rect 32956 21490 33008 21496
rect 33140 21548 33192 21554
rect 33140 21490 33192 21496
rect 33232 21548 33284 21554
rect 33232 21490 33284 21496
rect 32968 21350 32996 21490
rect 32956 21344 33008 21350
rect 32956 21286 33008 21292
rect 32680 20936 32732 20942
rect 32680 20878 32732 20884
rect 32864 20936 32916 20942
rect 32864 20878 32916 20884
rect 32680 20052 32732 20058
rect 32680 19994 32732 20000
rect 32496 19848 32548 19854
rect 32496 19790 32548 19796
rect 32692 19514 32720 19994
rect 32876 19854 32904 20878
rect 32968 19922 32996 21286
rect 33152 20602 33180 21490
rect 33244 21146 33272 21490
rect 33232 21140 33284 21146
rect 33232 21082 33284 21088
rect 34164 20942 34192 25094
rect 34256 22098 34284 25774
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35348 23520 35400 23526
rect 35348 23462 35400 23468
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 35360 23118 35388 23462
rect 35348 23112 35400 23118
rect 35348 23054 35400 23060
rect 35360 22710 35388 23054
rect 35348 22704 35400 22710
rect 35348 22646 35400 22652
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34244 22092 34296 22098
rect 34244 22034 34296 22040
rect 34256 21078 34284 22034
rect 35072 22024 35124 22030
rect 35072 21966 35124 21972
rect 35084 21418 35112 21966
rect 35072 21412 35124 21418
rect 35072 21354 35124 21360
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34244 21072 34296 21078
rect 34244 21014 34296 21020
rect 33692 20936 33744 20942
rect 33692 20878 33744 20884
rect 34152 20936 34204 20942
rect 34152 20878 34204 20884
rect 33140 20596 33192 20602
rect 33140 20538 33192 20544
rect 33704 20466 33732 20878
rect 33876 20868 33928 20874
rect 33876 20810 33928 20816
rect 33888 20466 33916 20810
rect 33692 20460 33744 20466
rect 33692 20402 33744 20408
rect 33876 20460 33928 20466
rect 33876 20402 33928 20408
rect 34520 20460 34572 20466
rect 34520 20402 34572 20408
rect 33704 20058 33732 20402
rect 33888 20346 33916 20402
rect 33888 20318 34008 20346
rect 33876 20256 33928 20262
rect 33876 20198 33928 20204
rect 33692 20052 33744 20058
rect 33692 19994 33744 20000
rect 32956 19916 33008 19922
rect 32956 19858 33008 19864
rect 32864 19848 32916 19854
rect 32864 19790 32916 19796
rect 32864 19712 32916 19718
rect 32864 19654 32916 19660
rect 32680 19508 32732 19514
rect 32680 19450 32732 19456
rect 32496 16992 32548 16998
rect 32496 16934 32548 16940
rect 32404 16516 32456 16522
rect 32404 16458 32456 16464
rect 32416 16250 32444 16458
rect 32404 16244 32456 16250
rect 32404 16186 32456 16192
rect 32508 16114 32536 16934
rect 32692 16114 32720 19450
rect 32876 19446 32904 19654
rect 32864 19440 32916 19446
rect 32864 19382 32916 19388
rect 33692 19372 33744 19378
rect 33692 19314 33744 19320
rect 33600 19236 33652 19242
rect 33600 19178 33652 19184
rect 33140 18828 33192 18834
rect 33140 18770 33192 18776
rect 33152 18222 33180 18770
rect 33612 18426 33640 19178
rect 33704 18698 33732 19314
rect 33784 18828 33836 18834
rect 33784 18770 33836 18776
rect 33692 18692 33744 18698
rect 33692 18634 33744 18640
rect 33600 18420 33652 18426
rect 33600 18362 33652 18368
rect 32956 18216 33008 18222
rect 32956 18158 33008 18164
rect 33140 18216 33192 18222
rect 33140 18158 33192 18164
rect 33324 18216 33376 18222
rect 33324 18158 33376 18164
rect 32968 17882 32996 18158
rect 33336 18086 33364 18158
rect 33324 18080 33376 18086
rect 33324 18022 33376 18028
rect 32956 17876 33008 17882
rect 32956 17818 33008 17824
rect 33324 17196 33376 17202
rect 33324 17138 33376 17144
rect 33336 16726 33364 17138
rect 33704 17134 33732 18634
rect 33796 18340 33824 18770
rect 33888 18766 33916 20198
rect 33980 19990 34008 20318
rect 34152 20052 34204 20058
rect 34152 19994 34204 20000
rect 34244 20052 34296 20058
rect 34244 19994 34296 20000
rect 33968 19984 34020 19990
rect 33968 19926 34020 19932
rect 33980 19378 34008 19926
rect 33968 19372 34020 19378
rect 33968 19314 34020 19320
rect 34164 19174 34192 19994
rect 34256 19718 34284 19994
rect 34532 19854 34560 20402
rect 34796 20392 34848 20398
rect 34796 20334 34848 20340
rect 34520 19848 34572 19854
rect 34520 19790 34572 19796
rect 34244 19712 34296 19718
rect 34244 19654 34296 19660
rect 34152 19168 34204 19174
rect 34152 19110 34204 19116
rect 34428 19168 34480 19174
rect 34428 19110 34480 19116
rect 34152 18964 34204 18970
rect 34152 18906 34204 18912
rect 33876 18760 33928 18766
rect 33876 18702 33928 18708
rect 33968 18624 34020 18630
rect 33968 18566 34020 18572
rect 33876 18352 33928 18358
rect 33796 18312 33876 18340
rect 33876 18294 33928 18300
rect 33980 18086 34008 18566
rect 34060 18284 34112 18290
rect 34060 18226 34112 18232
rect 33968 18080 34020 18086
rect 33968 18022 34020 18028
rect 34072 17882 34100 18226
rect 34164 18154 34192 18906
rect 34440 18834 34468 19110
rect 34520 18896 34572 18902
rect 34520 18838 34572 18844
rect 34428 18828 34480 18834
rect 34428 18770 34480 18776
rect 34152 18148 34204 18154
rect 34152 18090 34204 18096
rect 34060 17876 34112 17882
rect 34060 17818 34112 17824
rect 33692 17128 33744 17134
rect 33692 17070 33744 17076
rect 34072 17066 34100 17818
rect 34532 17354 34560 18838
rect 34808 18834 34836 20334
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35452 20058 35480 25774
rect 35636 21690 35664 45426
rect 40604 44946 40632 45426
rect 40592 44940 40644 44946
rect 40592 44882 40644 44888
rect 40040 44872 40092 44878
rect 40040 44814 40092 44820
rect 40052 44334 40080 44814
rect 40040 44328 40092 44334
rect 40040 44270 40092 44276
rect 36544 43852 36596 43858
rect 36544 43794 36596 43800
rect 36556 43314 36584 43794
rect 36544 43308 36596 43314
rect 36544 43250 36596 43256
rect 35716 42220 35768 42226
rect 35716 42162 35768 42168
rect 35728 41682 35756 42162
rect 35716 41676 35768 41682
rect 35716 41618 35768 41624
rect 36636 37256 36688 37262
rect 36636 37198 36688 37204
rect 35900 33516 35952 33522
rect 35900 33458 35952 33464
rect 35912 28558 35940 33458
rect 36648 33454 36676 37198
rect 36636 33448 36688 33454
rect 36636 33390 36688 33396
rect 36648 32502 36676 33390
rect 36636 32496 36688 32502
rect 36636 32438 36688 32444
rect 40604 31754 40632 44882
rect 40604 31726 40816 31754
rect 38016 29164 38068 29170
rect 38016 29106 38068 29112
rect 35900 28552 35952 28558
rect 35900 28494 35952 28500
rect 35716 27464 35768 27470
rect 35716 27406 35768 27412
rect 35728 27130 35756 27406
rect 35808 27328 35860 27334
rect 35808 27270 35860 27276
rect 35716 27124 35768 27130
rect 35716 27066 35768 27072
rect 35716 26444 35768 26450
rect 35716 26386 35768 26392
rect 35728 24818 35756 26386
rect 35820 26382 35848 27270
rect 35912 26518 35940 28494
rect 36176 27464 36228 27470
rect 36176 27406 36228 27412
rect 36188 26790 36216 27406
rect 36452 27396 36504 27402
rect 36452 27338 36504 27344
rect 36176 26784 36228 26790
rect 36176 26726 36228 26732
rect 35900 26512 35952 26518
rect 35900 26454 35952 26460
rect 35808 26376 35860 26382
rect 35808 26318 35860 26324
rect 36084 26376 36136 26382
rect 36084 26318 36136 26324
rect 35992 26308 36044 26314
rect 35992 26250 36044 26256
rect 36004 24818 36032 26250
rect 36096 25974 36124 26318
rect 36188 25974 36216 26726
rect 36084 25968 36136 25974
rect 36084 25910 36136 25916
rect 36176 25968 36228 25974
rect 36176 25910 36228 25916
rect 35716 24812 35768 24818
rect 35716 24754 35768 24760
rect 35992 24812 36044 24818
rect 35992 24754 36044 24760
rect 36004 24274 36032 24754
rect 36096 24750 36124 25910
rect 36188 25362 36216 25910
rect 36464 25362 36492 27338
rect 38028 26994 38056 29106
rect 38476 29028 38528 29034
rect 38476 28970 38528 28976
rect 38108 28484 38160 28490
rect 38108 28426 38160 28432
rect 38120 27470 38148 28426
rect 38108 27464 38160 27470
rect 38108 27406 38160 27412
rect 37648 26988 37700 26994
rect 37648 26930 37700 26936
rect 38016 26988 38068 26994
rect 38016 26930 38068 26936
rect 37660 26382 37688 26930
rect 36544 26376 36596 26382
rect 36544 26318 36596 26324
rect 37648 26376 37700 26382
rect 37648 26318 37700 26324
rect 36556 25770 36584 26318
rect 38120 25838 38148 27406
rect 38384 27056 38436 27062
rect 38384 26998 38436 27004
rect 38396 26382 38424 26998
rect 38488 26466 38516 28970
rect 38568 27396 38620 27402
rect 38568 27338 38620 27344
rect 38580 27130 38608 27338
rect 39488 27328 39540 27334
rect 39488 27270 39540 27276
rect 38568 27124 38620 27130
rect 38568 27066 38620 27072
rect 39500 26994 39528 27270
rect 38936 26988 38988 26994
rect 38936 26930 38988 26936
rect 39488 26988 39540 26994
rect 39488 26930 39540 26936
rect 38844 26784 38896 26790
rect 38844 26726 38896 26732
rect 38856 26518 38884 26726
rect 38844 26512 38896 26518
rect 38488 26438 38608 26466
rect 38844 26454 38896 26460
rect 38580 26382 38608 26438
rect 38292 26376 38344 26382
rect 38292 26318 38344 26324
rect 38384 26376 38436 26382
rect 38384 26318 38436 26324
rect 38568 26376 38620 26382
rect 38568 26318 38620 26324
rect 38304 25906 38332 26318
rect 38396 25906 38424 26318
rect 38292 25900 38344 25906
rect 38292 25842 38344 25848
rect 38384 25900 38436 25906
rect 38384 25842 38436 25848
rect 38568 25900 38620 25906
rect 38568 25842 38620 25848
rect 38752 25900 38804 25906
rect 38752 25842 38804 25848
rect 37280 25832 37332 25838
rect 37280 25774 37332 25780
rect 38108 25832 38160 25838
rect 38108 25774 38160 25780
rect 36544 25764 36596 25770
rect 36544 25706 36596 25712
rect 36728 25764 36780 25770
rect 36728 25706 36780 25712
rect 36176 25356 36228 25362
rect 36176 25298 36228 25304
rect 36452 25356 36504 25362
rect 36452 25298 36504 25304
rect 36360 25288 36412 25294
rect 36360 25230 36412 25236
rect 36372 24886 36400 25230
rect 36452 25220 36504 25226
rect 36452 25162 36504 25168
rect 36360 24880 36412 24886
rect 36360 24822 36412 24828
rect 36464 24818 36492 25162
rect 36740 24818 36768 25706
rect 36912 25696 36964 25702
rect 36912 25638 36964 25644
rect 36924 25294 36952 25638
rect 37292 25294 37320 25774
rect 38200 25696 38252 25702
rect 38200 25638 38252 25644
rect 36912 25288 36964 25294
rect 36912 25230 36964 25236
rect 37280 25288 37332 25294
rect 37280 25230 37332 25236
rect 36452 24812 36504 24818
rect 36452 24754 36504 24760
rect 36728 24812 36780 24818
rect 36728 24754 36780 24760
rect 36084 24744 36136 24750
rect 36084 24686 36136 24692
rect 36360 24608 36412 24614
rect 36360 24550 36412 24556
rect 35992 24268 36044 24274
rect 35992 24210 36044 24216
rect 36372 24206 36400 24550
rect 36360 24200 36412 24206
rect 36360 24142 36412 24148
rect 36464 24070 36492 24754
rect 36452 24064 36504 24070
rect 36452 24006 36504 24012
rect 36464 23730 36492 24006
rect 36452 23724 36504 23730
rect 36452 23666 36504 23672
rect 36268 23112 36320 23118
rect 36268 23054 36320 23060
rect 35808 22976 35860 22982
rect 35808 22918 35860 22924
rect 35820 22642 35848 22918
rect 35808 22636 35860 22642
rect 35808 22578 35860 22584
rect 35900 22636 35952 22642
rect 35900 22578 35952 22584
rect 35912 22098 35940 22578
rect 36084 22568 36136 22574
rect 36084 22510 36136 22516
rect 36176 22568 36228 22574
rect 36176 22510 36228 22516
rect 35900 22092 35952 22098
rect 35900 22034 35952 22040
rect 35624 21684 35676 21690
rect 35624 21626 35676 21632
rect 35624 20596 35676 20602
rect 35624 20538 35676 20544
rect 35636 20330 35664 20538
rect 35624 20324 35676 20330
rect 35624 20266 35676 20272
rect 35440 20052 35492 20058
rect 35440 19994 35492 20000
rect 35440 19916 35492 19922
rect 35440 19858 35492 19864
rect 35348 19712 35400 19718
rect 35348 19654 35400 19660
rect 35360 19378 35388 19654
rect 35348 19372 35400 19378
rect 35348 19314 35400 19320
rect 35256 19304 35308 19310
rect 35452 19258 35480 19858
rect 35624 19780 35676 19786
rect 35624 19722 35676 19728
rect 35532 19440 35584 19446
rect 35532 19382 35584 19388
rect 35308 19252 35480 19258
rect 35256 19246 35480 19252
rect 35268 19230 35480 19246
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35452 18970 35480 19230
rect 35544 18970 35572 19382
rect 35440 18964 35492 18970
rect 35440 18906 35492 18912
rect 35532 18964 35584 18970
rect 35532 18906 35584 18912
rect 35636 18834 35664 19722
rect 35716 19712 35768 19718
rect 35716 19654 35768 19660
rect 35728 19514 35756 19654
rect 35716 19508 35768 19514
rect 35716 19450 35768 19456
rect 35808 19440 35860 19446
rect 35808 19382 35860 19388
rect 34796 18828 34848 18834
rect 34796 18770 34848 18776
rect 35624 18828 35676 18834
rect 35624 18770 35676 18776
rect 35820 18766 35848 19382
rect 35912 19310 35940 22034
rect 36096 21894 36124 22510
rect 36084 21888 36136 21894
rect 36084 21830 36136 21836
rect 36188 21554 36216 22510
rect 36176 21548 36228 21554
rect 36176 21490 36228 21496
rect 36280 21350 36308 23054
rect 36464 23050 36492 23666
rect 36544 23520 36596 23526
rect 36544 23462 36596 23468
rect 36556 23118 36584 23462
rect 36544 23112 36596 23118
rect 36544 23054 36596 23060
rect 36452 23044 36504 23050
rect 36452 22986 36504 22992
rect 36544 22432 36596 22438
rect 36544 22374 36596 22380
rect 36556 21962 36584 22374
rect 36544 21956 36596 21962
rect 36544 21898 36596 21904
rect 36740 21894 36768 24754
rect 37292 24274 37320 25230
rect 38016 25220 38068 25226
rect 38016 25162 38068 25168
rect 38028 24954 38056 25162
rect 38016 24948 38068 24954
rect 38016 24890 38068 24896
rect 37372 24880 37424 24886
rect 37372 24822 37424 24828
rect 37280 24268 37332 24274
rect 37280 24210 37332 24216
rect 37188 22160 37240 22166
rect 37188 22102 37240 22108
rect 36728 21888 36780 21894
rect 36728 21830 36780 21836
rect 37200 21554 37228 22102
rect 37292 22030 37320 24210
rect 37384 23730 37412 24822
rect 38212 24818 38240 25638
rect 38200 24812 38252 24818
rect 38200 24754 38252 24760
rect 37372 23724 37424 23730
rect 37372 23666 37424 23672
rect 37384 22982 37412 23666
rect 37372 22976 37424 22982
rect 37372 22918 37424 22924
rect 37280 22024 37332 22030
rect 37280 21966 37332 21972
rect 37188 21548 37240 21554
rect 37188 21490 37240 21496
rect 36268 21344 36320 21350
rect 36268 21286 36320 21292
rect 35992 19780 36044 19786
rect 35992 19722 36044 19728
rect 36004 19514 36032 19722
rect 35992 19508 36044 19514
rect 35992 19450 36044 19456
rect 35900 19304 35952 19310
rect 35900 19246 35952 19252
rect 35912 18902 35940 19246
rect 36280 18970 36308 21286
rect 37292 19854 37320 21966
rect 38108 21344 38160 21350
rect 38108 21286 38160 21292
rect 38120 20942 38148 21286
rect 38108 20936 38160 20942
rect 38108 20878 38160 20884
rect 38304 20806 38332 25842
rect 38476 25152 38528 25158
rect 38476 25094 38528 25100
rect 38488 24750 38516 25094
rect 38476 24744 38528 24750
rect 38476 24686 38528 24692
rect 38384 24608 38436 24614
rect 38384 24550 38436 24556
rect 37924 20800 37976 20806
rect 37924 20742 37976 20748
rect 38292 20800 38344 20806
rect 38292 20742 38344 20748
rect 37740 20460 37792 20466
rect 37740 20402 37792 20408
rect 37752 20058 37780 20402
rect 37740 20052 37792 20058
rect 37740 19994 37792 20000
rect 37936 19854 37964 20742
rect 38200 20256 38252 20262
rect 38200 20198 38252 20204
rect 38212 19922 38240 20198
rect 38200 19916 38252 19922
rect 38200 19858 38252 19864
rect 37280 19848 37332 19854
rect 37280 19790 37332 19796
rect 37924 19848 37976 19854
rect 37924 19790 37976 19796
rect 37464 19712 37516 19718
rect 37464 19654 37516 19660
rect 37476 19446 37504 19654
rect 38212 19446 38240 19858
rect 38396 19786 38424 24550
rect 38476 22636 38528 22642
rect 38476 22578 38528 22584
rect 38488 22030 38516 22578
rect 38476 22024 38528 22030
rect 38476 21966 38528 21972
rect 38580 21350 38608 25842
rect 38764 22778 38792 25842
rect 38856 24614 38884 26454
rect 38844 24608 38896 24614
rect 38844 24550 38896 24556
rect 38752 22772 38804 22778
rect 38752 22714 38804 22720
rect 38948 22642 38976 26930
rect 40684 26376 40736 26382
rect 40684 26318 40736 26324
rect 39028 26240 39080 26246
rect 39028 26182 39080 26188
rect 39040 25974 39068 26182
rect 40696 26042 40724 26318
rect 40684 26036 40736 26042
rect 40604 25996 40684 26024
rect 39028 25968 39080 25974
rect 39028 25910 39080 25916
rect 39764 24336 39816 24342
rect 39764 24278 39816 24284
rect 39396 24200 39448 24206
rect 39396 24142 39448 24148
rect 39408 23866 39436 24142
rect 39776 23866 39804 24278
rect 39396 23860 39448 23866
rect 39396 23802 39448 23808
rect 39764 23860 39816 23866
rect 39764 23802 39816 23808
rect 39948 23656 40000 23662
rect 39948 23598 40000 23604
rect 39120 23112 39172 23118
rect 39120 23054 39172 23060
rect 39396 23112 39448 23118
rect 39396 23054 39448 23060
rect 39132 22710 39160 23054
rect 39120 22704 39172 22710
rect 39120 22646 39172 22652
rect 38936 22636 38988 22642
rect 38936 22578 38988 22584
rect 39304 22636 39356 22642
rect 39304 22578 39356 22584
rect 39212 22568 39264 22574
rect 39212 22510 39264 22516
rect 39224 22030 39252 22510
rect 39316 22234 39344 22578
rect 39408 22234 39436 23054
rect 39580 23044 39632 23050
rect 39580 22986 39632 22992
rect 39592 22642 39620 22986
rect 39672 22772 39724 22778
rect 39672 22714 39724 22720
rect 39580 22636 39632 22642
rect 39580 22578 39632 22584
rect 39304 22228 39356 22234
rect 39304 22170 39356 22176
rect 39396 22228 39448 22234
rect 39396 22170 39448 22176
rect 39684 22094 39712 22714
rect 39592 22066 39712 22094
rect 39212 22024 39264 22030
rect 39212 21966 39264 21972
rect 39488 21888 39540 21894
rect 39488 21830 39540 21836
rect 39500 21554 39528 21830
rect 39488 21548 39540 21554
rect 39488 21490 39540 21496
rect 38568 21344 38620 21350
rect 38568 21286 38620 21292
rect 38936 21344 38988 21350
rect 38936 21286 38988 21292
rect 38752 20868 38804 20874
rect 38752 20810 38804 20816
rect 38384 19780 38436 19786
rect 38384 19722 38436 19728
rect 37464 19440 37516 19446
rect 37464 19382 37516 19388
rect 38200 19440 38252 19446
rect 38200 19382 38252 19388
rect 36636 19168 36688 19174
rect 36636 19110 36688 19116
rect 36268 18964 36320 18970
rect 36268 18906 36320 18912
rect 35900 18896 35952 18902
rect 35900 18838 35952 18844
rect 35808 18760 35860 18766
rect 35808 18702 35860 18708
rect 36648 18698 36676 19110
rect 38292 18964 38344 18970
rect 38292 18906 38344 18912
rect 37188 18896 37240 18902
rect 37188 18838 37240 18844
rect 34888 18692 34940 18698
rect 34888 18634 34940 18640
rect 36636 18692 36688 18698
rect 36636 18634 36688 18640
rect 34900 18154 34928 18634
rect 35900 18624 35952 18630
rect 35900 18566 35952 18572
rect 35912 18358 35940 18566
rect 36648 18426 36676 18634
rect 36636 18420 36688 18426
rect 36636 18362 36688 18368
rect 35900 18352 35952 18358
rect 35900 18294 35952 18300
rect 34888 18148 34940 18154
rect 34888 18090 34940 18096
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35912 17882 35940 18294
rect 36452 18284 36504 18290
rect 36452 18226 36504 18232
rect 35900 17876 35952 17882
rect 35900 17818 35952 17824
rect 36464 17678 36492 18226
rect 36648 18170 36676 18362
rect 37200 18358 37228 18838
rect 37188 18352 37240 18358
rect 37188 18294 37240 18300
rect 37004 18284 37056 18290
rect 37004 18226 37056 18232
rect 36648 18142 36768 18170
rect 36636 18080 36688 18086
rect 36636 18022 36688 18028
rect 34612 17672 34664 17678
rect 34612 17614 34664 17620
rect 35992 17672 36044 17678
rect 35992 17614 36044 17620
rect 36452 17672 36504 17678
rect 36452 17614 36504 17620
rect 34440 17326 34560 17354
rect 33416 17060 33468 17066
rect 33416 17002 33468 17008
rect 34060 17060 34112 17066
rect 34060 17002 34112 17008
rect 33324 16720 33376 16726
rect 33324 16662 33376 16668
rect 33336 16454 33364 16662
rect 33324 16448 33376 16454
rect 33324 16390 33376 16396
rect 33336 16114 33364 16390
rect 33428 16114 33456 17002
rect 34440 16998 34468 17326
rect 34624 17270 34652 17614
rect 35808 17604 35860 17610
rect 35808 17546 35860 17552
rect 35348 17536 35400 17542
rect 35348 17478 35400 17484
rect 34612 17264 34664 17270
rect 34612 17206 34664 17212
rect 34796 17264 34848 17270
rect 34796 17206 34848 17212
rect 34520 17196 34572 17202
rect 34520 17138 34572 17144
rect 34428 16992 34480 16998
rect 34428 16934 34480 16940
rect 34532 16454 34560 17138
rect 34704 16992 34756 16998
rect 34704 16934 34756 16940
rect 34716 16794 34744 16934
rect 34704 16788 34756 16794
rect 34704 16730 34756 16736
rect 34716 16522 34744 16730
rect 34808 16590 34836 17206
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35072 16720 35124 16726
rect 35072 16662 35124 16668
rect 34796 16584 34848 16590
rect 34796 16526 34848 16532
rect 34704 16516 34756 16522
rect 34704 16458 34756 16464
rect 34152 16448 34204 16454
rect 34152 16390 34204 16396
rect 34520 16448 34572 16454
rect 34520 16390 34572 16396
rect 34164 16114 34192 16390
rect 32496 16108 32548 16114
rect 32496 16050 32548 16056
rect 32680 16108 32732 16114
rect 32680 16050 32732 16056
rect 33324 16108 33376 16114
rect 33324 16050 33376 16056
rect 33416 16108 33468 16114
rect 33416 16050 33468 16056
rect 33600 16108 33652 16114
rect 33600 16050 33652 16056
rect 34152 16108 34204 16114
rect 34152 16050 34204 16056
rect 33232 15904 33284 15910
rect 33232 15846 33284 15852
rect 33244 15502 33272 15846
rect 33232 15496 33284 15502
rect 33232 15438 33284 15444
rect 32680 15020 32732 15026
rect 32680 14962 32732 14968
rect 32588 14816 32640 14822
rect 32588 14758 32640 14764
rect 32496 14408 32548 14414
rect 32496 14350 32548 14356
rect 32312 13864 32364 13870
rect 32312 13806 32364 13812
rect 32324 12918 32352 13806
rect 32508 13394 32536 14350
rect 32600 14006 32628 14758
rect 32588 14000 32640 14006
rect 32588 13942 32640 13948
rect 32692 13530 32720 14962
rect 32772 14952 32824 14958
rect 32772 14894 32824 14900
rect 32680 13524 32732 13530
rect 32680 13466 32732 13472
rect 32496 13388 32548 13394
rect 32496 13330 32548 13336
rect 32312 12912 32364 12918
rect 32312 12854 32364 12860
rect 32508 12850 32536 13330
rect 32496 12844 32548 12850
rect 32496 12786 32548 12792
rect 32784 12434 32812 14894
rect 33428 13326 33456 16050
rect 33612 13530 33640 16050
rect 34532 15434 34560 16390
rect 34716 16182 34744 16458
rect 34704 16176 34756 16182
rect 34704 16118 34756 16124
rect 34808 15910 34836 16526
rect 35084 16522 35112 16662
rect 35360 16658 35388 17478
rect 35532 17264 35584 17270
rect 35532 17206 35584 17212
rect 35544 16794 35572 17206
rect 35820 16998 35848 17546
rect 36004 17202 36032 17614
rect 35992 17196 36044 17202
rect 35992 17138 36044 17144
rect 35808 16992 35860 16998
rect 35808 16934 35860 16940
rect 35532 16788 35584 16794
rect 35532 16730 35584 16736
rect 35348 16652 35400 16658
rect 35348 16594 35400 16600
rect 35072 16516 35124 16522
rect 35072 16458 35124 16464
rect 35360 16250 35388 16594
rect 36648 16590 36676 18022
rect 36740 17814 36768 18142
rect 36728 17808 36780 17814
rect 36728 17750 36780 17756
rect 37016 17746 37044 18226
rect 37004 17740 37056 17746
rect 37004 17682 37056 17688
rect 36912 17672 36964 17678
rect 36912 17614 36964 17620
rect 36728 17536 36780 17542
rect 36728 17478 36780 17484
rect 36740 16794 36768 17478
rect 36820 17196 36872 17202
rect 36820 17138 36872 17144
rect 36832 16794 36860 17138
rect 36924 17134 36952 17614
rect 36912 17128 36964 17134
rect 36912 17070 36964 17076
rect 36728 16788 36780 16794
rect 36728 16730 36780 16736
rect 36820 16788 36872 16794
rect 36820 16730 36872 16736
rect 35716 16584 35768 16590
rect 35716 16526 35768 16532
rect 36636 16584 36688 16590
rect 36636 16526 36688 16532
rect 35728 16454 35756 16526
rect 35716 16448 35768 16454
rect 35716 16390 35768 16396
rect 35348 16244 35400 16250
rect 35348 16186 35400 16192
rect 34796 15904 34848 15910
rect 34796 15846 34848 15852
rect 35716 15904 35768 15910
rect 35716 15846 35768 15852
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 35728 15570 35756 15846
rect 35716 15564 35768 15570
rect 35716 15506 35768 15512
rect 37096 15496 37148 15502
rect 37096 15438 37148 15444
rect 34520 15428 34572 15434
rect 34520 15370 34572 15376
rect 35716 15428 35768 15434
rect 35716 15370 35768 15376
rect 35440 15360 35492 15366
rect 35440 15302 35492 15308
rect 35452 15094 35480 15302
rect 35728 15162 35756 15370
rect 35716 15156 35768 15162
rect 35716 15098 35768 15104
rect 35440 15088 35492 15094
rect 35440 15030 35492 15036
rect 33692 14884 33744 14890
rect 33692 14826 33744 14832
rect 33704 14482 33732 14826
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 33692 14476 33744 14482
rect 33692 14418 33744 14424
rect 33784 13728 33836 13734
rect 33784 13670 33836 13676
rect 33600 13524 33652 13530
rect 33600 13466 33652 13472
rect 33416 13320 33468 13326
rect 33416 13262 33468 13268
rect 33048 12912 33100 12918
rect 33048 12854 33100 12860
rect 33060 12434 33088 12854
rect 32692 12406 32812 12434
rect 32876 12406 33088 12434
rect 32692 12306 32720 12406
rect 32680 12300 32732 12306
rect 32680 12242 32732 12248
rect 32404 11620 32456 11626
rect 32404 11562 32456 11568
rect 32312 11552 32364 11558
rect 32312 11494 32364 11500
rect 32324 11082 32352 11494
rect 32416 11082 32444 11562
rect 32588 11552 32640 11558
rect 32588 11494 32640 11500
rect 32312 11076 32364 11082
rect 32312 11018 32364 11024
rect 32404 11076 32456 11082
rect 32404 11018 32456 11024
rect 32600 10266 32628 11494
rect 32588 10260 32640 10266
rect 32588 10202 32640 10208
rect 32404 9920 32456 9926
rect 32404 9862 32456 9868
rect 32416 9586 32444 9862
rect 32404 9580 32456 9586
rect 32404 9522 32456 9528
rect 32220 8424 32272 8430
rect 32220 8366 32272 8372
rect 32312 3528 32364 3534
rect 32312 3470 32364 3476
rect 32324 3058 32352 3470
rect 32496 3392 32548 3398
rect 32496 3334 32548 3340
rect 32508 3126 32536 3334
rect 32496 3120 32548 3126
rect 32496 3062 32548 3068
rect 32312 3052 32364 3058
rect 32312 2994 32364 3000
rect 32220 2984 32272 2990
rect 32220 2926 32272 2932
rect 28356 2848 28408 2854
rect 28356 2790 28408 2796
rect 29000 2372 29052 2378
rect 29000 2314 29052 2320
rect 29012 800 29040 2314
rect 32232 800 32260 2926
rect 32692 2774 32720 12242
rect 32876 11150 32904 12406
rect 33612 11830 33640 13466
rect 33796 13326 33824 13670
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 37108 13326 37136 15438
rect 37200 14346 37228 18294
rect 37556 18284 37608 18290
rect 37556 18226 37608 18232
rect 37924 18284 37976 18290
rect 37924 18226 37976 18232
rect 37568 18170 37596 18226
rect 37568 18142 37688 18170
rect 37280 18080 37332 18086
rect 37280 18022 37332 18028
rect 37292 16658 37320 18022
rect 37372 17672 37424 17678
rect 37372 17614 37424 17620
rect 37464 17672 37516 17678
rect 37464 17614 37516 17620
rect 37384 17270 37412 17614
rect 37372 17264 37424 17270
rect 37372 17206 37424 17212
rect 37280 16652 37332 16658
rect 37280 16594 37332 16600
rect 37384 16590 37412 17206
rect 37476 17134 37504 17614
rect 37464 17128 37516 17134
rect 37464 17070 37516 17076
rect 37476 16658 37504 17070
rect 37660 16998 37688 18142
rect 37648 16992 37700 16998
rect 37648 16934 37700 16940
rect 37464 16652 37516 16658
rect 37464 16594 37516 16600
rect 37372 16584 37424 16590
rect 37372 16526 37424 16532
rect 37372 15360 37424 15366
rect 37372 15302 37424 15308
rect 37384 15094 37412 15302
rect 37372 15088 37424 15094
rect 37372 15030 37424 15036
rect 37476 15026 37504 16594
rect 37464 15020 37516 15026
rect 37464 14962 37516 14968
rect 37936 14550 37964 18226
rect 38304 16726 38332 18906
rect 38476 18760 38528 18766
rect 38476 18702 38528 18708
rect 38488 18426 38516 18702
rect 38660 18624 38712 18630
rect 38660 18566 38712 18572
rect 38476 18420 38528 18426
rect 38476 18362 38528 18368
rect 38672 17678 38700 18566
rect 38764 18290 38792 20810
rect 38948 18290 38976 21286
rect 39028 19780 39080 19786
rect 39028 19722 39080 19728
rect 39040 18970 39068 19722
rect 39488 19304 39540 19310
rect 39488 19246 39540 19252
rect 39028 18964 39080 18970
rect 39028 18906 39080 18912
rect 39120 18760 39172 18766
rect 39120 18702 39172 18708
rect 38752 18284 38804 18290
rect 38752 18226 38804 18232
rect 38936 18284 38988 18290
rect 38936 18226 38988 18232
rect 38660 17672 38712 17678
rect 38660 17614 38712 17620
rect 38292 16720 38344 16726
rect 38292 16662 38344 16668
rect 38948 15502 38976 18226
rect 39132 17882 39160 18702
rect 39120 17876 39172 17882
rect 39120 17818 39172 17824
rect 39132 17338 39160 17818
rect 39120 17332 39172 17338
rect 39120 17274 39172 17280
rect 39500 17202 39528 19246
rect 39488 17196 39540 17202
rect 39488 17138 39540 17144
rect 39500 16590 39528 17138
rect 39488 16584 39540 16590
rect 39488 16526 39540 16532
rect 39500 16182 39528 16526
rect 39488 16176 39540 16182
rect 39488 16118 39540 16124
rect 39304 16108 39356 16114
rect 39304 16050 39356 16056
rect 39316 15706 39344 16050
rect 39304 15700 39356 15706
rect 39304 15642 39356 15648
rect 38936 15496 38988 15502
rect 38936 15438 38988 15444
rect 38936 15360 38988 15366
rect 38936 15302 38988 15308
rect 38200 14816 38252 14822
rect 38200 14758 38252 14764
rect 37924 14544 37976 14550
rect 37924 14486 37976 14492
rect 38212 14414 38240 14758
rect 38948 14618 38976 15302
rect 38936 14612 38988 14618
rect 38936 14554 38988 14560
rect 38948 14414 38976 14554
rect 38200 14408 38252 14414
rect 38200 14350 38252 14356
rect 38752 14408 38804 14414
rect 38752 14350 38804 14356
rect 38936 14408 38988 14414
rect 38936 14350 38988 14356
rect 37188 14340 37240 14346
rect 37188 14282 37240 14288
rect 38016 14068 38068 14074
rect 38016 14010 38068 14016
rect 37556 13932 37608 13938
rect 37556 13874 37608 13880
rect 37568 13530 37596 13874
rect 37556 13524 37608 13530
rect 37556 13466 37608 13472
rect 38028 13326 38056 14010
rect 38212 13326 38240 14350
rect 33784 13320 33836 13326
rect 33784 13262 33836 13268
rect 36820 13320 36872 13326
rect 36820 13262 36872 13268
rect 37096 13320 37148 13326
rect 37096 13262 37148 13268
rect 38016 13320 38068 13326
rect 38016 13262 38068 13268
rect 38200 13320 38252 13326
rect 38200 13262 38252 13268
rect 36728 13252 36780 13258
rect 36728 13194 36780 13200
rect 33784 13184 33836 13190
rect 33784 13126 33836 13132
rect 33796 12238 33824 13126
rect 34152 12844 34204 12850
rect 34152 12786 34204 12792
rect 36360 12844 36412 12850
rect 36360 12786 36412 12792
rect 34164 12442 34192 12786
rect 34520 12640 34572 12646
rect 34520 12582 34572 12588
rect 34152 12436 34204 12442
rect 34152 12378 34204 12384
rect 33784 12232 33836 12238
rect 33784 12174 33836 12180
rect 34532 12170 34560 12582
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 36372 12306 36400 12786
rect 36740 12782 36768 13194
rect 36452 12776 36504 12782
rect 36452 12718 36504 12724
rect 36728 12776 36780 12782
rect 36728 12718 36780 12724
rect 36464 12374 36492 12718
rect 36832 12646 36860 13262
rect 36820 12640 36872 12646
rect 36820 12582 36872 12588
rect 36832 12434 36860 12582
rect 36740 12406 36860 12434
rect 36452 12368 36504 12374
rect 36452 12310 36504 12316
rect 36360 12300 36412 12306
rect 36360 12242 36412 12248
rect 35716 12232 35768 12238
rect 35716 12174 35768 12180
rect 33968 12164 34020 12170
rect 33968 12106 34020 12112
rect 34520 12164 34572 12170
rect 34520 12106 34572 12112
rect 33980 11898 34008 12106
rect 33968 11892 34020 11898
rect 33968 11834 34020 11840
rect 33600 11824 33652 11830
rect 33600 11766 33652 11772
rect 33784 11756 33836 11762
rect 33784 11698 33836 11704
rect 32864 11144 32916 11150
rect 32864 11086 32916 11092
rect 32772 11008 32824 11014
rect 32772 10950 32824 10956
rect 32784 10674 32812 10950
rect 32772 10668 32824 10674
rect 32772 10610 32824 10616
rect 32784 9722 32812 10610
rect 32876 10198 32904 11086
rect 33140 11008 33192 11014
rect 33140 10950 33192 10956
rect 33152 10674 33180 10950
rect 33140 10668 33192 10674
rect 33140 10610 33192 10616
rect 32864 10192 32916 10198
rect 32864 10134 32916 10140
rect 33152 10062 33180 10610
rect 33796 10266 33824 11698
rect 34532 11218 34560 12106
rect 35440 12096 35492 12102
rect 35440 12038 35492 12044
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 35452 11218 35480 12038
rect 34520 11212 34572 11218
rect 34520 11154 34572 11160
rect 35440 11212 35492 11218
rect 35440 11154 35492 11160
rect 34060 11008 34112 11014
rect 34060 10950 34112 10956
rect 35532 11008 35584 11014
rect 35532 10950 35584 10956
rect 34072 10742 34100 10950
rect 35544 10742 35572 10950
rect 34060 10736 34112 10742
rect 34060 10678 34112 10684
rect 35532 10736 35584 10742
rect 35532 10678 35584 10684
rect 33784 10260 33836 10266
rect 33784 10202 33836 10208
rect 34072 10198 34100 10678
rect 35728 10674 35756 12174
rect 36372 11830 36400 12242
rect 36360 11824 36412 11830
rect 36360 11766 36412 11772
rect 35900 11756 35952 11762
rect 35900 11698 35952 11704
rect 35808 11280 35860 11286
rect 35808 11222 35860 11228
rect 35820 10810 35848 11222
rect 35912 11150 35940 11698
rect 36372 11354 36400 11766
rect 36464 11558 36492 12310
rect 36740 11694 36768 12406
rect 37108 12170 37136 13262
rect 37280 13252 37332 13258
rect 37280 13194 37332 13200
rect 37292 12306 37320 13194
rect 37464 13184 37516 13190
rect 37464 13126 37516 13132
rect 37476 12850 37504 13126
rect 37464 12844 37516 12850
rect 37464 12786 37516 12792
rect 37648 12844 37700 12850
rect 37648 12786 37700 12792
rect 37660 12442 37688 12786
rect 37648 12436 37700 12442
rect 37648 12378 37700 12384
rect 37280 12300 37332 12306
rect 37280 12242 37332 12248
rect 37096 12164 37148 12170
rect 37096 12106 37148 12112
rect 37292 11898 37320 12242
rect 38764 12238 38792 14350
rect 38752 12232 38804 12238
rect 38752 12174 38804 12180
rect 37280 11892 37332 11898
rect 37280 11834 37332 11840
rect 38016 11756 38068 11762
rect 38016 11698 38068 11704
rect 38384 11756 38436 11762
rect 38384 11698 38436 11704
rect 36728 11688 36780 11694
rect 36728 11630 36780 11636
rect 36452 11552 36504 11558
rect 36452 11494 36504 11500
rect 36360 11348 36412 11354
rect 36360 11290 36412 11296
rect 35900 11144 35952 11150
rect 35900 11086 35952 11092
rect 35808 10804 35860 10810
rect 35912 10792 35940 11086
rect 35912 10764 36032 10792
rect 35808 10746 35860 10752
rect 35624 10668 35676 10674
rect 35624 10610 35676 10616
rect 35716 10668 35768 10674
rect 35716 10610 35768 10616
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 35636 10266 35664 10610
rect 35624 10260 35676 10266
rect 35624 10202 35676 10208
rect 34060 10192 34112 10198
rect 34060 10134 34112 10140
rect 33140 10056 33192 10062
rect 33140 9998 33192 10004
rect 32772 9716 32824 9722
rect 32772 9658 32824 9664
rect 35636 9450 35664 10202
rect 35728 9722 35756 10610
rect 35900 10464 35952 10470
rect 35900 10406 35952 10412
rect 35912 10062 35940 10406
rect 35900 10056 35952 10062
rect 35900 9998 35952 10004
rect 35716 9716 35768 9722
rect 35716 9658 35768 9664
rect 36004 9518 36032 10764
rect 36740 10606 36768 11630
rect 37832 11552 37884 11558
rect 37832 11494 37884 11500
rect 37844 10742 37872 11494
rect 38028 11150 38056 11698
rect 38292 11552 38344 11558
rect 38292 11494 38344 11500
rect 38108 11212 38160 11218
rect 38108 11154 38160 11160
rect 37924 11144 37976 11150
rect 37924 11086 37976 11092
rect 38016 11144 38068 11150
rect 38016 11086 38068 11092
rect 37936 10996 37964 11086
rect 38120 10996 38148 11154
rect 37936 10968 38148 10996
rect 37832 10736 37884 10742
rect 37832 10678 37884 10684
rect 36728 10600 36780 10606
rect 36728 10542 36780 10548
rect 38200 10532 38252 10538
rect 38200 10474 38252 10480
rect 36912 10464 36964 10470
rect 36912 10406 36964 10412
rect 36924 10130 36952 10406
rect 36912 10124 36964 10130
rect 36912 10066 36964 10072
rect 38212 10062 38240 10474
rect 38304 10470 38332 11494
rect 38396 10742 38424 11698
rect 38568 11552 38620 11558
rect 38568 11494 38620 11500
rect 38476 11144 38528 11150
rect 38476 11086 38528 11092
rect 38384 10736 38436 10742
rect 38384 10678 38436 10684
rect 38488 10606 38516 11086
rect 38580 10810 38608 11494
rect 38660 11008 38712 11014
rect 38660 10950 38712 10956
rect 38672 10810 38700 10950
rect 38568 10804 38620 10810
rect 38568 10746 38620 10752
rect 38660 10804 38712 10810
rect 38660 10746 38712 10752
rect 38476 10600 38528 10606
rect 38476 10542 38528 10548
rect 38292 10464 38344 10470
rect 38292 10406 38344 10412
rect 38304 10266 38332 10406
rect 38292 10260 38344 10266
rect 38292 10202 38344 10208
rect 38200 10056 38252 10062
rect 38200 9998 38252 10004
rect 38016 9920 38068 9926
rect 38016 9862 38068 9868
rect 38028 9586 38056 9862
rect 38016 9580 38068 9586
rect 38016 9522 38068 9528
rect 35992 9512 36044 9518
rect 35992 9454 36044 9460
rect 38488 9450 38516 10542
rect 38764 10062 38792 12174
rect 38948 11694 38976 14350
rect 38936 11688 38988 11694
rect 38936 11630 38988 11636
rect 38948 10674 38976 11630
rect 39120 11348 39172 11354
rect 39120 11290 39172 11296
rect 39132 11150 39160 11290
rect 39120 11144 39172 11150
rect 39120 11086 39172 11092
rect 38936 10668 38988 10674
rect 38936 10610 38988 10616
rect 39212 10600 39264 10606
rect 39212 10542 39264 10548
rect 38568 10056 38620 10062
rect 38568 9998 38620 10004
rect 38752 10056 38804 10062
rect 38752 9998 38804 10004
rect 38580 9722 38608 9998
rect 38568 9716 38620 9722
rect 38568 9658 38620 9664
rect 35624 9444 35676 9450
rect 35624 9386 35676 9392
rect 38476 9444 38528 9450
rect 38476 9386 38528 9392
rect 38764 9382 38792 9998
rect 39224 9994 39252 10542
rect 39212 9988 39264 9994
rect 39212 9930 39264 9936
rect 39224 9382 39252 9930
rect 39396 9920 39448 9926
rect 39396 9862 39448 9868
rect 39408 9586 39436 9862
rect 39396 9580 39448 9586
rect 39396 9522 39448 9528
rect 39488 9580 39540 9586
rect 39488 9522 39540 9528
rect 38752 9376 38804 9382
rect 38752 9318 38804 9324
rect 39212 9376 39264 9382
rect 39212 9318 39264 9324
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 38764 9042 38792 9318
rect 38752 9036 38804 9042
rect 38752 8978 38804 8984
rect 39224 8974 39252 9318
rect 39500 9178 39528 9522
rect 39488 9172 39540 9178
rect 39488 9114 39540 9120
rect 39212 8968 39264 8974
rect 39212 8910 39264 8916
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 39212 6112 39264 6118
rect 39212 6054 39264 6060
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 39028 5704 39080 5710
rect 39028 5646 39080 5652
rect 39040 5234 39068 5646
rect 39224 5302 39252 6054
rect 39212 5296 39264 5302
rect 39212 5238 39264 5244
rect 39028 5228 39080 5234
rect 39028 5170 39080 5176
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 39304 3664 39356 3670
rect 39304 3606 39356 3612
rect 32692 2746 32904 2774
rect 32876 2310 32904 2746
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 38660 2440 38712 2446
rect 38660 2382 38712 2388
rect 32864 2304 32916 2310
rect 32864 2246 32916 2252
rect 38672 800 38700 2382
rect 39316 800 39344 3606
rect 39592 2582 39620 22066
rect 39764 22024 39816 22030
rect 39764 21966 39816 21972
rect 39776 21552 39804 21966
rect 39856 21616 39908 21622
rect 39856 21558 39908 21564
rect 39764 21546 39816 21552
rect 39764 21488 39816 21494
rect 39868 20398 39896 21558
rect 39856 20392 39908 20398
rect 39856 20334 39908 20340
rect 39960 19990 39988 23598
rect 40040 23180 40092 23186
rect 40040 23122 40092 23128
rect 40052 22778 40080 23122
rect 40604 23118 40632 25996
rect 40684 25978 40736 25984
rect 40684 23656 40736 23662
rect 40684 23598 40736 23604
rect 40696 23322 40724 23598
rect 40684 23316 40736 23322
rect 40684 23258 40736 23264
rect 40316 23112 40368 23118
rect 40316 23054 40368 23060
rect 40592 23112 40644 23118
rect 40592 23054 40644 23060
rect 40040 22772 40092 22778
rect 40040 22714 40092 22720
rect 40052 22642 40080 22714
rect 40040 22636 40092 22642
rect 40040 22578 40092 22584
rect 40224 22500 40276 22506
rect 40224 22442 40276 22448
rect 40040 22432 40092 22438
rect 40040 22374 40092 22380
rect 40052 21962 40080 22374
rect 40132 22228 40184 22234
rect 40132 22170 40184 22176
rect 40144 22098 40172 22170
rect 40132 22092 40184 22098
rect 40132 22034 40184 22040
rect 40040 21956 40092 21962
rect 40040 21898 40092 21904
rect 40040 20936 40092 20942
rect 40040 20878 40092 20884
rect 40052 20534 40080 20878
rect 40040 20528 40092 20534
rect 40040 20470 40092 20476
rect 39948 19984 40000 19990
rect 39948 19926 40000 19932
rect 39960 19378 39988 19926
rect 40144 19514 40172 22034
rect 40236 21962 40264 22442
rect 40328 22094 40356 23054
rect 40604 22642 40632 23054
rect 40592 22636 40644 22642
rect 40592 22578 40644 22584
rect 40500 22228 40552 22234
rect 40500 22170 40552 22176
rect 40328 22066 40448 22094
rect 40420 21978 40448 22066
rect 40512 22080 40540 22170
rect 40512 22052 40632 22080
rect 40224 21956 40276 21962
rect 40420 21950 40540 21978
rect 40224 21898 40276 21904
rect 40316 21344 40368 21350
rect 40316 21286 40368 21292
rect 40328 20942 40356 21286
rect 40316 20936 40368 20942
rect 40316 20878 40368 20884
rect 40512 20534 40540 21950
rect 40604 21672 40632 22052
rect 40604 21644 40724 21672
rect 40592 21548 40644 21554
rect 40592 21490 40644 21496
rect 40604 21418 40632 21490
rect 40592 21412 40644 21418
rect 40592 21354 40644 21360
rect 40408 20528 40460 20534
rect 40408 20470 40460 20476
rect 40500 20528 40552 20534
rect 40500 20470 40552 20476
rect 40316 20460 40368 20466
rect 40316 20402 40368 20408
rect 40224 20052 40276 20058
rect 40224 19994 40276 20000
rect 40132 19508 40184 19514
rect 40132 19450 40184 19456
rect 39948 19372 40000 19378
rect 39948 19314 40000 19320
rect 39672 18148 39724 18154
rect 39672 18090 39724 18096
rect 39684 9178 39712 18090
rect 39960 17134 39988 19314
rect 40144 18766 40172 19450
rect 40132 18760 40184 18766
rect 40132 18702 40184 18708
rect 39948 17128 40000 17134
rect 39948 17070 40000 17076
rect 39764 16040 39816 16046
rect 39764 15982 39816 15988
rect 39776 14006 39804 15982
rect 40132 15904 40184 15910
rect 40236 15892 40264 19994
rect 40328 19310 40356 20402
rect 40420 19922 40448 20470
rect 40604 20466 40632 21354
rect 40592 20460 40644 20466
rect 40592 20402 40644 20408
rect 40408 19916 40460 19922
rect 40408 19858 40460 19864
rect 40316 19304 40368 19310
rect 40316 19246 40368 19252
rect 40420 18222 40448 19858
rect 40604 18358 40632 20402
rect 40696 20058 40724 21644
rect 40788 21593 40816 31726
rect 41340 30326 41368 45426
rect 41328 30320 41380 30326
rect 41328 30262 41380 30268
rect 42904 24410 42932 47126
rect 45376 47048 45428 47054
rect 45376 46990 45428 46996
rect 45388 46594 45416 46990
rect 45560 46980 45612 46986
rect 45560 46922 45612 46928
rect 45388 46566 45508 46594
rect 45376 46504 45428 46510
rect 45376 46446 45428 46452
rect 45388 46170 45416 46446
rect 45376 46164 45428 46170
rect 45376 46106 45428 46112
rect 45480 45490 45508 46566
rect 45572 46170 45600 46922
rect 46400 46918 46428 49200
rect 47214 49056 47270 49065
rect 47214 48991 47270 49000
rect 47228 47122 47256 48991
rect 47216 47116 47268 47122
rect 47216 47058 47268 47064
rect 46388 46912 46440 46918
rect 46388 46854 46440 46860
rect 46940 46912 46992 46918
rect 46940 46854 46992 46860
rect 46664 46368 46716 46374
rect 46570 46336 46626 46345
rect 46664 46310 46716 46316
rect 46570 46271 46626 46280
rect 45560 46164 45612 46170
rect 45560 46106 45612 46112
rect 45836 45960 45888 45966
rect 45836 45902 45888 45908
rect 46480 45960 46532 45966
rect 46480 45902 46532 45908
rect 45848 45554 45876 45902
rect 45928 45554 45980 45558
rect 45848 45552 45980 45554
rect 45848 45526 45928 45552
rect 45468 45484 45520 45490
rect 45468 45426 45520 45432
rect 45848 44878 45876 45526
rect 45928 45494 45980 45500
rect 46492 45490 46520 45902
rect 46584 45830 46612 46271
rect 46676 46034 46704 46310
rect 46664 46028 46716 46034
rect 46664 45970 46716 45976
rect 46572 45824 46624 45830
rect 46572 45766 46624 45772
rect 46480 45484 46532 45490
rect 46480 45426 46532 45432
rect 46480 45280 46532 45286
rect 46480 45222 46532 45228
rect 46492 44946 46520 45222
rect 46480 44940 46532 44946
rect 46480 44882 46532 44888
rect 45836 44872 45888 44878
rect 45836 44814 45888 44820
rect 46480 42016 46532 42022
rect 46480 41958 46532 41964
rect 46492 41682 46520 41958
rect 46480 41676 46532 41682
rect 46480 41618 46532 41624
rect 46020 41608 46072 41614
rect 46020 41550 46072 41556
rect 46032 41206 46060 41550
rect 46020 41200 46072 41206
rect 46020 41142 46072 41148
rect 46952 41070 46980 46854
rect 47032 46504 47084 46510
rect 47032 46446 47084 46452
rect 47044 45558 47072 46446
rect 47032 45552 47084 45558
rect 47032 45494 47084 45500
rect 47400 43308 47452 43314
rect 47400 43250 47452 43256
rect 47216 43104 47268 43110
rect 47216 43046 47268 43052
rect 47228 42770 47256 43046
rect 47216 42764 47268 42770
rect 47216 42706 47268 42712
rect 45928 41064 45980 41070
rect 45928 41006 45980 41012
rect 46940 41064 46992 41070
rect 46940 41006 46992 41012
rect 45940 40730 45968 41006
rect 46480 40928 46532 40934
rect 46480 40870 46532 40876
rect 45928 40724 45980 40730
rect 45928 40666 45980 40672
rect 46492 40594 46520 40870
rect 46480 40588 46532 40594
rect 46480 40530 46532 40536
rect 47124 40452 47176 40458
rect 47124 40394 47176 40400
rect 47032 40384 47084 40390
rect 47032 40326 47084 40332
rect 47044 40050 47072 40326
rect 47136 40050 47164 40394
rect 47032 40044 47084 40050
rect 47032 39986 47084 39992
rect 47124 40044 47176 40050
rect 47124 39986 47176 39992
rect 46480 39840 46532 39846
rect 46480 39782 46532 39788
rect 46492 39506 46520 39782
rect 46480 39500 46532 39506
rect 46480 39442 46532 39448
rect 47308 38956 47360 38962
rect 47308 38898 47360 38904
rect 46662 37496 46718 37505
rect 46662 37431 46718 37440
rect 46480 36576 46532 36582
rect 46480 36518 46532 36524
rect 46492 36242 46520 36518
rect 46480 36236 46532 36242
rect 46480 36178 46532 36184
rect 46480 30048 46532 30054
rect 46480 29990 46532 29996
rect 46492 29714 46520 29990
rect 46480 29708 46532 29714
rect 46480 29650 46532 29656
rect 46480 26784 46532 26790
rect 46480 26726 46532 26732
rect 46492 26450 46520 26726
rect 46480 26444 46532 26450
rect 46480 26386 46532 26392
rect 46480 25696 46532 25702
rect 46480 25638 46532 25644
rect 46492 25362 46520 25638
rect 46480 25356 46532 25362
rect 46480 25298 46532 25304
rect 42892 24404 42944 24410
rect 42892 24346 42944 24352
rect 40868 24064 40920 24070
rect 40868 24006 40920 24012
rect 40880 23730 40908 24006
rect 40868 23724 40920 23730
rect 40868 23666 40920 23672
rect 46296 23724 46348 23730
rect 46296 23666 46348 23672
rect 40880 22778 40908 23666
rect 45928 23112 45980 23118
rect 45928 23054 45980 23060
rect 40868 22772 40920 22778
rect 40868 22714 40920 22720
rect 43076 22636 43128 22642
rect 43076 22578 43128 22584
rect 43812 22636 43864 22642
rect 43812 22578 43864 22584
rect 42892 22568 42944 22574
rect 42892 22510 42944 22516
rect 41512 22432 41564 22438
rect 41512 22374 41564 22380
rect 41524 22098 41552 22374
rect 42904 22166 42932 22510
rect 42892 22160 42944 22166
rect 42892 22102 42944 22108
rect 40960 22092 41012 22098
rect 40960 22034 41012 22040
rect 41512 22092 41564 22098
rect 41512 22034 41564 22040
rect 40868 21956 40920 21962
rect 40868 21898 40920 21904
rect 40880 21690 40908 21898
rect 40868 21684 40920 21690
rect 40868 21626 40920 21632
rect 40774 21584 40830 21593
rect 40830 21528 40908 21536
rect 40774 21519 40776 21528
rect 40828 21508 40908 21528
rect 40776 21490 40828 21496
rect 40788 21459 40816 21490
rect 40880 20482 40908 21508
rect 40972 21418 41000 22034
rect 41052 22024 41104 22030
rect 41052 21966 41104 21972
rect 40960 21412 41012 21418
rect 40960 21354 41012 21360
rect 41064 21146 41092 21966
rect 42800 21480 42852 21486
rect 42800 21422 42852 21428
rect 41052 21140 41104 21146
rect 41052 21082 41104 21088
rect 42708 21004 42760 21010
rect 42708 20946 42760 20952
rect 41880 20596 41932 20602
rect 41880 20538 41932 20544
rect 40880 20454 41000 20482
rect 40868 20392 40920 20398
rect 40868 20334 40920 20340
rect 40684 20052 40736 20058
rect 40684 19994 40736 20000
rect 40880 18902 40908 20334
rect 40868 18896 40920 18902
rect 40868 18838 40920 18844
rect 40776 18760 40828 18766
rect 40776 18702 40828 18708
rect 40592 18352 40644 18358
rect 40592 18294 40644 18300
rect 40684 18284 40736 18290
rect 40684 18226 40736 18232
rect 40408 18216 40460 18222
rect 40408 18158 40460 18164
rect 40420 16658 40448 18158
rect 40696 17882 40724 18226
rect 40684 17876 40736 17882
rect 40684 17818 40736 17824
rect 40788 17610 40816 18702
rect 40776 17604 40828 17610
rect 40776 17546 40828 17552
rect 40408 16652 40460 16658
rect 40408 16594 40460 16600
rect 40776 16652 40828 16658
rect 40776 16594 40828 16600
rect 40184 15864 40264 15892
rect 40132 15846 40184 15852
rect 40040 15428 40092 15434
rect 40040 15370 40092 15376
rect 39764 14000 39816 14006
rect 39764 13942 39816 13948
rect 40052 13394 40080 15370
rect 40236 15094 40264 15864
rect 40788 15706 40816 16594
rect 40776 15700 40828 15706
rect 40776 15642 40828 15648
rect 40788 15570 40816 15642
rect 40776 15564 40828 15570
rect 40776 15506 40828 15512
rect 40500 15496 40552 15502
rect 40500 15438 40552 15444
rect 40224 15088 40276 15094
rect 40224 15030 40276 15036
rect 40512 14822 40540 15438
rect 40500 14816 40552 14822
rect 40500 14758 40552 14764
rect 40776 14340 40828 14346
rect 40776 14282 40828 14288
rect 40788 14074 40816 14282
rect 40776 14068 40828 14074
rect 40776 14010 40828 14016
rect 40132 13932 40184 13938
rect 40132 13874 40184 13880
rect 40224 13932 40276 13938
rect 40224 13874 40276 13880
rect 40040 13388 40092 13394
rect 40040 13330 40092 13336
rect 40144 12986 40172 13874
rect 40132 12980 40184 12986
rect 40132 12922 40184 12928
rect 40236 12850 40264 13874
rect 40408 13524 40460 13530
rect 40408 13466 40460 13472
rect 40316 13184 40368 13190
rect 40316 13126 40368 13132
rect 40328 12918 40356 13126
rect 40316 12912 40368 12918
rect 40316 12854 40368 12860
rect 40420 12850 40448 13466
rect 40788 12986 40816 14010
rect 40868 14000 40920 14006
rect 40868 13942 40920 13948
rect 40880 13394 40908 13942
rect 40868 13388 40920 13394
rect 40868 13330 40920 13336
rect 40776 12980 40828 12986
rect 40776 12922 40828 12928
rect 40224 12844 40276 12850
rect 40224 12786 40276 12792
rect 40408 12844 40460 12850
rect 40408 12786 40460 12792
rect 40420 12646 40448 12786
rect 40788 12782 40816 12922
rect 40776 12776 40828 12782
rect 40776 12718 40828 12724
rect 40408 12640 40460 12646
rect 40408 12582 40460 12588
rect 40420 12434 40448 12582
rect 40420 12406 40632 12434
rect 40316 11212 40368 11218
rect 40316 11154 40368 11160
rect 40132 10804 40184 10810
rect 40132 10746 40184 10752
rect 40144 9586 40172 10746
rect 40328 10674 40356 11154
rect 40316 10668 40368 10674
rect 40316 10610 40368 10616
rect 40408 10464 40460 10470
rect 40408 10406 40460 10412
rect 40224 10056 40276 10062
rect 40224 9998 40276 10004
rect 40236 9654 40264 9998
rect 40316 9988 40368 9994
rect 40316 9930 40368 9936
rect 40224 9648 40276 9654
rect 40224 9590 40276 9596
rect 40132 9580 40184 9586
rect 40132 9522 40184 9528
rect 40328 9518 40356 9930
rect 40420 9586 40448 10406
rect 40604 9926 40632 12406
rect 40868 11212 40920 11218
rect 40868 11154 40920 11160
rect 40880 10674 40908 11154
rect 40868 10668 40920 10674
rect 40868 10610 40920 10616
rect 40880 10266 40908 10610
rect 40868 10260 40920 10266
rect 40868 10202 40920 10208
rect 40592 9920 40644 9926
rect 40592 9862 40644 9868
rect 40604 9586 40632 9862
rect 40684 9716 40736 9722
rect 40684 9658 40736 9664
rect 40696 9586 40724 9658
rect 40408 9580 40460 9586
rect 40408 9522 40460 9528
rect 40592 9580 40644 9586
rect 40592 9522 40644 9528
rect 40684 9580 40736 9586
rect 40684 9522 40736 9528
rect 40316 9512 40368 9518
rect 40316 9454 40368 9460
rect 39672 9172 39724 9178
rect 39672 9114 39724 9120
rect 40040 5160 40092 5166
rect 40040 5102 40092 5108
rect 39948 4480 40000 4486
rect 39948 4422 40000 4428
rect 39960 4146 39988 4422
rect 39948 4140 40000 4146
rect 39948 4082 40000 4088
rect 40052 3670 40080 5102
rect 40132 3936 40184 3942
rect 40132 3878 40184 3884
rect 40776 3936 40828 3942
rect 40776 3878 40828 3884
rect 40040 3664 40092 3670
rect 40040 3606 40092 3612
rect 39948 3528 40000 3534
rect 39948 3470 40000 3476
rect 39960 3058 39988 3470
rect 40144 3126 40172 3878
rect 40788 3602 40816 3878
rect 40776 3596 40828 3602
rect 40776 3538 40828 3544
rect 40972 3466 41000 20454
rect 41892 19718 41920 20538
rect 42720 20534 42748 20946
rect 42812 20942 42840 21422
rect 42904 21146 42932 22102
rect 43088 21690 43116 22578
rect 43628 22432 43680 22438
rect 43628 22374 43680 22380
rect 43076 21684 43128 21690
rect 43076 21626 43128 21632
rect 43640 21554 43668 22374
rect 43824 21690 43852 22578
rect 44364 22432 44416 22438
rect 44364 22374 44416 22380
rect 45468 22432 45520 22438
rect 45468 22374 45520 22380
rect 44088 22160 44140 22166
rect 44088 22102 44140 22108
rect 44100 21894 44128 22102
rect 43996 21888 44048 21894
rect 43996 21830 44048 21836
rect 44088 21888 44140 21894
rect 44088 21830 44140 21836
rect 43812 21684 43864 21690
rect 43812 21626 43864 21632
rect 43076 21548 43128 21554
rect 43076 21490 43128 21496
rect 43352 21548 43404 21554
rect 43352 21490 43404 21496
rect 43628 21548 43680 21554
rect 43628 21490 43680 21496
rect 42892 21140 42944 21146
rect 42892 21082 42944 21088
rect 42800 20936 42852 20942
rect 42800 20878 42852 20884
rect 42984 20936 43036 20942
rect 42984 20878 43036 20884
rect 42708 20528 42760 20534
rect 42708 20470 42760 20476
rect 42156 19848 42208 19854
rect 42156 19790 42208 19796
rect 41880 19712 41932 19718
rect 41880 19654 41932 19660
rect 41892 19378 41920 19654
rect 41880 19372 41932 19378
rect 41880 19314 41932 19320
rect 42168 18970 42196 19790
rect 42156 18964 42208 18970
rect 42156 18906 42208 18912
rect 42616 18420 42668 18426
rect 42616 18362 42668 18368
rect 41696 18352 41748 18358
rect 41696 18294 41748 18300
rect 41708 17678 41736 18294
rect 42628 18290 42656 18362
rect 42064 18284 42116 18290
rect 42064 18226 42116 18232
rect 42616 18284 42668 18290
rect 42616 18226 42668 18232
rect 42076 17678 42104 18226
rect 42720 18222 42748 20470
rect 42800 19372 42852 19378
rect 42800 19314 42852 19320
rect 42812 18766 42840 19314
rect 42800 18760 42852 18766
rect 42800 18702 42852 18708
rect 42892 18760 42944 18766
rect 42892 18702 42944 18708
rect 42708 18216 42760 18222
rect 42708 18158 42760 18164
rect 41052 17672 41104 17678
rect 41052 17614 41104 17620
rect 41696 17672 41748 17678
rect 41696 17614 41748 17620
rect 42064 17672 42116 17678
rect 42064 17614 42116 17620
rect 41064 17338 41092 17614
rect 41604 17536 41656 17542
rect 41604 17478 41656 17484
rect 41052 17332 41104 17338
rect 41052 17274 41104 17280
rect 41616 17202 41644 17478
rect 41604 17196 41656 17202
rect 41604 17138 41656 17144
rect 41788 16652 41840 16658
rect 41788 16594 41840 16600
rect 41604 16244 41656 16250
rect 41604 16186 41656 16192
rect 41616 15502 41644 16186
rect 41800 16114 41828 16594
rect 41880 16176 41932 16182
rect 41880 16118 41932 16124
rect 41788 16108 41840 16114
rect 41788 16050 41840 16056
rect 41696 15904 41748 15910
rect 41696 15846 41748 15852
rect 41604 15496 41656 15502
rect 41604 15438 41656 15444
rect 41420 15360 41472 15366
rect 41420 15302 41472 15308
rect 41432 15162 41460 15302
rect 41420 15156 41472 15162
rect 41420 15098 41472 15104
rect 41616 14770 41644 15438
rect 41708 14890 41736 15846
rect 41800 15570 41828 16050
rect 41892 15570 41920 16118
rect 42076 15978 42104 17614
rect 42800 17536 42852 17542
rect 42800 17478 42852 17484
rect 42708 17060 42760 17066
rect 42708 17002 42760 17008
rect 42064 15972 42116 15978
rect 42064 15914 42116 15920
rect 41972 15904 42024 15910
rect 41972 15846 42024 15852
rect 41788 15564 41840 15570
rect 41788 15506 41840 15512
rect 41880 15564 41932 15570
rect 41880 15506 41932 15512
rect 41984 15502 42012 15846
rect 42720 15706 42748 17002
rect 42812 16590 42840 17478
rect 42904 17202 42932 18702
rect 42996 18290 43024 20878
rect 43088 20874 43116 21490
rect 43076 20868 43128 20874
rect 43076 20810 43128 20816
rect 43364 20806 43392 21490
rect 43444 21412 43496 21418
rect 43444 21354 43496 21360
rect 43456 21146 43484 21354
rect 44008 21146 44036 21830
rect 44376 21554 44404 22374
rect 45480 22030 45508 22374
rect 45940 22098 45968 23054
rect 46112 23044 46164 23050
rect 46112 22986 46164 22992
rect 46124 22778 46152 22986
rect 46112 22772 46164 22778
rect 46112 22714 46164 22720
rect 46308 22642 46336 23666
rect 46388 23520 46440 23526
rect 46388 23462 46440 23468
rect 46296 22636 46348 22642
rect 46296 22578 46348 22584
rect 46400 22098 46428 23462
rect 46570 22536 46626 22545
rect 46570 22471 46626 22480
rect 46584 22166 46612 22471
rect 46572 22160 46624 22166
rect 46572 22102 46624 22108
rect 46676 22098 46704 37431
rect 47320 32774 47348 38898
rect 47412 35698 47440 43250
rect 47492 39976 47544 39982
rect 47492 39918 47544 39924
rect 47400 35692 47452 35698
rect 47400 35634 47452 35640
rect 47308 32768 47360 32774
rect 47308 32710 47360 32716
rect 47412 32586 47440 35634
rect 47136 32558 47440 32586
rect 47136 26234 47164 32558
rect 47308 30252 47360 30258
rect 47308 30194 47360 30200
rect 47216 28960 47268 28966
rect 47216 28902 47268 28908
rect 47228 28626 47256 28902
rect 47216 28620 47268 28626
rect 47216 28562 47268 28568
rect 47216 27872 47268 27878
rect 47216 27814 47268 27820
rect 47228 27538 47256 27814
rect 47216 27532 47268 27538
rect 47216 27474 47268 27480
rect 47044 26206 47164 26234
rect 47044 24818 47072 26206
rect 47124 25220 47176 25226
rect 47124 25162 47176 25168
rect 47136 24818 47164 25162
rect 47032 24812 47084 24818
rect 47032 24754 47084 24760
rect 47124 24812 47176 24818
rect 47124 24754 47176 24760
rect 46848 24676 46900 24682
rect 46848 24618 46900 24624
rect 46860 23905 46888 24618
rect 46940 24608 46992 24614
rect 46940 24550 46992 24556
rect 46846 23896 46902 23905
rect 46846 23831 46902 23840
rect 46952 23798 46980 24550
rect 46940 23792 46992 23798
rect 46940 23734 46992 23740
rect 46848 22636 46900 22642
rect 46848 22578 46900 22584
rect 45928 22092 45980 22098
rect 45928 22034 45980 22040
rect 46388 22092 46440 22098
rect 46388 22034 46440 22040
rect 46664 22092 46716 22098
rect 46664 22034 46716 22040
rect 45468 22024 45520 22030
rect 45468 21966 45520 21972
rect 45192 21888 45244 21894
rect 45192 21830 45244 21836
rect 45204 21622 45232 21830
rect 45192 21616 45244 21622
rect 45192 21558 45244 21564
rect 44364 21548 44416 21554
rect 44364 21490 44416 21496
rect 43444 21140 43496 21146
rect 43444 21082 43496 21088
rect 43996 21140 44048 21146
rect 43996 21082 44048 21088
rect 43352 20800 43404 20806
rect 43352 20742 43404 20748
rect 44272 20800 44324 20806
rect 44272 20742 44324 20748
rect 43364 19802 43392 20742
rect 44284 19854 44312 20742
rect 44272 19848 44324 19854
rect 43364 19786 43484 19802
rect 44272 19790 44324 19796
rect 43364 19780 43496 19786
rect 43364 19774 43444 19780
rect 43444 19722 43496 19728
rect 43352 19712 43404 19718
rect 43352 19654 43404 19660
rect 43364 19378 43392 19654
rect 43456 19446 43484 19722
rect 44180 19712 44232 19718
rect 44180 19654 44232 19660
rect 43536 19508 43588 19514
rect 43536 19450 43588 19456
rect 43812 19508 43864 19514
rect 43812 19450 43864 19456
rect 43444 19440 43496 19446
rect 43444 19382 43496 19388
rect 43352 19372 43404 19378
rect 43352 19314 43404 19320
rect 43076 19168 43128 19174
rect 43076 19110 43128 19116
rect 43088 18766 43116 19110
rect 43076 18760 43128 18766
rect 43076 18702 43128 18708
rect 43548 18698 43576 19450
rect 43352 18692 43404 18698
rect 43352 18634 43404 18640
rect 43536 18692 43588 18698
rect 43536 18634 43588 18640
rect 42984 18284 43036 18290
rect 42984 18226 43036 18232
rect 43260 18080 43312 18086
rect 43260 18022 43312 18028
rect 43272 17542 43300 18022
rect 43260 17536 43312 17542
rect 43260 17478 43312 17484
rect 42892 17196 42944 17202
rect 42892 17138 42944 17144
rect 42800 16584 42852 16590
rect 42800 16526 42852 16532
rect 42904 16402 42932 17138
rect 43272 17134 43300 17478
rect 43260 17128 43312 17134
rect 43260 17070 43312 17076
rect 42812 16374 42932 16402
rect 42708 15700 42760 15706
rect 42708 15642 42760 15648
rect 42720 15570 42748 15642
rect 42708 15564 42760 15570
rect 42708 15506 42760 15512
rect 41972 15496 42024 15502
rect 41972 15438 42024 15444
rect 41696 14884 41748 14890
rect 41696 14826 41748 14832
rect 41616 14742 41736 14770
rect 41512 14000 41564 14006
rect 41512 13942 41564 13948
rect 41524 13326 41552 13942
rect 41604 13932 41656 13938
rect 41604 13874 41656 13880
rect 41616 13326 41644 13874
rect 41512 13320 41564 13326
rect 41512 13262 41564 13268
rect 41604 13320 41656 13326
rect 41604 13262 41656 13268
rect 41708 12986 41736 14742
rect 41984 14618 42012 15438
rect 42812 15094 42840 16374
rect 43076 15428 43128 15434
rect 43076 15370 43128 15376
rect 43088 15162 43116 15370
rect 43076 15156 43128 15162
rect 43076 15098 43128 15104
rect 42800 15088 42852 15094
rect 42800 15030 42852 15036
rect 43364 15042 43392 18634
rect 43824 18426 43852 19450
rect 44192 18834 44220 19654
rect 44284 19446 44312 19790
rect 44272 19440 44324 19446
rect 44272 19382 44324 19388
rect 44272 19168 44324 19174
rect 44272 19110 44324 19116
rect 44180 18828 44232 18834
rect 44180 18770 44232 18776
rect 44284 18766 44312 19110
rect 44272 18760 44324 18766
rect 44272 18702 44324 18708
rect 44180 18692 44232 18698
rect 44180 18634 44232 18640
rect 43812 18420 43864 18426
rect 43812 18362 43864 18368
rect 43996 18352 44048 18358
rect 43996 18294 44048 18300
rect 43444 18080 43496 18086
rect 43444 18022 43496 18028
rect 43456 17746 43484 18022
rect 43444 17740 43496 17746
rect 43444 17682 43496 17688
rect 43456 17338 43484 17682
rect 44008 17610 44036 18294
rect 43996 17604 44048 17610
rect 43996 17546 44048 17552
rect 43444 17332 43496 17338
rect 43444 17274 43496 17280
rect 43628 17196 43680 17202
rect 43628 17138 43680 17144
rect 43640 16794 43668 17138
rect 44192 16998 44220 18634
rect 44376 18290 44404 21490
rect 45480 21010 45508 21966
rect 45940 21690 45968 22034
rect 45928 21684 45980 21690
rect 45928 21626 45980 21632
rect 45468 21004 45520 21010
rect 45468 20946 45520 20952
rect 45940 20942 45968 21626
rect 46664 21344 46716 21350
rect 46664 21286 46716 21292
rect 46676 21010 46704 21286
rect 46664 21004 46716 21010
rect 46664 20946 46716 20952
rect 45928 20936 45980 20942
rect 45928 20878 45980 20884
rect 46860 20466 46888 22578
rect 47044 22522 47072 24754
rect 46952 22494 47072 22522
rect 46572 20460 46624 20466
rect 46572 20402 46624 20408
rect 46848 20460 46900 20466
rect 46848 20402 46900 20408
rect 44456 19916 44508 19922
rect 44456 19858 44508 19864
rect 44468 19378 44496 19858
rect 44548 19848 44600 19854
rect 44548 19790 44600 19796
rect 44456 19372 44508 19378
rect 44456 19314 44508 19320
rect 44468 18902 44496 19314
rect 44456 18896 44508 18902
rect 44456 18838 44508 18844
rect 44468 18426 44496 18838
rect 44456 18420 44508 18426
rect 44456 18362 44508 18368
rect 44364 18284 44416 18290
rect 44364 18226 44416 18232
rect 44376 17270 44404 18226
rect 44364 17264 44416 17270
rect 44364 17206 44416 17212
rect 43812 16992 43864 16998
rect 43812 16934 43864 16940
rect 44180 16992 44232 16998
rect 44180 16934 44232 16940
rect 43628 16788 43680 16794
rect 43628 16730 43680 16736
rect 41972 14612 42024 14618
rect 41972 14554 42024 14560
rect 41984 13938 42012 14554
rect 41972 13932 42024 13938
rect 41972 13874 42024 13880
rect 41788 13864 41840 13870
rect 41788 13806 41840 13812
rect 41800 13326 41828 13806
rect 41788 13320 41840 13326
rect 41788 13262 41840 13268
rect 42248 13320 42300 13326
rect 42248 13262 42300 13268
rect 41696 12980 41748 12986
rect 41696 12922 41748 12928
rect 41144 12844 41196 12850
rect 41144 12786 41196 12792
rect 41236 12844 41288 12850
rect 41236 12786 41288 12792
rect 41156 12238 41184 12786
rect 41248 12306 41276 12786
rect 41328 12708 41380 12714
rect 41328 12650 41380 12656
rect 41236 12300 41288 12306
rect 41236 12242 41288 12248
rect 41144 12232 41196 12238
rect 41144 12174 41196 12180
rect 41156 11898 41184 12174
rect 41340 12102 41368 12650
rect 41800 12442 41828 13262
rect 42260 12918 42288 13262
rect 42248 12912 42300 12918
rect 42248 12854 42300 12860
rect 42812 12730 42840 15030
rect 43364 15026 43484 15042
rect 43364 15020 43496 15026
rect 43364 15014 43444 15020
rect 42892 14408 42944 14414
rect 42892 14350 42944 14356
rect 42904 13938 42932 14350
rect 42892 13932 42944 13938
rect 42892 13874 42944 13880
rect 42904 13326 42932 13874
rect 43364 13530 43392 15014
rect 43444 14962 43496 14968
rect 43720 15020 43772 15026
rect 43720 14962 43772 14968
rect 43732 14482 43760 14962
rect 43720 14476 43772 14482
rect 43720 14418 43772 14424
rect 43732 13938 43760 14418
rect 43720 13932 43772 13938
rect 43720 13874 43772 13880
rect 43628 13864 43680 13870
rect 43680 13812 43760 13818
rect 43628 13806 43760 13812
rect 43536 13796 43588 13802
rect 43640 13790 43760 13806
rect 43536 13738 43588 13744
rect 43352 13524 43404 13530
rect 43352 13466 43404 13472
rect 43548 13326 43576 13738
rect 43628 13728 43680 13734
rect 43628 13670 43680 13676
rect 42892 13320 42944 13326
rect 42892 13262 42944 13268
rect 43536 13320 43588 13326
rect 43536 13262 43588 13268
rect 42904 13002 42932 13262
rect 43168 13184 43220 13190
rect 43168 13126 43220 13132
rect 42904 12974 43024 13002
rect 42996 12850 43024 12974
rect 43180 12850 43208 13126
rect 42892 12844 42944 12850
rect 42892 12786 42944 12792
rect 42984 12844 43036 12850
rect 42984 12786 43036 12792
rect 43168 12844 43220 12850
rect 43168 12786 43220 12792
rect 42720 12702 42840 12730
rect 42720 12646 42748 12702
rect 42708 12640 42760 12646
rect 42708 12582 42760 12588
rect 42800 12640 42852 12646
rect 42800 12582 42852 12588
rect 42812 12442 42840 12582
rect 42904 12442 42932 12786
rect 41788 12436 41840 12442
rect 41788 12378 41840 12384
rect 42800 12436 42852 12442
rect 42800 12378 42852 12384
rect 42892 12436 42944 12442
rect 42892 12378 42944 12384
rect 42904 12102 42932 12378
rect 41328 12096 41380 12102
rect 41328 12038 41380 12044
rect 42892 12096 42944 12102
rect 42892 12038 42944 12044
rect 41144 11892 41196 11898
rect 41144 11834 41196 11840
rect 41340 11286 41368 12038
rect 42800 11688 42852 11694
rect 42800 11630 42852 11636
rect 41328 11280 41380 11286
rect 41328 11222 41380 11228
rect 42812 11014 42840 11630
rect 42996 11150 43024 12786
rect 43260 12708 43312 12714
rect 43260 12650 43312 12656
rect 43272 12238 43300 12650
rect 43260 12232 43312 12238
rect 43260 12174 43312 12180
rect 43076 11756 43128 11762
rect 43076 11698 43128 11704
rect 43088 11354 43116 11698
rect 43272 11694 43300 12174
rect 43640 11762 43668 13670
rect 43732 13326 43760 13790
rect 43720 13320 43772 13326
rect 43720 13262 43772 13268
rect 43720 13184 43772 13190
rect 43720 13126 43772 13132
rect 43732 12170 43760 13126
rect 43824 12481 43852 16934
rect 44560 16726 44588 19790
rect 44640 18624 44692 18630
rect 44640 18566 44692 18572
rect 44652 18358 44680 18566
rect 46480 18420 46532 18426
rect 46480 18362 46532 18368
rect 44640 18352 44692 18358
rect 44640 18294 44692 18300
rect 46492 17746 46520 18362
rect 46584 18290 46612 20402
rect 46664 20256 46716 20262
rect 46664 20198 46716 20204
rect 46676 19922 46704 20198
rect 46664 19916 46716 19922
rect 46664 19858 46716 19864
rect 46572 18284 46624 18290
rect 46572 18226 46624 18232
rect 46480 17740 46532 17746
rect 46480 17682 46532 17688
rect 46388 17128 46440 17134
rect 46388 17070 46440 17076
rect 44548 16720 44600 16726
rect 44548 16662 44600 16668
rect 44088 15360 44140 15366
rect 44088 15302 44140 15308
rect 44100 15026 44128 15302
rect 44088 15020 44140 15026
rect 44088 14962 44140 14968
rect 44180 15020 44232 15026
rect 44180 14962 44232 14968
rect 44192 14482 44220 14962
rect 44364 14952 44416 14958
rect 44364 14894 44416 14900
rect 44456 14952 44508 14958
rect 44456 14894 44508 14900
rect 44272 14816 44324 14822
rect 44272 14758 44324 14764
rect 44284 14618 44312 14758
rect 44376 14618 44404 14894
rect 44272 14612 44324 14618
rect 44272 14554 44324 14560
rect 44364 14612 44416 14618
rect 44364 14554 44416 14560
rect 44284 14498 44312 14554
rect 44180 14476 44232 14482
rect 44284 14470 44404 14498
rect 44180 14418 44232 14424
rect 44192 14074 44220 14418
rect 44272 14408 44324 14414
rect 44272 14350 44324 14356
rect 44180 14068 44232 14074
rect 44180 14010 44232 14016
rect 44192 13326 44220 14010
rect 44180 13320 44232 13326
rect 44180 13262 44232 13268
rect 44180 12844 44232 12850
rect 44284 12832 44312 14350
rect 44232 12804 44312 12832
rect 44180 12786 44232 12792
rect 43810 12472 43866 12481
rect 44192 12442 44220 12786
rect 44376 12782 44404 14470
rect 44468 14414 44496 14894
rect 44456 14408 44508 14414
rect 44456 14350 44508 14356
rect 44364 12776 44416 12782
rect 44364 12718 44416 12724
rect 43810 12407 43866 12416
rect 44180 12436 44232 12442
rect 43720 12164 43772 12170
rect 43720 12106 43772 12112
rect 43628 11756 43680 11762
rect 43628 11698 43680 11704
rect 43260 11688 43312 11694
rect 43260 11630 43312 11636
rect 43076 11348 43128 11354
rect 43076 11290 43128 11296
rect 42984 11144 43036 11150
rect 42984 11086 43036 11092
rect 42800 11008 42852 11014
rect 42800 10950 42852 10956
rect 41052 10804 41104 10810
rect 41052 10746 41104 10752
rect 41604 10804 41656 10810
rect 41604 10746 41656 10752
rect 41064 10538 41092 10746
rect 41052 10532 41104 10538
rect 41052 10474 41104 10480
rect 41144 10464 41196 10470
rect 41144 10406 41196 10412
rect 41156 9654 41184 10406
rect 41616 10198 41644 10746
rect 42616 10532 42668 10538
rect 42616 10474 42668 10480
rect 41604 10192 41656 10198
rect 41604 10134 41656 10140
rect 41616 9654 41644 10134
rect 42628 10130 42656 10474
rect 43536 10464 43588 10470
rect 43536 10406 43588 10412
rect 42616 10124 42668 10130
rect 42616 10066 42668 10072
rect 42064 10056 42116 10062
rect 42064 9998 42116 10004
rect 41144 9648 41196 9654
rect 41144 9590 41196 9596
rect 41604 9648 41656 9654
rect 41604 9590 41656 9596
rect 42076 9518 42104 9998
rect 42628 9586 42656 10066
rect 43548 10062 43576 10406
rect 43824 10062 43852 12407
rect 44180 12378 44232 12384
rect 44456 11756 44508 11762
rect 44456 11698 44508 11704
rect 44180 11552 44232 11558
rect 44180 11494 44232 11500
rect 43904 11212 43956 11218
rect 43904 11154 43956 11160
rect 43916 10130 43944 11154
rect 44192 11082 44220 11494
rect 44468 11354 44496 11698
rect 44456 11348 44508 11354
rect 44456 11290 44508 11296
rect 44456 11144 44508 11150
rect 44456 11086 44508 11092
rect 44180 11076 44232 11082
rect 44180 11018 44232 11024
rect 44192 10674 44220 11018
rect 44180 10668 44232 10674
rect 44180 10610 44232 10616
rect 44088 10600 44140 10606
rect 44088 10542 44140 10548
rect 43904 10124 43956 10130
rect 43904 10066 43956 10072
rect 43536 10056 43588 10062
rect 43536 9998 43588 10004
rect 43812 10056 43864 10062
rect 43812 9998 43864 10004
rect 43260 9920 43312 9926
rect 43260 9862 43312 9868
rect 43272 9654 43300 9862
rect 43824 9722 43852 9998
rect 43916 9722 43944 10066
rect 44100 10062 44128 10542
rect 44192 10130 44220 10610
rect 44468 10606 44496 11086
rect 44560 10674 44588 16662
rect 46400 16046 46428 17070
rect 46480 16992 46532 16998
rect 46480 16934 46532 16940
rect 46492 16658 46520 16934
rect 46480 16652 46532 16658
rect 46480 16594 46532 16600
rect 46388 16040 46440 16046
rect 46388 15982 46440 15988
rect 45468 14068 45520 14074
rect 45468 14010 45520 14016
rect 44640 13864 44692 13870
rect 44640 13806 44692 13812
rect 45100 13864 45152 13870
rect 45100 13806 45152 13812
rect 44652 10742 44680 13806
rect 44916 13456 44968 13462
rect 44916 13398 44968 13404
rect 44732 12640 44784 12646
rect 44732 12582 44784 12588
rect 44744 11830 44772 12582
rect 44732 11824 44784 11830
rect 44732 11766 44784 11772
rect 44744 11626 44772 11766
rect 44928 11762 44956 13398
rect 45112 13394 45140 13806
rect 45100 13388 45152 13394
rect 45100 13330 45152 13336
rect 45112 13274 45140 13330
rect 45480 13326 45508 14010
rect 45744 13932 45796 13938
rect 45744 13874 45796 13880
rect 45756 13530 45784 13874
rect 45744 13524 45796 13530
rect 45744 13466 45796 13472
rect 45468 13320 45520 13326
rect 45008 13252 45060 13258
rect 45112 13246 45232 13274
rect 45468 13262 45520 13268
rect 45560 13320 45612 13326
rect 45560 13262 45612 13268
rect 45008 13194 45060 13200
rect 45020 12986 45048 13194
rect 45008 12980 45060 12986
rect 45008 12922 45060 12928
rect 45008 12096 45060 12102
rect 45008 12038 45060 12044
rect 44916 11756 44968 11762
rect 44916 11698 44968 11704
rect 44732 11620 44784 11626
rect 44732 11562 44784 11568
rect 44916 11008 44968 11014
rect 44916 10950 44968 10956
rect 44928 10810 44956 10950
rect 44916 10804 44968 10810
rect 44916 10746 44968 10752
rect 44640 10736 44692 10742
rect 44640 10678 44692 10684
rect 44928 10674 44956 10746
rect 44548 10668 44600 10674
rect 44548 10610 44600 10616
rect 44916 10668 44968 10674
rect 44916 10610 44968 10616
rect 44456 10600 44508 10606
rect 44456 10542 44508 10548
rect 44824 10600 44876 10606
rect 44824 10542 44876 10548
rect 44836 10470 44864 10542
rect 44824 10464 44876 10470
rect 44824 10406 44876 10412
rect 44180 10124 44232 10130
rect 44180 10066 44232 10072
rect 44088 10056 44140 10062
rect 44088 9998 44140 10004
rect 43812 9716 43864 9722
rect 43812 9658 43864 9664
rect 43904 9716 43956 9722
rect 43904 9658 43956 9664
rect 43260 9648 43312 9654
rect 43260 9590 43312 9596
rect 42616 9580 42668 9586
rect 42616 9522 42668 9528
rect 42064 9512 42116 9518
rect 42064 9454 42116 9460
rect 41328 9444 41380 9450
rect 41328 9386 41380 9392
rect 41340 8974 41368 9386
rect 43916 9042 43944 9658
rect 44100 9586 44128 9998
rect 44836 9926 44864 10406
rect 44928 10062 44956 10610
rect 44916 10056 44968 10062
rect 44916 9998 44968 10004
rect 44824 9920 44876 9926
rect 44824 9862 44876 9868
rect 44088 9580 44140 9586
rect 44088 9522 44140 9528
rect 44100 9110 44128 9522
rect 44836 9382 44864 9862
rect 45020 9450 45048 12038
rect 45100 11552 45152 11558
rect 45100 11494 45152 11500
rect 45112 11150 45140 11494
rect 45100 11144 45152 11150
rect 45100 11086 45152 11092
rect 45204 10674 45232 13246
rect 45572 12481 45600 13262
rect 45558 12472 45614 12481
rect 45558 12407 45614 12416
rect 45572 11150 45600 12407
rect 45652 11212 45704 11218
rect 45652 11154 45704 11160
rect 45560 11144 45612 11150
rect 45560 11086 45612 11092
rect 45376 10736 45428 10742
rect 45376 10678 45428 10684
rect 45192 10668 45244 10674
rect 45192 10610 45244 10616
rect 45388 9994 45416 10678
rect 45664 10266 45692 11154
rect 45744 11008 45796 11014
rect 45744 10950 45796 10956
rect 45756 10742 45784 10950
rect 45744 10736 45796 10742
rect 45744 10678 45796 10684
rect 45652 10260 45704 10266
rect 45652 10202 45704 10208
rect 45376 9988 45428 9994
rect 45376 9930 45428 9936
rect 45008 9444 45060 9450
rect 45008 9386 45060 9392
rect 44824 9376 44876 9382
rect 44824 9318 44876 9324
rect 44088 9104 44140 9110
rect 44088 9046 44140 9052
rect 43904 9036 43956 9042
rect 43904 8978 43956 8984
rect 45388 8974 45416 9930
rect 45664 9654 45692 10202
rect 45652 9648 45704 9654
rect 45652 9590 45704 9596
rect 41328 8968 41380 8974
rect 41328 8910 41380 8916
rect 45376 8968 45428 8974
rect 45376 8910 45428 8916
rect 43076 6112 43128 6118
rect 43076 6054 43128 6060
rect 46480 6112 46532 6118
rect 46480 6054 46532 6060
rect 43088 4146 43116 6054
rect 46020 5704 46072 5710
rect 46020 5646 46072 5652
rect 46032 5166 46060 5646
rect 46020 5160 46072 5166
rect 46020 5102 46072 5108
rect 44272 5024 44324 5030
rect 44272 4966 44324 4972
rect 45376 5024 45428 5030
rect 45376 4966 45428 4972
rect 44284 4690 44312 4966
rect 45388 4690 45416 4966
rect 44272 4684 44324 4690
rect 44272 4626 44324 4632
rect 45376 4684 45428 4690
rect 45376 4626 45428 4632
rect 45652 4684 45704 4690
rect 45652 4626 45704 4632
rect 44640 4616 44692 4622
rect 44640 4558 44692 4564
rect 43260 4480 43312 4486
rect 43260 4422 43312 4428
rect 43272 4214 43300 4422
rect 43260 4208 43312 4214
rect 43260 4150 43312 4156
rect 43076 4140 43128 4146
rect 43076 4082 43128 4088
rect 41604 4072 41656 4078
rect 41604 4014 41656 4020
rect 41420 3936 41472 3942
rect 41420 3878 41472 3884
rect 41236 3664 41288 3670
rect 41236 3606 41288 3612
rect 40960 3460 41012 3466
rect 40960 3402 41012 3408
rect 40132 3120 40184 3126
rect 40132 3062 40184 3068
rect 39948 3052 40000 3058
rect 39948 2994 40000 3000
rect 40592 2984 40644 2990
rect 40592 2926 40644 2932
rect 39580 2576 39632 2582
rect 39580 2518 39632 2524
rect 40604 800 40632 2926
rect 41248 800 41276 3606
rect 41432 3602 41460 3878
rect 41420 3596 41472 3602
rect 41420 3538 41472 3544
rect 41616 2446 41644 4014
rect 42616 3528 42668 3534
rect 42616 3470 42668 3476
rect 42628 3058 42656 3470
rect 42616 3052 42668 3058
rect 42616 2994 42668 3000
rect 42892 2984 42944 2990
rect 42892 2926 42944 2932
rect 41880 2916 41932 2922
rect 41880 2858 41932 2864
rect 41604 2440 41656 2446
rect 41604 2382 41656 2388
rect 41892 800 41920 2858
rect 42904 2650 42932 2926
rect 42892 2644 42944 2650
rect 42892 2586 42944 2592
rect 44652 2514 44680 4558
rect 44916 4072 44968 4078
rect 44916 4014 44968 4020
rect 44928 3738 44956 4014
rect 44916 3732 44968 3738
rect 44916 3674 44968 3680
rect 44916 3528 44968 3534
rect 44916 3470 44968 3476
rect 44928 3058 44956 3470
rect 45100 3392 45152 3398
rect 45100 3334 45152 3340
rect 45112 3126 45140 3334
rect 45100 3120 45152 3126
rect 45100 3062 45152 3068
rect 44916 3052 44968 3058
rect 44916 2994 44968 3000
rect 45664 2922 45692 4626
rect 46112 3936 46164 3942
rect 46112 3878 46164 3884
rect 46124 3602 46152 3878
rect 46112 3596 46164 3602
rect 46112 3538 46164 3544
rect 45744 2984 45796 2990
rect 45744 2926 45796 2932
rect 45100 2916 45152 2922
rect 45100 2858 45152 2864
rect 45652 2916 45704 2922
rect 45652 2858 45704 2864
rect 44640 2508 44692 2514
rect 44640 2450 44692 2456
rect 43812 2372 43864 2378
rect 43812 2314 43864 2320
rect 43824 800 43852 2314
rect 45112 800 45140 2858
rect 45756 800 45784 2926
rect 46492 2514 46520 6054
rect 46584 3466 46612 18226
rect 46756 18148 46808 18154
rect 46756 18090 46808 18096
rect 46664 18080 46716 18086
rect 46664 18022 46716 18028
rect 46676 17746 46704 18022
rect 46664 17740 46716 17746
rect 46664 17682 46716 17688
rect 46768 16522 46796 18090
rect 46848 17128 46900 17134
rect 46846 17096 46848 17105
rect 46900 17096 46902 17105
rect 46846 17031 46902 17040
rect 46756 16516 46808 16522
rect 46756 16458 46808 16464
rect 46952 16114 46980 22494
rect 47032 21548 47084 21554
rect 47032 21490 47084 21496
rect 46940 16108 46992 16114
rect 46940 16050 46992 16056
rect 47044 15026 47072 21490
rect 47320 19378 47348 30194
rect 47504 28082 47532 39918
rect 47492 28076 47544 28082
rect 47492 28018 47544 28024
rect 47400 24880 47452 24886
rect 47400 24822 47452 24828
rect 47308 19372 47360 19378
rect 47308 19314 47360 19320
rect 47124 19168 47176 19174
rect 47124 19110 47176 19116
rect 47136 18834 47164 19110
rect 47124 18828 47176 18834
rect 47124 18770 47176 18776
rect 47124 17264 47176 17270
rect 47124 17206 47176 17212
rect 47136 16250 47164 17206
rect 47124 16244 47176 16250
rect 47124 16186 47176 16192
rect 47124 15428 47176 15434
rect 47124 15370 47176 15376
rect 47136 15162 47164 15370
rect 47124 15156 47176 15162
rect 47124 15098 47176 15104
rect 47032 15020 47084 15026
rect 47032 14962 47084 14968
rect 47044 13938 47072 14962
rect 47032 13932 47084 13938
rect 47032 13874 47084 13880
rect 47044 6322 47072 13874
rect 47124 13728 47176 13734
rect 47124 13670 47176 13676
rect 47136 13394 47164 13670
rect 47124 13388 47176 13394
rect 47124 13330 47176 13336
rect 47320 12850 47348 19314
rect 47308 12844 47360 12850
rect 47308 12786 47360 12792
rect 47124 12640 47176 12646
rect 47124 12582 47176 12588
rect 47136 12306 47164 12582
rect 47124 12300 47176 12306
rect 47124 12242 47176 12248
rect 47032 6316 47084 6322
rect 47032 6258 47084 6264
rect 47216 6112 47268 6118
rect 47216 6054 47268 6060
rect 47228 5778 47256 6054
rect 47216 5772 47268 5778
rect 47216 5714 47268 5720
rect 47216 5160 47268 5166
rect 47216 5102 47268 5108
rect 46940 4480 46992 4486
rect 46940 4422 46992 4428
rect 46952 4078 46980 4422
rect 46940 4072 46992 4078
rect 46940 4014 46992 4020
rect 47032 3596 47084 3602
rect 47032 3538 47084 3544
rect 46572 3460 46624 3466
rect 46572 3402 46624 3408
rect 46480 2508 46532 2514
rect 46480 2450 46532 2456
rect 46848 2508 46900 2514
rect 46848 2450 46900 2456
rect 46860 2145 46888 2450
rect 46846 2136 46902 2145
rect 46846 2071 46902 2080
rect 47044 800 47072 3538
rect 47228 1465 47256 5102
rect 47412 4146 47440 24822
rect 47596 23186 47624 49286
rect 48290 49200 48402 49800
rect 48934 49200 49046 49800
rect 49578 49200 49690 49800
rect 48226 47016 48282 47025
rect 48226 46951 48282 46960
rect 48044 46912 48096 46918
rect 48044 46854 48096 46860
rect 47768 46572 47820 46578
rect 47768 46514 47820 46520
rect 47780 45490 47808 46514
rect 47768 45484 47820 45490
rect 47768 45426 47820 45432
rect 47768 45348 47820 45354
rect 47768 45290 47820 45296
rect 47780 44402 47808 45290
rect 47860 44804 47912 44810
rect 47860 44746 47912 44752
rect 47872 44538 47900 44746
rect 47860 44532 47912 44538
rect 47860 44474 47912 44480
rect 47768 44396 47820 44402
rect 47768 44338 47820 44344
rect 47780 42226 47808 44338
rect 47860 43104 47912 43110
rect 47860 43046 47912 43052
rect 47872 42634 47900 43046
rect 47860 42628 47912 42634
rect 47860 42570 47912 42576
rect 47768 42220 47820 42226
rect 47768 42162 47820 42168
rect 47676 38344 47728 38350
rect 47676 38286 47728 38292
rect 47688 37126 47716 38286
rect 47780 37874 47808 42162
rect 47860 42016 47912 42022
rect 47860 41958 47912 41964
rect 47872 41682 47900 41958
rect 47860 41676 47912 41682
rect 47860 41618 47912 41624
rect 47860 39364 47912 39370
rect 47860 39306 47912 39312
rect 47872 39098 47900 39306
rect 47860 39092 47912 39098
rect 47860 39034 47912 39040
rect 47768 37868 47820 37874
rect 47768 37810 47820 37816
rect 47860 37664 47912 37670
rect 47860 37606 47912 37612
rect 47872 37194 47900 37606
rect 47860 37188 47912 37194
rect 47860 37130 47912 37136
rect 47676 37120 47728 37126
rect 47676 37062 47728 37068
rect 47860 36100 47912 36106
rect 47860 36042 47912 36048
rect 47872 35834 47900 36042
rect 47860 35828 47912 35834
rect 47860 35770 47912 35776
rect 47952 33312 48004 33318
rect 47952 33254 48004 33260
rect 47964 32978 47992 33254
rect 47952 32972 48004 32978
rect 47952 32914 48004 32920
rect 47860 32836 47912 32842
rect 47860 32778 47912 32784
rect 47872 32570 47900 32778
rect 47860 32564 47912 32570
rect 47860 32506 47912 32512
rect 47676 30320 47728 30326
rect 47676 30262 47728 30268
rect 47688 29170 47716 30262
rect 47860 30048 47912 30054
rect 47860 29990 47912 29996
rect 47872 29714 47900 29990
rect 47860 29708 47912 29714
rect 47860 29650 47912 29656
rect 47676 29164 47728 29170
rect 47676 29106 47728 29112
rect 47584 23180 47636 23186
rect 47584 23122 47636 23128
rect 47688 18290 47716 29106
rect 47860 28960 47912 28966
rect 47860 28902 47912 28908
rect 47872 28490 47900 28902
rect 47860 28484 47912 28490
rect 47860 28426 47912 28432
rect 47768 28076 47820 28082
rect 47768 28018 47820 28024
rect 47780 25906 47808 28018
rect 47860 27872 47912 27878
rect 47860 27814 47912 27820
rect 47872 27402 47900 27814
rect 47860 27396 47912 27402
rect 47860 27338 47912 27344
rect 47860 26308 47912 26314
rect 47860 26250 47912 26256
rect 47872 26042 47900 26250
rect 47860 26036 47912 26042
rect 47860 25978 47912 25984
rect 47768 25900 47820 25906
rect 47768 25842 47820 25848
rect 47780 24886 47808 25842
rect 47768 24880 47820 24886
rect 47768 24822 47820 24828
rect 47952 21344 48004 21350
rect 47952 21286 48004 21292
rect 47964 21078 47992 21286
rect 48056 21146 48084 46854
rect 48240 46034 48268 46951
rect 48332 46646 48360 49200
rect 48976 47054 49004 49200
rect 48964 47048 49016 47054
rect 48964 46990 49016 46996
rect 48320 46640 48372 46646
rect 48320 46582 48372 46588
rect 48228 46028 48280 46034
rect 48228 45970 48280 45976
rect 48226 44976 48282 44985
rect 48226 44911 48228 44920
rect 48280 44911 48282 44920
rect 48228 44882 48280 44888
rect 48226 42936 48282 42945
rect 48226 42871 48282 42880
rect 48240 42770 48268 42871
rect 48228 42764 48280 42770
rect 48228 42706 48280 42712
rect 48228 41676 48280 41682
rect 48228 41618 48280 41624
rect 48240 41585 48268 41618
rect 48226 41576 48282 41585
rect 48226 41511 48282 41520
rect 48320 40452 48372 40458
rect 48320 40394 48372 40400
rect 48332 40225 48360 40394
rect 48318 40216 48374 40225
rect 48318 40151 48374 40160
rect 48226 39536 48282 39545
rect 48226 39471 48228 39480
rect 48280 39471 48282 39480
rect 48228 39442 48280 39448
rect 48226 38176 48282 38185
rect 48226 38111 48282 38120
rect 48240 37330 48268 38111
rect 48228 37324 48280 37330
rect 48228 37266 48280 37272
rect 48228 36236 48280 36242
rect 48228 36178 48280 36184
rect 48240 36145 48268 36178
rect 48226 36136 48282 36145
rect 48226 36071 48282 36080
rect 48320 32836 48372 32842
rect 48320 32778 48372 32784
rect 48136 32768 48188 32774
rect 48332 32745 48360 32778
rect 48136 32710 48188 32716
rect 48318 32736 48374 32745
rect 48148 32434 48176 32710
rect 48318 32671 48374 32680
rect 48136 32428 48188 32434
rect 48136 32370 48188 32376
rect 48044 21140 48096 21146
rect 48044 21082 48096 21088
rect 47952 21072 48004 21078
rect 47952 21014 48004 21020
rect 47952 20256 48004 20262
rect 47952 20198 48004 20204
rect 47964 19990 47992 20198
rect 47952 19984 48004 19990
rect 47952 19926 48004 19932
rect 47952 19168 48004 19174
rect 47952 19110 48004 19116
rect 47964 18902 47992 19110
rect 47952 18896 48004 18902
rect 47952 18838 48004 18844
rect 47676 18284 47728 18290
rect 47676 18226 47728 18232
rect 47492 12844 47544 12850
rect 47492 12786 47544 12792
rect 47504 5370 47532 12786
rect 47584 5636 47636 5642
rect 47584 5578 47636 5584
rect 47492 5364 47544 5370
rect 47492 5306 47544 5312
rect 47504 4622 47532 5306
rect 47596 4826 47624 5578
rect 47584 4820 47636 4826
rect 47584 4762 47636 4768
rect 47688 4758 47716 18226
rect 48044 17740 48096 17746
rect 48044 17682 48096 17688
rect 47952 15564 48004 15570
rect 47952 15506 48004 15512
rect 47964 15026 47992 15506
rect 47952 15020 48004 15026
rect 47952 14962 48004 14968
rect 47952 13728 48004 13734
rect 47952 13670 48004 13676
rect 47964 13462 47992 13670
rect 47952 13456 48004 13462
rect 47952 13398 48004 13404
rect 47952 12640 48004 12646
rect 47952 12582 48004 12588
rect 47964 12374 47992 12582
rect 47952 12368 48004 12374
rect 48056 12345 48084 17682
rect 47952 12310 48004 12316
rect 48042 12336 48098 12345
rect 48042 12271 48098 12280
rect 47950 8936 48006 8945
rect 47950 8871 47952 8880
rect 48004 8871 48006 8880
rect 47952 8842 48004 8848
rect 47860 8492 47912 8498
rect 47860 8434 47912 8440
rect 47872 8265 47900 8434
rect 47858 8256 47914 8265
rect 47858 8191 47914 8200
rect 47952 7200 48004 7206
rect 47952 7142 48004 7148
rect 47964 6866 47992 7142
rect 47952 6860 48004 6866
rect 47952 6802 48004 6808
rect 47860 6724 47912 6730
rect 47860 6666 47912 6672
rect 47872 6458 47900 6666
rect 47860 6452 47912 6458
rect 47860 6394 47912 6400
rect 47768 6316 47820 6322
rect 47768 6258 47820 6264
rect 47780 5234 47808 6258
rect 47768 5228 47820 5234
rect 47768 5170 47820 5176
rect 47676 4752 47728 4758
rect 47676 4694 47728 4700
rect 48148 4622 48176 32370
rect 48320 29572 48372 29578
rect 48320 29514 48372 29520
rect 48332 29345 48360 29514
rect 48318 29336 48374 29345
rect 48318 29271 48374 29280
rect 48226 28656 48282 28665
rect 48226 28591 48228 28600
rect 48280 28591 48282 28600
rect 48228 28562 48280 28568
rect 48226 27976 48282 27985
rect 48226 27911 48282 27920
rect 48240 27538 48268 27911
rect 48228 27532 48280 27538
rect 48228 27474 48280 27480
rect 48226 26616 48282 26625
rect 48226 26551 48282 26560
rect 48240 26450 48268 26551
rect 48228 26444 48280 26450
rect 48228 26386 48280 26392
rect 48226 25936 48282 25945
rect 48226 25871 48282 25880
rect 48240 25362 48268 25871
rect 48228 25356 48280 25362
rect 48228 25298 48280 25304
rect 48228 24812 48280 24818
rect 48228 24754 48280 24760
rect 48240 24585 48268 24754
rect 48226 24576 48282 24585
rect 48226 24511 48282 24520
rect 48226 21856 48282 21865
rect 48226 21791 48282 21800
rect 48240 21010 48268 21791
rect 48228 21004 48280 21010
rect 48228 20946 48280 20952
rect 48226 20496 48282 20505
rect 48226 20431 48282 20440
rect 48240 19922 48268 20431
rect 48228 19916 48280 19922
rect 48228 19858 48280 19864
rect 48226 19136 48282 19145
rect 48226 19071 48282 19080
rect 48240 18834 48268 19071
rect 48228 18828 48280 18834
rect 48228 18770 48280 18776
rect 48226 17776 48282 17785
rect 48226 17711 48282 17720
rect 48240 16658 48268 17711
rect 48228 16652 48280 16658
rect 48228 16594 48280 16600
rect 48228 15564 48280 15570
rect 48228 15506 48280 15512
rect 48240 15065 48268 15506
rect 48226 15056 48282 15065
rect 48226 14991 48282 15000
rect 48226 13696 48282 13705
rect 48226 13631 48282 13640
rect 48240 13394 48268 13631
rect 48228 13388 48280 13394
rect 48228 13330 48280 13336
rect 48226 13016 48282 13025
rect 48226 12951 48282 12960
rect 48240 12306 48268 12951
rect 48228 12300 48280 12306
rect 48228 12242 48280 12248
rect 48226 6896 48282 6905
rect 48226 6831 48228 6840
rect 48280 6831 48282 6840
rect 48228 6802 48280 6808
rect 48228 5772 48280 5778
rect 48228 5714 48280 5720
rect 48240 5545 48268 5714
rect 48226 5536 48282 5545
rect 48226 5471 48282 5480
rect 47492 4616 47544 4622
rect 47492 4558 47544 4564
rect 48136 4616 48188 4622
rect 48136 4558 48188 4564
rect 48148 4282 48176 4558
rect 48136 4276 48188 4282
rect 48136 4218 48188 4224
rect 47400 4140 47452 4146
rect 47400 4082 47452 4088
rect 47676 4072 47728 4078
rect 47676 4014 47728 4020
rect 47214 1456 47270 1465
rect 47214 1391 47270 1400
rect 47688 800 47716 4014
rect 47952 4004 48004 4010
rect 47952 3946 48004 3952
rect 47964 2650 47992 3946
rect 48320 3732 48372 3738
rect 48320 3674 48372 3680
rect 48042 3496 48098 3505
rect 48042 3431 48098 3440
rect 48056 3058 48084 3431
rect 48044 3052 48096 3058
rect 48044 2994 48096 3000
rect 47952 2644 48004 2650
rect 47952 2586 48004 2592
rect 2778 776 2834 785
rect 2778 711 2834 720
rect 3210 200 3322 800
rect 4498 200 4610 800
rect 5142 200 5254 800
rect 6430 200 6542 800
rect 7074 200 7186 800
rect 7718 200 7830 800
rect 9006 200 9118 800
rect 9650 200 9762 800
rect 10938 200 11050 800
rect 11582 200 11694 800
rect 12870 200 12982 800
rect 13514 200 13626 800
rect 14158 200 14270 800
rect 15446 200 15558 800
rect 16090 200 16202 800
rect 17378 200 17490 800
rect 18022 200 18134 800
rect 19310 200 19422 800
rect 19954 200 20066 800
rect 20598 200 20710 800
rect 21886 200 21998 800
rect 22530 200 22642 800
rect 23818 200 23930 800
rect 24462 200 24574 800
rect 25750 200 25862 800
rect 26394 200 26506 800
rect 27682 200 27794 800
rect 28326 200 28438 800
rect 28970 200 29082 800
rect 30258 200 30370 800
rect 30902 200 31014 800
rect 32190 200 32302 800
rect 32834 200 32946 800
rect 34122 200 34234 800
rect 34766 200 34878 800
rect 35410 200 35522 800
rect 36698 200 36810 800
rect 37342 200 37454 800
rect 38630 200 38742 800
rect 39274 200 39386 800
rect 40562 200 40674 800
rect 41206 200 41318 800
rect 41850 200 41962 800
rect 43138 200 43250 800
rect 43782 200 43894 800
rect 45070 200 45182 800
rect 45714 200 45826 800
rect 47002 200 47114 800
rect 47646 200 47758 800
rect 48332 105 48360 3674
rect 48964 3188 49016 3194
rect 48964 3130 49016 3136
rect 48976 800 49004 3130
rect 48934 200 49046 800
rect 49578 200 49690 800
rect 48318 96 48374 105
rect 48318 31 48374 40
<< via2 >>
rect 1582 38800 1638 38856
rect 2778 48320 2834 48376
rect 2962 47640 3018 47696
rect 2870 46280 2926 46336
rect 2778 45600 2834 45656
rect 2778 43560 2834 43616
rect 1582 36760 1638 36816
rect 1582 34040 1638 34096
rect 1582 32000 1638 32056
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 2778 41520 2834 41576
rect 2778 32680 2834 32736
rect 2778 25200 2834 25256
rect 2778 21800 2834 21856
rect 2962 20440 3018 20496
rect 2778 18400 2834 18456
rect 2778 17040 2834 17096
rect 3514 40840 3570 40896
rect 2778 15000 2834 15056
rect 2778 14320 2834 14376
rect 2778 11636 2780 11656
rect 2780 11636 2832 11656
rect 2832 11636 2834 11656
rect 2778 11600 2834 11636
rect 2778 9560 2834 9616
rect 2778 7520 2834 7576
rect 3146 10240 3202 10296
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4066 23840 4122 23896
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 2778 6860 2834 6896
rect 2778 6840 2780 6860
rect 2780 6840 2832 6860
rect 2832 6840 2834 6860
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 2962 4800 3018 4856
rect 3514 5480 3570 5536
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 2778 3440 2834 3496
rect 2778 2760 2834 2816
rect 2870 1400 2926 1456
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 10414 21548 10470 21584
rect 10414 21528 10416 21548
rect 10416 21528 10468 21548
rect 10468 21528 10470 21548
rect 19706 46980 19762 47016
rect 19706 46960 19708 46980
rect 19708 46960 19760 46980
rect 19760 46960 19762 46980
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 20074 36896 20130 36952
rect 19430 36760 19486 36816
rect 19890 36624 19946 36680
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 20534 36644 20590 36680
rect 20534 36624 20536 36644
rect 20536 36624 20588 36644
rect 20588 36624 20590 36644
rect 20626 35944 20682 36000
rect 22926 37848 22982 37904
rect 23846 37868 23902 37904
rect 23846 37848 23848 37868
rect 23848 37848 23900 37868
rect 23900 37848 23902 37868
rect 23386 37712 23442 37768
rect 23938 37748 23940 37768
rect 23940 37748 23992 37768
rect 23992 37748 23994 37768
rect 23018 36896 23074 36952
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 22466 31320 22522 31376
rect 23938 37712 23994 37748
rect 24582 36780 24638 36816
rect 24582 36760 24584 36780
rect 24584 36760 24636 36780
rect 24636 36760 24638 36780
rect 22650 24384 22706 24440
rect 23202 24404 23258 24440
rect 23202 24384 23204 24404
rect 23204 24384 23256 24404
rect 23256 24384 23258 24404
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 27158 11756 27214 11792
rect 27158 11736 27160 11756
rect 27160 11736 27212 11756
rect 27212 11736 27214 11756
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 28998 21256 29054 21312
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 28630 11756 28686 11792
rect 28630 11736 28632 11756
rect 28632 11736 28684 11756
rect 28684 11736 28686 11756
rect 32494 21256 32550 21312
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 47214 49000 47270 49056
rect 46570 46280 46626 46336
rect 46662 37440 46718 37496
rect 40774 21548 40830 21584
rect 40774 21528 40776 21548
rect 40776 21528 40828 21548
rect 40828 21528 40830 21548
rect 46570 22480 46626 22536
rect 46846 23840 46902 23896
rect 43810 12416 43866 12472
rect 45558 12416 45614 12472
rect 46846 17076 46848 17096
rect 46848 17076 46900 17096
rect 46900 17076 46902 17096
rect 46846 17040 46902 17076
rect 46846 2080 46902 2136
rect 48226 46960 48282 47016
rect 48226 44940 48282 44976
rect 48226 44920 48228 44940
rect 48228 44920 48280 44940
rect 48280 44920 48282 44940
rect 48226 42880 48282 42936
rect 48226 41520 48282 41576
rect 48318 40160 48374 40216
rect 48226 39500 48282 39536
rect 48226 39480 48228 39500
rect 48228 39480 48280 39500
rect 48280 39480 48282 39500
rect 48226 38120 48282 38176
rect 48226 36080 48282 36136
rect 48318 32680 48374 32736
rect 48042 12280 48098 12336
rect 47950 8900 48006 8936
rect 47950 8880 47952 8900
rect 47952 8880 48004 8900
rect 48004 8880 48006 8900
rect 47858 8200 47914 8256
rect 48318 29280 48374 29336
rect 48226 28620 48282 28656
rect 48226 28600 48228 28620
rect 48228 28600 48280 28620
rect 48280 28600 48282 28620
rect 48226 27920 48282 27976
rect 48226 26560 48282 26616
rect 48226 25880 48282 25936
rect 48226 24520 48282 24576
rect 48226 21800 48282 21856
rect 48226 20440 48282 20496
rect 48226 19080 48282 19136
rect 48226 17720 48282 17776
rect 48226 15000 48282 15056
rect 48226 13640 48282 13696
rect 48226 12960 48282 13016
rect 48226 6860 48282 6896
rect 48226 6840 48228 6860
rect 48228 6840 48280 6860
rect 48280 6840 48282 6860
rect 48226 5480 48282 5536
rect 47214 1400 47270 1456
rect 48042 3440 48098 3496
rect 2778 720 2834 776
rect 48318 40 48374 96
<< metal3 >>
rect 200 49588 800 49828
rect 47209 49058 47275 49061
rect 49200 49058 49800 49148
rect 47209 49056 49800 49058
rect 47209 49000 47214 49056
rect 47270 49000 49800 49056
rect 47209 48998 49800 49000
rect 47209 48995 47275 48998
rect 49200 48908 49800 48998
rect 200 48378 800 48468
rect 2773 48378 2839 48381
rect 200 48376 2839 48378
rect 200 48320 2778 48376
rect 2834 48320 2839 48376
rect 200 48318 2839 48320
rect 200 48228 800 48318
rect 2773 48315 2839 48318
rect 49200 48228 49800 48468
rect 200 47698 800 47788
rect 2957 47698 3023 47701
rect 200 47696 3023 47698
rect 200 47640 2962 47696
rect 3018 47640 3023 47696
rect 200 47638 3023 47640
rect 200 47548 800 47638
rect 2957 47635 3023 47638
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 19701 47018 19767 47021
rect 20110 47018 20116 47020
rect 19701 47016 20116 47018
rect 19701 46960 19706 47016
rect 19762 46960 20116 47016
rect 19701 46958 20116 46960
rect 19701 46955 19767 46958
rect 20110 46956 20116 46958
rect 20180 46956 20186 47020
rect 48221 47018 48287 47021
rect 49200 47018 49800 47108
rect 48221 47016 49800 47018
rect 48221 46960 48226 47016
rect 48282 46960 49800 47016
rect 48221 46958 49800 46960
rect 48221 46955 48287 46958
rect 49200 46868 49800 46958
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 200 46338 800 46428
rect 2865 46338 2931 46341
rect 200 46336 2931 46338
rect 200 46280 2870 46336
rect 2926 46280 2931 46336
rect 200 46278 2931 46280
rect 200 46188 800 46278
rect 2865 46275 2931 46278
rect 46565 46338 46631 46341
rect 49200 46338 49800 46428
rect 46565 46336 49800 46338
rect 46565 46280 46570 46336
rect 46626 46280 49800 46336
rect 46565 46278 49800 46280
rect 46565 46275 46631 46278
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 49200 46188 49800 46278
rect 200 45658 800 45748
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 2773 45658 2839 45661
rect 200 45656 2839 45658
rect 200 45600 2778 45656
rect 2834 45600 2839 45656
rect 200 45598 2839 45600
rect 200 45508 800 45598
rect 2773 45595 2839 45598
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 48221 44978 48287 44981
rect 49200 44978 49800 45068
rect 48221 44976 49800 44978
rect 48221 44920 48226 44976
rect 48282 44920 49800 44976
rect 48221 44918 49800 44920
rect 48221 44915 48287 44918
rect 49200 44828 49800 44918
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 200 44148 800 44388
rect 49200 44148 49800 44388
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 200 43618 800 43708
rect 2773 43618 2839 43621
rect 200 43616 2839 43618
rect 200 43560 2778 43616
rect 2834 43560 2839 43616
rect 200 43558 2839 43560
rect 200 43468 800 43558
rect 2773 43555 2839 43558
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 200 42788 800 43028
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 48221 42938 48287 42941
rect 49200 42938 49800 43028
rect 48221 42936 49800 42938
rect 48221 42880 48226 42936
rect 48282 42880 49800 42936
rect 48221 42878 49800 42880
rect 48221 42875 48287 42878
rect 49200 42788 49800 42878
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 49200 42108 49800 42348
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 200 41578 800 41668
rect 2773 41578 2839 41581
rect 200 41576 2839 41578
rect 200 41520 2778 41576
rect 2834 41520 2839 41576
rect 200 41518 2839 41520
rect 200 41428 800 41518
rect 2773 41515 2839 41518
rect 48221 41578 48287 41581
rect 49200 41578 49800 41668
rect 48221 41576 49800 41578
rect 48221 41520 48226 41576
rect 48282 41520 49800 41576
rect 48221 41518 49800 41520
rect 48221 41515 48287 41518
rect 49200 41428 49800 41518
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 200 40898 800 40988
rect 3509 40898 3575 40901
rect 200 40896 3575 40898
rect 200 40840 3514 40896
rect 3570 40840 3575 40896
rect 200 40838 3575 40840
rect 200 40748 800 40838
rect 3509 40835 3575 40838
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 48313 40218 48379 40221
rect 49200 40218 49800 40308
rect 48313 40216 49800 40218
rect 48313 40160 48318 40216
rect 48374 40160 49800 40216
rect 48313 40158 49800 40160
rect 48313 40155 48379 40158
rect 49200 40068 49800 40158
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 200 39388 800 39628
rect 48221 39538 48287 39541
rect 49200 39538 49800 39628
rect 48221 39536 49800 39538
rect 48221 39480 48226 39536
rect 48282 39480 49800 39536
rect 48221 39478 49800 39480
rect 48221 39475 48287 39478
rect 49200 39388 49800 39478
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 200 38858 800 38948
rect 1577 38858 1643 38861
rect 200 38856 1643 38858
rect 200 38800 1582 38856
rect 1638 38800 1643 38856
rect 200 38798 1643 38800
rect 200 38708 800 38798
rect 1577 38795 1643 38798
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 48221 38178 48287 38181
rect 49200 38178 49800 38268
rect 48221 38176 49800 38178
rect 48221 38120 48226 38176
rect 48282 38120 49800 38176
rect 48221 38118 49800 38120
rect 48221 38115 48287 38118
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 49200 38028 49800 38118
rect 22921 37906 22987 37909
rect 23841 37906 23907 37909
rect 22921 37904 23907 37906
rect 22921 37848 22926 37904
rect 22982 37848 23846 37904
rect 23902 37848 23907 37904
rect 22921 37846 23907 37848
rect 22921 37843 22987 37846
rect 23841 37843 23907 37846
rect 23381 37770 23447 37773
rect 23933 37770 23999 37773
rect 23381 37768 23999 37770
rect 23381 37712 23386 37768
rect 23442 37712 23938 37768
rect 23994 37712 23999 37768
rect 23381 37710 23999 37712
rect 23381 37707 23447 37710
rect 23933 37707 23999 37710
rect 200 37348 800 37588
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 46657 37498 46723 37501
rect 49200 37498 49800 37588
rect 46657 37496 49800 37498
rect 46657 37440 46662 37496
rect 46718 37440 49800 37496
rect 46657 37438 49800 37440
rect 46657 37435 46723 37438
rect 49200 37348 49800 37438
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 20069 36954 20135 36957
rect 23013 36954 23079 36957
rect 20069 36952 23079 36954
rect 200 36818 800 36908
rect 20069 36896 20074 36952
rect 20130 36896 23018 36952
rect 23074 36896 23079 36952
rect 20069 36894 23079 36896
rect 20069 36891 20135 36894
rect 23013 36891 23079 36894
rect 1577 36818 1643 36821
rect 200 36816 1643 36818
rect 200 36760 1582 36816
rect 1638 36760 1643 36816
rect 200 36758 1643 36760
rect 200 36668 800 36758
rect 1577 36755 1643 36758
rect 19425 36818 19491 36821
rect 24577 36818 24643 36821
rect 19425 36816 24643 36818
rect 19425 36760 19430 36816
rect 19486 36760 24582 36816
rect 24638 36760 24643 36816
rect 19425 36758 24643 36760
rect 19425 36755 19491 36758
rect 24577 36755 24643 36758
rect 19885 36682 19951 36685
rect 20529 36682 20595 36685
rect 19885 36680 20595 36682
rect 19885 36624 19890 36680
rect 19946 36624 20534 36680
rect 20590 36624 20595 36680
rect 19885 36622 20595 36624
rect 19885 36619 19951 36622
rect 20529 36619 20595 36622
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 200 35988 800 36228
rect 48221 36138 48287 36141
rect 49200 36138 49800 36228
rect 48221 36136 49800 36138
rect 48221 36080 48226 36136
rect 48282 36080 49800 36136
rect 48221 36078 49800 36080
rect 48221 36075 48287 36078
rect 20621 36004 20687 36005
rect 20621 36000 20668 36004
rect 20732 36002 20738 36004
rect 20621 35944 20626 36000
rect 20621 35940 20668 35944
rect 20732 35942 20778 36002
rect 49200 35988 49800 36078
rect 20732 35940 20738 35942
rect 20621 35939 20687 35940
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 49200 35308 49800 35548
rect 200 34628 800 34868
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 49200 34628 49800 34868
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 200 34098 800 34188
rect 1577 34098 1643 34101
rect 200 34096 1643 34098
rect 200 34040 1582 34096
rect 1638 34040 1643 34096
rect 200 34038 1643 34040
rect 200 33948 800 34038
rect 1577 34035 1643 34038
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 49200 33268 49800 33508
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 200 32738 800 32828
rect 2773 32738 2839 32741
rect 200 32736 2839 32738
rect 200 32680 2778 32736
rect 2834 32680 2839 32736
rect 200 32678 2839 32680
rect 200 32588 800 32678
rect 2773 32675 2839 32678
rect 48313 32738 48379 32741
rect 49200 32738 49800 32828
rect 48313 32736 49800 32738
rect 48313 32680 48318 32736
rect 48374 32680 49800 32736
rect 48313 32678 49800 32680
rect 48313 32675 48379 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 49200 32588 49800 32678
rect 200 32058 800 32148
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 1577 32058 1643 32061
rect 200 32056 1643 32058
rect 200 32000 1582 32056
rect 1638 32000 1643 32056
rect 200 31998 1643 32000
rect 200 31908 800 31998
rect 1577 31995 1643 31998
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 20662 31316 20668 31380
rect 20732 31378 20738 31380
rect 22461 31378 22527 31381
rect 20732 31376 22527 31378
rect 20732 31320 22466 31376
rect 22522 31320 22527 31376
rect 20732 31318 22527 31320
rect 20732 31316 20738 31318
rect 22461 31315 22527 31318
rect 49200 31228 49800 31468
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 200 30548 800 30788
rect 49200 30548 49800 30788
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 200 29868 800 30108
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 200 29188 800 29428
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 48313 29338 48379 29341
rect 49200 29338 49800 29428
rect 48313 29336 49800 29338
rect 48313 29280 48318 29336
rect 48374 29280 49800 29336
rect 48313 29278 49800 29280
rect 48313 29275 48379 29278
rect 49200 29188 49800 29278
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 48221 28658 48287 28661
rect 49200 28658 49800 28748
rect 48221 28656 49800 28658
rect 48221 28600 48226 28656
rect 48282 28600 49800 28656
rect 48221 28598 49800 28600
rect 48221 28595 48287 28598
rect 49200 28508 49800 28598
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 200 27828 800 28068
rect 48221 27978 48287 27981
rect 49200 27978 49800 28068
rect 48221 27976 49800 27978
rect 48221 27920 48226 27976
rect 48282 27920 49800 27976
rect 48221 27918 49800 27920
rect 48221 27915 48287 27918
rect 49200 27828 49800 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 200 27148 800 27388
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 48221 26618 48287 26621
rect 49200 26618 49800 26708
rect 48221 26616 49800 26618
rect 48221 26560 48226 26616
rect 48282 26560 49800 26616
rect 48221 26558 49800 26560
rect 48221 26555 48287 26558
rect 49200 26468 49800 26558
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 200 25788 800 26028
rect 48221 25938 48287 25941
rect 49200 25938 49800 26028
rect 48221 25936 49800 25938
rect 48221 25880 48226 25936
rect 48282 25880 49800 25936
rect 48221 25878 49800 25880
rect 48221 25875 48287 25878
rect 49200 25788 49800 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 200 25258 800 25348
rect 2773 25258 2839 25261
rect 200 25256 2839 25258
rect 200 25200 2778 25256
rect 2834 25200 2839 25256
rect 200 25198 2839 25200
rect 200 25108 800 25198
rect 2773 25195 2839 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 48221 24578 48287 24581
rect 49200 24578 49800 24668
rect 48221 24576 49800 24578
rect 48221 24520 48226 24576
rect 48282 24520 49800 24576
rect 48221 24518 49800 24520
rect 48221 24515 48287 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 20110 24380 20116 24444
rect 20180 24442 20186 24444
rect 22645 24442 22711 24445
rect 23197 24442 23263 24445
rect 20180 24440 23263 24442
rect 20180 24384 22650 24440
rect 22706 24384 23202 24440
rect 23258 24384 23263 24440
rect 49200 24428 49800 24518
rect 20180 24382 23263 24384
rect 20180 24380 20186 24382
rect 22645 24379 22711 24382
rect 23197 24379 23263 24382
rect 200 23898 800 23988
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 4061 23898 4127 23901
rect 200 23896 4127 23898
rect 200 23840 4066 23896
rect 4122 23840 4127 23896
rect 200 23838 4127 23840
rect 200 23748 800 23838
rect 4061 23835 4127 23838
rect 46841 23898 46907 23901
rect 49200 23898 49800 23988
rect 46841 23896 49800 23898
rect 46841 23840 46846 23896
rect 46902 23840 49800 23896
rect 46841 23838 49800 23840
rect 46841 23835 46907 23838
rect 49200 23748 49800 23838
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 200 23068 800 23308
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 46565 22538 46631 22541
rect 49200 22538 49800 22628
rect 46565 22536 49800 22538
rect 46565 22480 46570 22536
rect 46626 22480 49800 22536
rect 46565 22478 49800 22480
rect 46565 22475 46631 22478
rect 49200 22388 49800 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 200 21858 800 21948
rect 2773 21858 2839 21861
rect 200 21856 2839 21858
rect 200 21800 2778 21856
rect 2834 21800 2839 21856
rect 200 21798 2839 21800
rect 200 21708 800 21798
rect 2773 21795 2839 21798
rect 48221 21858 48287 21861
rect 49200 21858 49800 21948
rect 48221 21856 49800 21858
rect 48221 21800 48226 21856
rect 48282 21800 49800 21856
rect 48221 21798 49800 21800
rect 48221 21795 48287 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 49200 21708 49800 21798
rect 10409 21586 10475 21589
rect 40769 21586 40835 21589
rect 10409 21584 40835 21586
rect 10409 21528 10414 21584
rect 10470 21528 40774 21584
rect 40830 21528 40835 21584
rect 10409 21526 40835 21528
rect 10409 21523 10475 21526
rect 40769 21523 40835 21526
rect 28993 21314 29059 21317
rect 32489 21314 32555 21317
rect 28993 21312 32555 21314
rect 200 21028 800 21268
rect 28993 21256 28998 21312
rect 29054 21256 32494 21312
rect 32550 21256 32555 21312
rect 28993 21254 32555 21256
rect 28993 21251 29059 21254
rect 32489 21251 32555 21254
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 200 20498 800 20588
rect 2957 20498 3023 20501
rect 200 20496 3023 20498
rect 200 20440 2962 20496
rect 3018 20440 3023 20496
rect 200 20438 3023 20440
rect 200 20348 800 20438
rect 2957 20435 3023 20438
rect 48221 20498 48287 20501
rect 49200 20498 49800 20588
rect 48221 20496 49800 20498
rect 48221 20440 48226 20496
rect 48282 20440 49800 20496
rect 48221 20438 49800 20440
rect 48221 20435 48287 20438
rect 49200 20348 49800 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 49200 19668 49800 19908
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 200 18988 800 19228
rect 48221 19138 48287 19141
rect 49200 19138 49800 19228
rect 48221 19136 49800 19138
rect 48221 19080 48226 19136
rect 48282 19080 49800 19136
rect 48221 19078 49800 19080
rect 48221 19075 48287 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 49200 18988 49800 19078
rect 200 18458 800 18548
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 2773 18458 2839 18461
rect 200 18456 2839 18458
rect 200 18400 2778 18456
rect 2834 18400 2839 18456
rect 200 18398 2839 18400
rect 200 18308 800 18398
rect 2773 18395 2839 18398
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 48221 17778 48287 17781
rect 49200 17778 49800 17868
rect 48221 17776 49800 17778
rect 48221 17720 48226 17776
rect 48282 17720 49800 17776
rect 48221 17718 49800 17720
rect 48221 17715 48287 17718
rect 49200 17628 49800 17718
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 200 17098 800 17188
rect 2773 17098 2839 17101
rect 200 17096 2839 17098
rect 200 17040 2778 17096
rect 2834 17040 2839 17096
rect 200 17038 2839 17040
rect 200 16948 800 17038
rect 2773 17035 2839 17038
rect 46841 17098 46907 17101
rect 49200 17098 49800 17188
rect 46841 17096 49800 17098
rect 46841 17040 46846 17096
rect 46902 17040 49800 17096
rect 46841 17038 49800 17040
rect 46841 17035 46907 17038
rect 49200 16948 49800 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 200 16268 800 16508
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 49200 15588 49800 15828
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 200 15058 800 15148
rect 2773 15058 2839 15061
rect 200 15056 2839 15058
rect 200 15000 2778 15056
rect 2834 15000 2839 15056
rect 200 14998 2839 15000
rect 200 14908 800 14998
rect 2773 14995 2839 14998
rect 48221 15058 48287 15061
rect 49200 15058 49800 15148
rect 48221 15056 49800 15058
rect 48221 15000 48226 15056
rect 48282 15000 49800 15056
rect 48221 14998 49800 15000
rect 48221 14995 48287 14998
rect 49200 14908 49800 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 200 14378 800 14468
rect 2773 14378 2839 14381
rect 200 14376 2839 14378
rect 200 14320 2778 14376
rect 2834 14320 2839 14376
rect 200 14318 2839 14320
rect 200 14228 800 14318
rect 2773 14315 2839 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 200 13548 800 13788
rect 48221 13698 48287 13701
rect 49200 13698 49800 13788
rect 48221 13696 49800 13698
rect 48221 13640 48226 13696
rect 48282 13640 49800 13696
rect 48221 13638 49800 13640
rect 48221 13635 48287 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 49200 13548 49800 13638
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 48221 13018 48287 13021
rect 49200 13018 49800 13108
rect 48221 13016 49800 13018
rect 48221 12960 48226 13016
rect 48282 12960 49800 13016
rect 48221 12958 49800 12960
rect 48221 12955 48287 12958
rect 49200 12868 49800 12958
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 43805 12474 43871 12477
rect 45553 12474 45619 12477
rect 43805 12472 45619 12474
rect 200 12188 800 12428
rect 43805 12416 43810 12472
rect 43866 12416 45558 12472
rect 45614 12416 45619 12472
rect 43805 12414 45619 12416
rect 43805 12411 43871 12414
rect 45553 12411 45619 12414
rect 48037 12338 48103 12341
rect 49200 12338 49800 12428
rect 48037 12336 49800 12338
rect 48037 12280 48042 12336
rect 48098 12280 49800 12336
rect 48037 12278 49800 12280
rect 48037 12275 48103 12278
rect 49200 12188 49800 12278
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 27153 11794 27219 11797
rect 28625 11794 28691 11797
rect 27153 11792 28691 11794
rect 200 11658 800 11748
rect 27153 11736 27158 11792
rect 27214 11736 28630 11792
rect 28686 11736 28691 11792
rect 27153 11734 28691 11736
rect 27153 11731 27219 11734
rect 28625 11731 28691 11734
rect 2773 11658 2839 11661
rect 200 11656 2839 11658
rect 200 11600 2778 11656
rect 2834 11600 2839 11656
rect 200 11598 2839 11600
rect 200 11508 800 11598
rect 2773 11595 2839 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 49200 10828 49800 11068
rect 200 10298 800 10388
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 3141 10298 3207 10301
rect 200 10296 3207 10298
rect 200 10240 3146 10296
rect 3202 10240 3207 10296
rect 200 10238 3207 10240
rect 200 10148 800 10238
rect 3141 10235 3207 10238
rect 49200 10148 49800 10388
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 200 9618 800 9708
rect 2773 9618 2839 9621
rect 200 9616 2839 9618
rect 200 9560 2778 9616
rect 2834 9560 2839 9616
rect 200 9558 2839 9560
rect 200 9468 800 9558
rect 2773 9555 2839 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 47945 8938 48011 8941
rect 49200 8938 49800 9028
rect 47945 8936 49800 8938
rect 47945 8880 47950 8936
rect 48006 8880 49800 8936
rect 47945 8878 49800 8880
rect 47945 8875 48011 8878
rect 49200 8788 49800 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 200 8108 800 8348
rect 47853 8258 47919 8261
rect 49200 8258 49800 8348
rect 47853 8256 49800 8258
rect 47853 8200 47858 8256
rect 47914 8200 49800 8256
rect 47853 8198 49800 8200
rect 47853 8195 47919 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 49200 8108 49800 8198
rect 200 7578 800 7668
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 2773 7578 2839 7581
rect 200 7576 2839 7578
rect 200 7520 2778 7576
rect 2834 7520 2839 7576
rect 200 7518 2839 7520
rect 200 7428 800 7518
rect 2773 7515 2839 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 200 6898 800 6988
rect 2773 6898 2839 6901
rect 200 6896 2839 6898
rect 200 6840 2778 6896
rect 2834 6840 2839 6896
rect 200 6838 2839 6840
rect 200 6748 800 6838
rect 2773 6835 2839 6838
rect 48221 6898 48287 6901
rect 49200 6898 49800 6988
rect 48221 6896 49800 6898
rect 48221 6840 48226 6896
rect 48282 6840 49800 6896
rect 48221 6838 49800 6840
rect 48221 6835 48287 6838
rect 49200 6748 49800 6838
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 49200 6068 49800 6308
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 200 5538 800 5628
rect 3509 5538 3575 5541
rect 200 5536 3575 5538
rect 200 5480 3514 5536
rect 3570 5480 3575 5536
rect 200 5478 3575 5480
rect 200 5388 800 5478
rect 3509 5475 3575 5478
rect 48221 5538 48287 5541
rect 49200 5538 49800 5628
rect 48221 5536 49800 5538
rect 48221 5480 48226 5536
rect 48282 5480 49800 5536
rect 48221 5478 49800 5480
rect 48221 5475 48287 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 49200 5388 49800 5478
rect 200 4858 800 4948
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 2957 4858 3023 4861
rect 200 4856 3023 4858
rect 200 4800 2962 4856
rect 3018 4800 3023 4856
rect 200 4798 3023 4800
rect 200 4708 800 4798
rect 2957 4795 3023 4798
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 49200 4028 49800 4268
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 200 3498 800 3588
rect 2773 3498 2839 3501
rect 200 3496 2839 3498
rect 200 3440 2778 3496
rect 2834 3440 2839 3496
rect 200 3438 2839 3440
rect 200 3348 800 3438
rect 2773 3435 2839 3438
rect 48037 3498 48103 3501
rect 49200 3498 49800 3588
rect 48037 3496 49800 3498
rect 48037 3440 48042 3496
rect 48098 3440 49800 3496
rect 48037 3438 49800 3440
rect 48037 3435 48103 3438
rect 49200 3348 49800 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 200 2818 800 2908
rect 2773 2818 2839 2821
rect 200 2816 2839 2818
rect 200 2760 2778 2816
rect 2834 2760 2839 2816
rect 200 2758 2839 2760
rect 200 2668 800 2758
rect 2773 2755 2839 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 46841 2138 46907 2141
rect 49200 2138 49800 2228
rect 46841 2136 49800 2138
rect 46841 2080 46846 2136
rect 46902 2080 49800 2136
rect 46841 2078 49800 2080
rect 46841 2075 46907 2078
rect 49200 1988 49800 2078
rect 200 1458 800 1548
rect 2865 1458 2931 1461
rect 200 1456 2931 1458
rect 200 1400 2870 1456
rect 2926 1400 2931 1456
rect 200 1398 2931 1400
rect 200 1308 800 1398
rect 2865 1395 2931 1398
rect 47209 1458 47275 1461
rect 49200 1458 49800 1548
rect 47209 1456 49800 1458
rect 47209 1400 47214 1456
rect 47270 1400 49800 1456
rect 47209 1398 49800 1400
rect 47209 1395 47275 1398
rect 49200 1308 49800 1398
rect 200 778 800 868
rect 2773 778 2839 781
rect 200 776 2839 778
rect 200 720 2778 776
rect 2834 720 2839 776
rect 200 718 2839 720
rect 200 628 800 718
rect 2773 715 2839 718
rect 48313 98 48379 101
rect 49200 98 49800 188
rect 48313 96 49800 98
rect 48313 40 48318 96
rect 48374 40 49800 96
rect 48313 38 49800 40
rect 48313 35 48379 38
rect 49200 -52 49800 38
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 20116 46956 20180 47020
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 20668 36000 20732 36004
rect 20668 35944 20682 36000
rect 20682 35944 20732 36000
rect 20668 35940 20732 35944
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 20668 31316 20732 31380
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 20116 24380 20180 24444
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 46816 19888 47376
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 20115 47020 20181 47021
rect 20115 46956 20116 47020
rect 20180 46956 20181 47020
rect 20115 46955 20181 46956
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 20118 24445 20178 46955
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 20667 36004 20733 36005
rect 20667 35940 20668 36004
rect 20732 35940 20733 36004
rect 20667 35939 20733 35940
rect 20670 31381 20730 35939
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 20667 31380 20733 31381
rect 20667 31316 20668 31380
rect 20732 31316 20733 31380
rect 20667 31315 20733 31316
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 20115 24444 20181 24445
rect 20115 24380 20116 24444
rect 20180 24380 20181 24444
rect 20115 24379 20181 24380
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17664 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1667941163
transform -1 0 17296 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1667941163
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1667941163
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1667941163
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1667941163
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119
timestamp 1667941163
transform 1 0 12052 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 13156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1667941163
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147
timestamp 1667941163
transform 1 0 14628 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_159
timestamp 1667941163
transform 1 0 15732 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1667941163
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_181
timestamp 1667941163
transform 1 0 17756 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_187
timestamp 1667941163
transform 1 0 18308 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_191
timestamp 1667941163
transform 1 0 18676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1667941163
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_202
timestamp 1667941163
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_212
timestamp 1667941163
transform 1 0 20608 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1667941163
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1667941163
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1667941163
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1667941163
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1667941163
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1667941163
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_315
timestamp 1667941163
transform 1 0 30084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_327
timestamp 1667941163
transform 1 0 31188 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1667941163
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1667941163
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1667941163
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1667941163
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1667941163
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_405
timestamp 1667941163
transform 1 0 38364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_413
timestamp 1667941163
transform 1 0 39100 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1667941163
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1667941163
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_433
timestamp 1667941163
transform 1 0 40940 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_439
timestamp 1667941163
transform 1 0 41492 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_443
timestamp 1667941163
transform 1 0 41860 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_447
timestamp 1667941163
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_449
timestamp 1667941163
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_461
timestamp 1667941163
transform 1 0 43516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_471
timestamp 1667941163
transform 1 0 44436 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1667941163
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_477
timestamp 1667941163
transform 1 0 44988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_502
timestamp 1667941163
transform 1 0 47288 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_505
timestamp 1667941163
transform 1 0 47564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_510
timestamp 1667941163
transform 1 0 48024 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7
timestamp 1667941163
transform 1 0 1748 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_29
timestamp 1667941163
transform 1 0 3772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1667941163
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_63
timestamp 1667941163
transform 1 0 6900 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_88
timestamp 1667941163
transform 1 0 9200 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_100
timestamp 1667941163
transform 1 0 10304 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1667941163
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1667941163
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_125
timestamp 1667941163
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_150
timestamp 1667941163
transform 1 0 14904 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_162
timestamp 1667941163
transform 1 0 16008 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_175
timestamp 1667941163
transform 1 0 17204 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_197
timestamp 1667941163
transform 1 0 19228 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1667941163
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1667941163
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_249
timestamp 1667941163
transform 1 0 24012 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1667941163
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_304
timestamp 1667941163
transform 1 0 29072 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_316
timestamp 1667941163
transform 1 0 30176 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_328
timestamp 1667941163
transform 1 0 31280 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_360
timestamp 1667941163
transform 1 0 34224 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_372
timestamp 1667941163
transform 1 0 35328 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_384
timestamp 1667941163
transform 1 0 36432 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_417
timestamp 1667941163
transform 1 0 39468 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_421
timestamp 1667941163
transform 1 0 39836 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_443
timestamp 1667941163
transform 1 0 41860 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1667941163
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_449
timestamp 1667941163
transform 1 0 42412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_472
timestamp 1667941163
transform 1 0 44528 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1667941163
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1667941163
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_505
timestamp 1667941163
transform 1 0 47564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_509
timestamp 1667941163
transform 1 0 47932 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_514
timestamp 1667941163
transform 1 0 48392 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_12
timestamp 1667941163
transform 1 0 2208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_19
timestamp 1667941163
transform 1 0 2852 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1667941163
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_35
timestamp 1667941163
transform 1 0 4324 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_42
timestamp 1667941163
transform 1 0 4968 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_49
timestamp 1667941163
transform 1 0 5612 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_74
timestamp 1667941163
transform 1 0 7912 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_81
timestamp 1667941163
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_101
timestamp 1667941163
transform 1 0 10396 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_123
timestamp 1667941163
transform 1 0 12420 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_132
timestamp 1667941163
transform 1 0 13248 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_153
timestamp 1667941163
transform 1 0 15180 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_161
timestamp 1667941163
transform 1 0 15916 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_166
timestamp 1667941163
transform 1 0 16376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_191
timestamp 1667941163
transform 1 0 18676 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1667941163
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_201
timestamp 1667941163
transform 1 0 19596 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_223
timestamp 1667941163
transform 1 0 21620 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_227
timestamp 1667941163
transform 1 0 21988 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_231
timestamp 1667941163
transform 1 0 22356 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_243
timestamp 1667941163
transform 1 0 23460 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1667941163
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_259
timestamp 1667941163
transform 1 0 24932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_266
timestamp 1667941163
transform 1 0 25576 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_291
timestamp 1667941163
transform 1 0 27876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_298
timestamp 1667941163
transform 1 0 28520 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp 1667941163
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_333
timestamp 1667941163
transform 1 0 31740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_337
timestamp 1667941163
transform 1 0 32108 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_344
timestamp 1667941163
transform 1 0 32752 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_356
timestamp 1667941163
transform 1 0 33856 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1667941163
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1667941163
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1667941163
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1667941163
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1667941163
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1667941163
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_426
timestamp 1667941163
transform 1 0 40296 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_430
timestamp 1667941163
transform 1 0 40664 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_452
timestamp 1667941163
transform 1 0 42688 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_459
timestamp 1667941163
transform 1 0 43332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_463
timestamp 1667941163
transform 1 0 43700 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_467
timestamp 1667941163
transform 1 0 44068 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_474
timestamp 1667941163
transform 1 0 44712 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_477
timestamp 1667941163
transform 1 0 44988 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_482
timestamp 1667941163
transform 1 0 45448 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_486
timestamp 1667941163
transform 1 0 45816 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_508
timestamp 1667941163
transform 1 0 47840 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_14
timestamp 1667941163
transform 1 0 2392 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_21
timestamp 1667941163
transform 1 0 3036 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_50
timestamp 1667941163
transform 1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_63
timestamp 1667941163
transform 1 0 6900 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_70
timestamp 1667941163
transform 1 0 7544 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_82
timestamp 1667941163
transform 1 0 8648 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_94
timestamp 1667941163
transform 1 0 9752 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1667941163
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1667941163
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_125
timestamp 1667941163
transform 1 0 12604 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_132
timestamp 1667941163
transform 1 0 13248 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_144
timestamp 1667941163
transform 1 0 14352 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_156
timestamp 1667941163
transform 1 0 15456 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_174
timestamp 1667941163
transform 1 0 17112 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_186
timestamp 1667941163
transform 1 0 18216 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_191
timestamp 1667941163
transform 1 0 18676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_197
timestamp 1667941163
transform 1 0 19228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_201
timestamp 1667941163
transform 1 0 19596 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_208
timestamp 1667941163
transform 1 0 20240 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_215
timestamp 1667941163
transform 1 0 20884 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1667941163
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_248
timestamp 1667941163
transform 1 0 23920 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_260
timestamp 1667941163
transform 1 0 25024 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_265
timestamp 1667941163
transform 1 0 25484 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_274
timestamp 1667941163
transform 1 0 26312 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_287
timestamp 1667941163
transform 1 0 27508 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_299
timestamp 1667941163
transform 1 0 28612 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_311
timestamp 1667941163
transform 1 0 29716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_323
timestamp 1667941163
transform 1 0 30820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1667941163
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1667941163
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1667941163
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1667941163
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_417
timestamp 1667941163
transform 1 0 39468 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_421
timestamp 1667941163
transform 1 0 39836 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_425
timestamp 1667941163
transform 1 0 40204 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_434
timestamp 1667941163
transform 1 0 41032 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1667941163
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1667941163
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_449
timestamp 1667941163
transform 1 0 42412 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_455
timestamp 1667941163
transform 1 0 42964 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_477
timestamp 1667941163
transform 1 0 44988 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_502
timestamp 1667941163
transform 1 0 47288 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_505
timestamp 1667941163
transform 1 0 47564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_510
timestamp 1667941163
transform 1 0 48024 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1667941163
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_34
timestamp 1667941163
transform 1 0 4232 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_43
timestamp 1667941163
transform 1 0 5060 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_59
timestamp 1667941163
transform 1 0 6532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_71
timestamp 1667941163
transform 1 0 7636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1667941163
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_93
timestamp 1667941163
transform 1 0 9660 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_116
timestamp 1667941163
transform 1 0 11776 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_128
timestamp 1667941163
transform 1 0 12880 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1667941163
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1667941163
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1667941163
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1667941163
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1667941163
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1667941163
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1667941163
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1667941163
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1667941163
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1667941163
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1667941163
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1667941163
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1667941163
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1667941163
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1667941163
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1667941163
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1667941163
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1667941163
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1667941163
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1667941163
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1667941163
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1667941163
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1667941163
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1667941163
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1667941163
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1667941163
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_457
timestamp 1667941163
transform 1 0 43148 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_463
timestamp 1667941163
transform 1 0 43700 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_467
timestamp 1667941163
transform 1 0 44068 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_474
timestamp 1667941163
transform 1 0 44712 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_477
timestamp 1667941163
transform 1 0 44988 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_500
timestamp 1667941163
transform 1 0 47104 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_507
timestamp 1667941163
transform 1 0 47748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_514
timestamp 1667941163
transform 1 0 48392 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_8
timestamp 1667941163
transform 1 0 1840 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_33
timestamp 1667941163
transform 1 0 4140 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_45
timestamp 1667941163
transform 1 0 5244 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1667941163
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1667941163
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1667941163
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1667941163
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1667941163
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1667941163
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1667941163
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1667941163
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1667941163
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1667941163
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1667941163
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1667941163
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1667941163
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1667941163
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1667941163
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1667941163
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1667941163
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1667941163
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1667941163
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1667941163
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1667941163
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1667941163
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1667941163
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1667941163
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1667941163
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1667941163
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1667941163
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_411
timestamp 1667941163
transform 1 0 38916 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_433
timestamp 1667941163
transform 1 0 40940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_445
timestamp 1667941163
transform 1 0 42044 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1667941163
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_461
timestamp 1667941163
transform 1 0 43516 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_470
timestamp 1667941163
transform 1 0 44344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_477
timestamp 1667941163
transform 1 0 44988 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_502
timestamp 1667941163
transform 1 0 47288 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_505
timestamp 1667941163
transform 1 0 47564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_510
timestamp 1667941163
transform 1 0 48024 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_9
timestamp 1667941163
transform 1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_16
timestamp 1667941163
transform 1 0 2576 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1667941163
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1667941163
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1667941163
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1667941163
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1667941163
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1667941163
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1667941163
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1667941163
transform 1 0 9476 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_95
timestamp 1667941163
transform 1 0 9844 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_102
timestamp 1667941163
transform 1 0 10488 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_114
timestamp 1667941163
transform 1 0 11592 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_126
timestamp 1667941163
transform 1 0 12696 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1667941163
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1667941163
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1667941163
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1667941163
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1667941163
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1667941163
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1667941163
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1667941163
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1667941163
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1667941163
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1667941163
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1667941163
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1667941163
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1667941163
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1667941163
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1667941163
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1667941163
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1667941163
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1667941163
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1667941163
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1667941163
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_401
timestamp 1667941163
transform 1 0 37996 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_409
timestamp 1667941163
transform 1 0 38732 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_415
timestamp 1667941163
transform 1 0 39284 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1667941163
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1667941163
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1667941163
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1667941163
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1667941163
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1667941163
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1667941163
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_477
timestamp 1667941163
transform 1 0 44988 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_485
timestamp 1667941163
transform 1 0 45724 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_489
timestamp 1667941163
transform 1 0 46092 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_514
timestamp 1667941163
transform 1 0 48392 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_14
timestamp 1667941163
transform 1 0 2392 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_21
timestamp 1667941163
transform 1 0 3036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_33
timestamp 1667941163
transform 1 0 4140 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_45
timestamp 1667941163
transform 1 0 5244 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_53
timestamp 1667941163
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1667941163
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1667941163
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1667941163
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1667941163
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1667941163
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1667941163
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1667941163
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1667941163
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1667941163
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1667941163
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1667941163
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1667941163
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1667941163
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1667941163
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1667941163
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1667941163
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1667941163
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1667941163
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1667941163
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1667941163
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1667941163
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1667941163
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1667941163
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1667941163
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1667941163
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1667941163
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1667941163
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1667941163
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_411
timestamp 1667941163
transform 1 0 38916 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_415
timestamp 1667941163
transform 1 0 39284 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_427
timestamp 1667941163
transform 1 0 40388 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_439
timestamp 1667941163
transform 1 0 41492 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1667941163
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1667941163
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1667941163
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1667941163
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_488
timestamp 1667941163
transform 1 0 46000 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_495
timestamp 1667941163
transform 1 0 46644 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_502
timestamp 1667941163
transform 1 0 47288 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_505
timestamp 1667941163
transform 1 0 47564 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_510
timestamp 1667941163
transform 1 0 48024 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1667941163
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1667941163
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1667941163
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1667941163
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1667941163
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1667941163
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1667941163
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1667941163
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1667941163
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1667941163
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1667941163
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1667941163
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1667941163
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1667941163
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1667941163
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1667941163
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1667941163
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1667941163
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1667941163
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1667941163
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1667941163
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1667941163
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1667941163
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1667941163
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1667941163
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1667941163
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1667941163
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1667941163
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1667941163
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1667941163
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1667941163
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1667941163
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1667941163
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1667941163
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1667941163
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1667941163
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1667941163
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1667941163
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1667941163
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_489
timestamp 1667941163
transform 1 0 46092 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_514
timestamp 1667941163
transform 1 0 48392 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_9
timestamp 1667941163
transform 1 0 1932 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_31
timestamp 1667941163
transform 1 0 3956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_43
timestamp 1667941163
transform 1 0 5060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1667941163
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1667941163
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1667941163
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1667941163
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1667941163
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1667941163
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1667941163
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1667941163
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1667941163
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1667941163
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1667941163
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1667941163
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1667941163
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1667941163
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1667941163
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1667941163
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1667941163
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1667941163
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1667941163
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1667941163
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1667941163
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1667941163
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1667941163
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1667941163
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1667941163
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1667941163
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1667941163
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1667941163
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1667941163
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1667941163
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1667941163
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1667941163
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1667941163
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1667941163
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1667941163
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1667941163
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1667941163
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1667941163
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_505
timestamp 1667941163
transform 1 0 47564 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_510
timestamp 1667941163
transform 1 0 48024 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_14
timestamp 1667941163
transform 1 0 2392 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_21
timestamp 1667941163
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1667941163
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1667941163
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1667941163
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1667941163
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1667941163
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1667941163
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1667941163
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1667941163
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1667941163
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1667941163
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1667941163
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1667941163
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1667941163
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1667941163
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1667941163
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1667941163
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1667941163
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1667941163
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1667941163
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1667941163
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1667941163
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1667941163
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1667941163
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1667941163
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1667941163
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1667941163
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1667941163
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1667941163
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1667941163
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1667941163
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1667941163
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1667941163
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1667941163
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1667941163
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1667941163
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1667941163
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1667941163
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1667941163
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1667941163
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1667941163
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1667941163
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1667941163
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_513
timestamp 1667941163
transform 1 0 48300 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1667941163
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1667941163
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1667941163
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1667941163
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1667941163
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1667941163
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1667941163
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1667941163
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1667941163
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1667941163
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1667941163
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1667941163
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1667941163
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1667941163
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1667941163
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1667941163
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1667941163
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1667941163
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1667941163
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1667941163
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1667941163
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1667941163
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1667941163
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1667941163
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1667941163
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1667941163
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1667941163
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1667941163
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1667941163
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1667941163
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1667941163
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1667941163
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1667941163
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1667941163
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1667941163
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1667941163
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1667941163
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1667941163
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1667941163
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1667941163
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_505
timestamp 1667941163
transform 1 0 47564 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_514
timestamp 1667941163
transform 1 0 48392 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_11
timestamp 1667941163
transform 1 0 2116 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1667941163
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1667941163
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1667941163
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1667941163
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1667941163
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1667941163
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1667941163
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1667941163
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1667941163
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1667941163
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1667941163
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1667941163
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1667941163
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1667941163
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1667941163
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1667941163
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1667941163
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1667941163
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1667941163
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1667941163
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1667941163
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1667941163
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1667941163
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1667941163
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1667941163
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1667941163
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1667941163
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_333
timestamp 1667941163
transform 1 0 31740 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_338
timestamp 1667941163
transform 1 0 32200 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_350
timestamp 1667941163
transform 1 0 33304 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_362
timestamp 1667941163
transform 1 0 34408 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1667941163
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1667941163
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_413
timestamp 1667941163
transform 1 0 39100 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_417
timestamp 1667941163
transform 1 0 39468 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1667941163
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1667941163
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1667941163
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_457
timestamp 1667941163
transform 1 0 43148 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_468
timestamp 1667941163
transform 1 0 44160 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1667941163
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1667941163
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_501
timestamp 1667941163
transform 1 0 47196 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_507
timestamp 1667941163
transform 1 0 47748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_514
timestamp 1667941163
transform 1 0 48392 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_9
timestamp 1667941163
transform 1 0 1932 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_31
timestamp 1667941163
transform 1 0 3956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_43
timestamp 1667941163
transform 1 0 5060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1667941163
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1667941163
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1667941163
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1667941163
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1667941163
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1667941163
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1667941163
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1667941163
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1667941163
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1667941163
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1667941163
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1667941163
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1667941163
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1667941163
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1667941163
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1667941163
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1667941163
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1667941163
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1667941163
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1667941163
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1667941163
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_289
timestamp 1667941163
transform 1 0 27692 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_294
timestamp 1667941163
transform 1 0 28152 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_305
timestamp 1667941163
transform 1 0 29164 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_315
timestamp 1667941163
transform 1 0 30084 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_327
timestamp 1667941163
transform 1 0 31188 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_334
timestamp 1667941163
transform 1 0 31832 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_346
timestamp 1667941163
transform 1 0 32936 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_358
timestamp 1667941163
transform 1 0 34040 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_370
timestamp 1667941163
transform 1 0 35144 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_380
timestamp 1667941163
transform 1 0 36064 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_411
timestamp 1667941163
transform 1 0 38916 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_418
timestamp 1667941163
transform 1 0 39560 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_424
timestamp 1667941163
transform 1 0 40112 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_433
timestamp 1667941163
transform 1 0 40940 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_444
timestamp 1667941163
transform 1 0 41952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_449
timestamp 1667941163
transform 1 0 42412 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_467
timestamp 1667941163
transform 1 0 44068 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_478
timestamp 1667941163
transform 1 0 45080 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_490
timestamp 1667941163
transform 1 0 46184 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_502
timestamp 1667941163
transform 1 0 47288 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_505
timestamp 1667941163
transform 1 0 47564 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_513
timestamp 1667941163
transform 1 0 48300 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_14
timestamp 1667941163
transform 1 0 2392 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1667941163
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1667941163
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1667941163
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1667941163
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1667941163
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1667941163
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1667941163
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1667941163
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1667941163
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1667941163
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1667941163
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1667941163
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1667941163
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1667941163
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1667941163
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1667941163
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1667941163
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_221
timestamp 1667941163
transform 1 0 21436 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_241
timestamp 1667941163
transform 1 0 23276 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_249
timestamp 1667941163
transform 1 0 24012 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_261
timestamp 1667941163
transform 1 0 25116 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_269
timestamp 1667941163
transform 1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_288
timestamp 1667941163
transform 1 0 27600 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_295
timestamp 1667941163
transform 1 0 28244 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_306
timestamp 1667941163
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_317
timestamp 1667941163
transform 1 0 30268 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_321
timestamp 1667941163
transform 1 0 30636 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_326
timestamp 1667941163
transform 1 0 31096 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_337
timestamp 1667941163
transform 1 0 32108 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_343
timestamp 1667941163
transform 1 0 32660 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_351
timestamp 1667941163
transform 1 0 33396 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_361
timestamp 1667941163
transform 1 0 34316 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_383
timestamp 1667941163
transform 1 0 36340 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_395
timestamp 1667941163
transform 1 0 37444 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_409
timestamp 1667941163
transform 1 0 38732 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_418
timestamp 1667941163
transform 1 0 39560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_421
timestamp 1667941163
transform 1 0 39836 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_441
timestamp 1667941163
transform 1 0 41676 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_448
timestamp 1667941163
transform 1 0 42320 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_456
timestamp 1667941163
transform 1 0 43056 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_466
timestamp 1667941163
transform 1 0 43976 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_474
timestamp 1667941163
transform 1 0 44712 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_477
timestamp 1667941163
transform 1 0 44988 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_484
timestamp 1667941163
transform 1 0 45632 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_496
timestamp 1667941163
transform 1 0 46736 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_508
timestamp 1667941163
transform 1 0 47840 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_15
timestamp 1667941163
transform 1 0 2484 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_38
timestamp 1667941163
transform 1 0 4600 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_50
timestamp 1667941163
transform 1 0 5704 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1667941163
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1667941163
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1667941163
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1667941163
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1667941163
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1667941163
transform 1 0 12236 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_143
timestamp 1667941163
transform 1 0 14260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_155
timestamp 1667941163
transform 1 0 15364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1667941163
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1667941163
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1667941163
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1667941163
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1667941163
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1667941163
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_231
timestamp 1667941163
transform 1 0 22356 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_238
timestamp 1667941163
transform 1 0 23000 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_246
timestamp 1667941163
transform 1 0 23736 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_264
timestamp 1667941163
transform 1 0 25392 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_276
timestamp 1667941163
transform 1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_292
timestamp 1667941163
transform 1 0 27968 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_300
timestamp 1667941163
transform 1 0 28704 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_305
timestamp 1667941163
transform 1 0 29164 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_309
timestamp 1667941163
transform 1 0 29532 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_315
timestamp 1667941163
transform 1 0 30084 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_321
timestamp 1667941163
transform 1 0 30636 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_325
timestamp 1667941163
transform 1 0 31004 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_334
timestamp 1667941163
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_352
timestamp 1667941163
transform 1 0 33488 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_364
timestamp 1667941163
transform 1 0 34592 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_379
timestamp 1667941163
transform 1 0 35972 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_385
timestamp 1667941163
transform 1 0 36524 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_390
timestamp 1667941163
transform 1 0 36984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_397
timestamp 1667941163
transform 1 0 37628 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_404
timestamp 1667941163
transform 1 0 38272 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_417
timestamp 1667941163
transform 1 0 39468 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_423
timestamp 1667941163
transform 1 0 40020 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_430
timestamp 1667941163
transform 1 0 40664 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_438
timestamp 1667941163
transform 1 0 41400 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_446
timestamp 1667941163
transform 1 0 42136 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1667941163
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_461
timestamp 1667941163
transform 1 0 43516 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_472
timestamp 1667941163
transform 1 0 44528 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_479
timestamp 1667941163
transform 1 0 45172 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_483
timestamp 1667941163
transform 1 0 45540 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_500
timestamp 1667941163
transform 1 0 47104 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_505
timestamp 1667941163
transform 1 0 47564 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_513
timestamp 1667941163
transform 1 0 48300 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_11
timestamp 1667941163
transform 1 0 2116 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_15
timestamp 1667941163
transform 1 0 2484 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_22
timestamp 1667941163
transform 1 0 3128 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_34
timestamp 1667941163
transform 1 0 4232 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_46
timestamp 1667941163
transform 1 0 5336 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_58
timestamp 1667941163
transform 1 0 6440 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_70
timestamp 1667941163
transform 1 0 7544 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1667941163
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1667941163
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1667941163
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_121
timestamp 1667941163
transform 1 0 12236 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_125
timestamp 1667941163
transform 1 0 12604 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_132
timestamp 1667941163
transform 1 0 13248 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1667941163
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1667941163
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1667941163
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1667941163
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1667941163
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1667941163
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_221
timestamp 1667941163
transform 1 0 21436 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_225
timestamp 1667941163
transform 1 0 21804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_242
timestamp 1667941163
transform 1 0 23368 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1667941163
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_272
timestamp 1667941163
transform 1 0 26128 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_284
timestamp 1667941163
transform 1 0 27232 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_290
timestamp 1667941163
transform 1 0 27784 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_299
timestamp 1667941163
transform 1 0 28612 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 1667941163
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_315
timestamp 1667941163
transform 1 0 30084 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_323
timestamp 1667941163
transform 1 0 30820 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_341
timestamp 1667941163
transform 1 0 32476 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_347
timestamp 1667941163
transform 1 0 33028 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_351
timestamp 1667941163
transform 1 0 33396 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_358
timestamp 1667941163
transform 1 0 34040 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_369
timestamp 1667941163
transform 1 0 35052 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_390
timestamp 1667941163
transform 1 0 36984 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_418
timestamp 1667941163
transform 1 0 39560 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1667941163
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1667941163
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_445
timestamp 1667941163
transform 1 0 42044 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_453
timestamp 1667941163
transform 1 0 42780 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_462
timestamp 1667941163
transform 1 0 43608 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_468
timestamp 1667941163
transform 1 0 44160 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_474
timestamp 1667941163
transform 1 0 44712 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_477
timestamp 1667941163
transform 1 0 44988 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_486
timestamp 1667941163
transform 1 0 45816 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_498
timestamp 1667941163
transform 1 0 46920 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_510
timestamp 1667941163
transform 1 0 48024 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_9
timestamp 1667941163
transform 1 0 1932 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_31
timestamp 1667941163
transform 1 0 3956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_43
timestamp 1667941163
transform 1 0 5060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1667941163
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1667941163
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1667941163
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1667941163
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1667941163
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1667941163
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1667941163
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1667941163
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1667941163
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1667941163
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1667941163
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1667941163
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1667941163
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1667941163
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1667941163
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1667941163
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_229
timestamp 1667941163
transform 1 0 22172 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_238
timestamp 1667941163
transform 1 0 23000 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_250
timestamp 1667941163
transform 1 0 24104 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_260
timestamp 1667941163
transform 1 0 25024 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_270
timestamp 1667941163
transform 1 0 25944 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1667941163
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_292
timestamp 1667941163
transform 1 0 27968 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_298
timestamp 1667941163
transform 1 0 28520 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_305
timestamp 1667941163
transform 1 0 29164 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_315
timestamp 1667941163
transform 1 0 30084 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_325
timestamp 1667941163
transform 1 0 31004 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_333
timestamp 1667941163
transform 1 0 31740 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_346
timestamp 1667941163
transform 1 0 32936 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_354
timestamp 1667941163
transform 1 0 33672 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_358
timestamp 1667941163
transform 1 0 34040 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_370
timestamp 1667941163
transform 1 0 35144 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_382
timestamp 1667941163
transform 1 0 36248 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_390
timestamp 1667941163
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_400
timestamp 1667941163
transform 1 0 37904 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_404
timestamp 1667941163
transform 1 0 38272 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_409
timestamp 1667941163
transform 1 0 38732 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_421
timestamp 1667941163
transform 1 0 39836 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_433
timestamp 1667941163
transform 1 0 40940 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_445
timestamp 1667941163
transform 1 0 42044 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_449
timestamp 1667941163
transform 1 0 42412 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_457
timestamp 1667941163
transform 1 0 43148 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_461
timestamp 1667941163
transform 1 0 43516 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_466
timestamp 1667941163
transform 1 0 43976 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_477
timestamp 1667941163
transform 1 0 44988 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_489
timestamp 1667941163
transform 1 0 46092 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_501
timestamp 1667941163
transform 1 0 47196 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_505
timestamp 1667941163
transform 1 0 47564 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_513
timestamp 1667941163
transform 1 0 48300 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_9
timestamp 1667941163
transform 1 0 1932 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_13
timestamp 1667941163
transform 1 0 2300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_25
timestamp 1667941163
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1667941163
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1667941163
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1667941163
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1667941163
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1667941163
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1667941163
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1667941163
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1667941163
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1667941163
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1667941163
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1667941163
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1667941163
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1667941163
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1667941163
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1667941163
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_209
timestamp 1667941163
transform 1 0 20332 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_229
timestamp 1667941163
transform 1 0 22172 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_241
timestamp 1667941163
transform 1 0 23276 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_249
timestamp 1667941163
transform 1 0 24012 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_259
timestamp 1667941163
transform 1 0 24932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_268
timestamp 1667941163
transform 1 0 25760 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_292
timestamp 1667941163
transform 1 0 27968 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_304
timestamp 1667941163
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1667941163
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1667941163
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_345
timestamp 1667941163
transform 1 0 32844 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_353
timestamp 1667941163
transform 1 0 33580 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_362
timestamp 1667941163
transform 1 0 34408 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_386
timestamp 1667941163
transform 1 0 36616 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_393
timestamp 1667941163
transform 1 0 37260 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_405
timestamp 1667941163
transform 1 0 38364 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_417
timestamp 1667941163
transform 1 0 39468 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1667941163
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_439
timestamp 1667941163
transform 1 0 41492 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_451
timestamp 1667941163
transform 1 0 42596 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_459
timestamp 1667941163
transform 1 0 43332 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_468
timestamp 1667941163
transform 1 0 44160 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1667941163
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_489
timestamp 1667941163
transform 1 0 46092 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_514
timestamp 1667941163
transform 1 0 48392 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1667941163
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1667941163
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1667941163
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1667941163
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1667941163
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1667941163
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1667941163
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1667941163
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1667941163
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1667941163
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1667941163
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1667941163
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1667941163
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1667941163
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1667941163
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1667941163
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1667941163
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1667941163
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1667941163
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1667941163
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_235
timestamp 1667941163
transform 1 0 22724 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_247
timestamp 1667941163
transform 1 0 23828 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_259
timestamp 1667941163
transform 1 0 24932 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_271
timestamp 1667941163
transform 1 0 26036 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1667941163
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1667941163
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1667941163
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1667941163
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1667941163
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_352
timestamp 1667941163
transform 1 0 33488 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_372
timestamp 1667941163
transform 1 0 35328 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_380
timestamp 1667941163
transform 1 0 36064 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_388
timestamp 1667941163
transform 1 0 36800 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_398
timestamp 1667941163
transform 1 0 37720 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_410
timestamp 1667941163
transform 1 0 38824 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_422
timestamp 1667941163
transform 1 0 39928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_431
timestamp 1667941163
transform 1 0 40756 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_443
timestamp 1667941163
transform 1 0 41860 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1667941163
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_449
timestamp 1667941163
transform 1 0 42412 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_453
timestamp 1667941163
transform 1 0 42780 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_458
timestamp 1667941163
transform 1 0 43240 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_466
timestamp 1667941163
transform 1 0 43976 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_472
timestamp 1667941163
transform 1 0 44528 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_479
timestamp 1667941163
transform 1 0 45172 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_491
timestamp 1667941163
transform 1 0 46276 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_502
timestamp 1667941163
transform 1 0 47288 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_505
timestamp 1667941163
transform 1 0 47564 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_510
timestamp 1667941163
transform 1 0 48024 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1667941163
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1667941163
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1667941163
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1667941163
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1667941163
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1667941163
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1667941163
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1667941163
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1667941163
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1667941163
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1667941163
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1667941163
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1667941163
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1667941163
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1667941163
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1667941163
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1667941163
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_209
timestamp 1667941163
transform 1 0 20332 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1667941163
transform 1 0 20700 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_230
timestamp 1667941163
transform 1 0 22264 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_240
timestamp 1667941163
transform 1 0 23184 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1667941163
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_277
timestamp 1667941163
transform 1 0 26588 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_285
timestamp 1667941163
transform 1 0 27324 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_296
timestamp 1667941163
transform 1 0 28336 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_317
timestamp 1667941163
transform 1 0 30268 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_326
timestamp 1667941163
transform 1 0 31096 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_346
timestamp 1667941163
transform 1 0 32936 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_356
timestamp 1667941163
transform 1 0 33856 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_397
timestamp 1667941163
transform 1 0 37628 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_406
timestamp 1667941163
transform 1 0 38456 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_418
timestamp 1667941163
transform 1 0 39560 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_421
timestamp 1667941163
transform 1 0 39836 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_435
timestamp 1667941163
transform 1 0 41124 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_443
timestamp 1667941163
transform 1 0 41860 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_450
timestamp 1667941163
transform 1 0 42504 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_458
timestamp 1667941163
transform 1 0 43240 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_464
timestamp 1667941163
transform 1 0 43792 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_471
timestamp 1667941163
transform 1 0 44436 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1667941163
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_477
timestamp 1667941163
transform 1 0 44988 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_486
timestamp 1667941163
transform 1 0 45816 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_492
timestamp 1667941163
transform 1 0 46368 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_514
timestamp 1667941163
transform 1 0 48392 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_14
timestamp 1667941163
transform 1 0 2392 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_21
timestamp 1667941163
transform 1 0 3036 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_33
timestamp 1667941163
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_45
timestamp 1667941163
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1667941163
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1667941163
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1667941163
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1667941163
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1667941163
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1667941163
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1667941163
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1667941163
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1667941163
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1667941163
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1667941163
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1667941163
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_205
timestamp 1667941163
transform 1 0 19964 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_213
timestamp 1667941163
transform 1 0 20700 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1667941163
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_235
timestamp 1667941163
transform 1 0 22724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_247
timestamp 1667941163
transform 1 0 23828 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_251
timestamp 1667941163
transform 1 0 24196 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_268
timestamp 1667941163
transform 1 0 25760 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_277
timestamp 1667941163
transform 1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_299
timestamp 1667941163
transform 1 0 28612 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_327
timestamp 1667941163
transform 1 0 31188 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1667941163
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_355
timestamp 1667941163
transform 1 0 33764 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_367
timestamp 1667941163
transform 1 0 34868 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_379
timestamp 1667941163
transform 1 0 35972 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1667941163
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_411
timestamp 1667941163
transform 1 0 38916 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_415
timestamp 1667941163
transform 1 0 39284 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_432
timestamp 1667941163
transform 1 0 40848 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_442
timestamp 1667941163
transform 1 0 41768 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_449
timestamp 1667941163
transform 1 0 42412 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_457
timestamp 1667941163
transform 1 0 43148 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_465
timestamp 1667941163
transform 1 0 43884 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_474
timestamp 1667941163
transform 1 0 44712 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_478
timestamp 1667941163
transform 1 0 45080 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_495
timestamp 1667941163
transform 1 0 46644 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_502
timestamp 1667941163
transform 1 0 47288 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_505
timestamp 1667941163
transform 1 0 47564 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_510
timestamp 1667941163
transform 1 0 48024 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1667941163
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_34
timestamp 1667941163
transform 1 0 4232 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_46
timestamp 1667941163
transform 1 0 5336 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_58
timestamp 1667941163
transform 1 0 6440 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_70
timestamp 1667941163
transform 1 0 7544 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1667941163
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1667941163
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1667941163
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1667941163
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1667941163
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1667941163
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_153
timestamp 1667941163
transform 1 0 15180 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_161
timestamp 1667941163
transform 1 0 15916 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_178
timestamp 1667941163
transform 1 0 17480 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_190
timestamp 1667941163
transform 1 0 18584 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1667941163
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1667941163
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_233
timestamp 1667941163
transform 1 0 22540 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_239
timestamp 1667941163
transform 1 0 23092 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_246
timestamp 1667941163
transform 1 0 23736 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_262
timestamp 1667941163
transform 1 0 25208 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_279
timestamp 1667941163
transform 1 0 26772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_289
timestamp 1667941163
transform 1 0 27692 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_297
timestamp 1667941163
transform 1 0 28428 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1667941163
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_317
timestamp 1667941163
transform 1 0 30268 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_329
timestamp 1667941163
transform 1 0 31372 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_337
timestamp 1667941163
transform 1 0 32108 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_345
timestamp 1667941163
transform 1 0 32844 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1667941163
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1667941163
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_389
timestamp 1667941163
transform 1 0 36892 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_397
timestamp 1667941163
transform 1 0 37628 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_405
timestamp 1667941163
transform 1 0 38364 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1667941163
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1667941163
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_421
timestamp 1667941163
transform 1 0 39836 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_429
timestamp 1667941163
transform 1 0 40572 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_436
timestamp 1667941163
transform 1 0 41216 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_448
timestamp 1667941163
transform 1 0 42320 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_456
timestamp 1667941163
transform 1 0 43056 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_465
timestamp 1667941163
transform 1 0 43884 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_474
timestamp 1667941163
transform 1 0 44712 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1667941163
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1667941163
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1667941163
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_513
timestamp 1667941163
transform 1 0 48300 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_14
timestamp 1667941163
transform 1 0 2392 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_21
timestamp 1667941163
transform 1 0 3036 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_50
timestamp 1667941163
transform 1 0 5704 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1667941163
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1667941163
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1667941163
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1667941163
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1667941163
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1667941163
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_137
timestamp 1667941163
transform 1 0 13708 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_154
timestamp 1667941163
transform 1 0 15272 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_162
timestamp 1667941163
transform 1 0 16008 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1667941163
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_177
timestamp 1667941163
transform 1 0 17388 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1667941163
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1667941163
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1667941163
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_237
timestamp 1667941163
transform 1 0 22908 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_248
timestamp 1667941163
transform 1 0 23920 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_260
timestamp 1667941163
transform 1 0 25024 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_272
timestamp 1667941163
transform 1 0 26128 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_286
timestamp 1667941163
transform 1 0 27416 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_298
timestamp 1667941163
transform 1 0 28520 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_316
timestamp 1667941163
transform 1 0 30176 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_328
timestamp 1667941163
transform 1 0 31280 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_347
timestamp 1667941163
transform 1 0 33028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_359
timestamp 1667941163
transform 1 0 34132 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_377
timestamp 1667941163
transform 1 0 35788 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_389
timestamp 1667941163
transform 1 0 36892 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_411
timestamp 1667941163
transform 1 0 38916 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_423
timestamp 1667941163
transform 1 0 40020 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1667941163
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1667941163
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1667941163
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_449
timestamp 1667941163
transform 1 0 42412 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_455
timestamp 1667941163
transform 1 0 42964 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_464
timestamp 1667941163
transform 1 0 43792 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_472
timestamp 1667941163
transform 1 0 44528 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_484
timestamp 1667941163
transform 1 0 45632 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_496
timestamp 1667941163
transform 1 0 46736 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_502
timestamp 1667941163
transform 1 0 47288 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_505
timestamp 1667941163
transform 1 0 47564 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_510
timestamp 1667941163
transform 1 0 48024 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1667941163
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1667941163
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1667941163
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1667941163
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1667941163
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1667941163
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1667941163
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1667941163
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_121
timestamp 1667941163
transform 1 0 12236 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_127
timestamp 1667941163
transform 1 0 12788 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_131
timestamp 1667941163
transform 1 0 13156 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1667941163
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_145
timestamp 1667941163
transform 1 0 14444 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_155
timestamp 1667941163
transform 1 0 15364 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_167
timestamp 1667941163
transform 1 0 16468 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_182
timestamp 1667941163
transform 1 0 17848 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_188
timestamp 1667941163
transform 1 0 18400 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1667941163
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_208
timestamp 1667941163
transform 1 0 20240 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_220
timestamp 1667941163
transform 1 0 21344 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_232
timestamp 1667941163
transform 1 0 22448 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1667941163
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_261
timestamp 1667941163
transform 1 0 25116 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_269
timestamp 1667941163
transform 1 0 25852 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_276
timestamp 1667941163
transform 1 0 26496 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_283
timestamp 1667941163
transform 1 0 27140 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_294
timestamp 1667941163
transform 1 0 28152 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1667941163
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1667941163
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_317
timestamp 1667941163
transform 1 0 30268 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_325
timestamp 1667941163
transform 1 0 31004 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_337
timestamp 1667941163
transform 1 0 32108 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_349
timestamp 1667941163
transform 1 0 33212 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_361
timestamp 1667941163
transform 1 0 34316 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_374
timestamp 1667941163
transform 1 0 35512 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_386
timestamp 1667941163
transform 1 0 36616 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_398
timestamp 1667941163
transform 1 0 37720 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_410
timestamp 1667941163
transform 1 0 38824 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_414
timestamp 1667941163
transform 1 0 39192 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_418
timestamp 1667941163
transform 1 0 39560 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_421
timestamp 1667941163
transform 1 0 39836 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_434
timestamp 1667941163
transform 1 0 41032 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_445
timestamp 1667941163
transform 1 0 42044 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_451
timestamp 1667941163
transform 1 0 42596 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_468
timestamp 1667941163
transform 1 0 44160 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1667941163
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_489
timestamp 1667941163
transform 1 0 46092 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_514
timestamp 1667941163
transform 1 0 48392 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_18
timestamp 1667941163
transform 1 0 2760 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_30
timestamp 1667941163
transform 1 0 3864 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_42
timestamp 1667941163
transform 1 0 4968 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1667941163
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1667941163
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1667941163
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1667941163
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1667941163
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1667941163
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_135
timestamp 1667941163
transform 1 0 13524 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_143
timestamp 1667941163
transform 1 0 14260 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_153
timestamp 1667941163
transform 1 0 15180 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_165
timestamp 1667941163
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_173
timestamp 1667941163
transform 1 0 17020 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_183
timestamp 1667941163
transform 1 0 17940 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_192
timestamp 1667941163
transform 1 0 18768 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_199
timestamp 1667941163
transform 1 0 19412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_211
timestamp 1667941163
transform 1 0 20516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1667941163
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_235
timestamp 1667941163
transform 1 0 22724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_247
timestamp 1667941163
transform 1 0 23828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_256
timestamp 1667941163
transform 1 0 24656 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_263
timestamp 1667941163
transform 1 0 25300 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_274
timestamp 1667941163
transform 1 0 26312 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1667941163
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1667941163
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_317
timestamp 1667941163
transform 1 0 30268 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_331
timestamp 1667941163
transform 1 0 31556 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1667941163
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_345
timestamp 1667941163
transform 1 0 32844 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_355
timestamp 1667941163
transform 1 0 33764 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_363
timestamp 1667941163
transform 1 0 34500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_370
timestamp 1667941163
transform 1 0 35144 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_378
timestamp 1667941163
transform 1 0 35880 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_390
timestamp 1667941163
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_417
timestamp 1667941163
transform 1 0 39468 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_436
timestamp 1667941163
transform 1 0 41216 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_443
timestamp 1667941163
transform 1 0 41860 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1667941163
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_449
timestamp 1667941163
transform 1 0 42412 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_456
timestamp 1667941163
transform 1 0 43056 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_468
timestamp 1667941163
transform 1 0 44160 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_480
timestamp 1667941163
transform 1 0 45264 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_492
timestamp 1667941163
transform 1 0 46368 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_498
timestamp 1667941163
transform 1 0 46920 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_502
timestamp 1667941163
transform 1 0 47288 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_505
timestamp 1667941163
transform 1 0 47564 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_510
timestamp 1667941163
transform 1 0 48024 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1667941163
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1667941163
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1667941163
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1667941163
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1667941163
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1667941163
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1667941163
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1667941163
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_121
timestamp 1667941163
transform 1 0 12236 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_125
timestamp 1667941163
transform 1 0 12604 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_135
timestamp 1667941163
transform 1 0 13524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1667941163
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1667941163
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_165
timestamp 1667941163
transform 1 0 16284 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_182
timestamp 1667941163
transform 1 0 17848 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1667941163
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_209
timestamp 1667941163
transform 1 0 20332 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_213
timestamp 1667941163
transform 1 0 20700 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_230
timestamp 1667941163
transform 1 0 22264 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_242
timestamp 1667941163
transform 1 0 23368 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_246
timestamp 1667941163
transform 1 0 23736 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_264
timestamp 1667941163
transform 1 0 25392 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_268
timestamp 1667941163
transform 1 0 25760 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_274
timestamp 1667941163
transform 1 0 26312 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_286
timestamp 1667941163
transform 1 0 27416 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_295
timestamp 1667941163
transform 1 0 28244 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1667941163
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_333
timestamp 1667941163
transform 1 0 31740 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_353
timestamp 1667941163
transform 1 0 33580 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_357
timestamp 1667941163
transform 1 0 33948 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_362
timestamp 1667941163
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_372
timestamp 1667941163
transform 1 0 35328 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_379
timestamp 1667941163
transform 1 0 35972 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_385
timestamp 1667941163
transform 1 0 36524 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_390
timestamp 1667941163
transform 1 0 36984 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_398
timestamp 1667941163
transform 1 0 37720 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_406
timestamp 1667941163
transform 1 0 38456 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_418
timestamp 1667941163
transform 1 0 39560 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1667941163
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1667941163
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1667941163
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_457
timestamp 1667941163
transform 1 0 43148 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_463
timestamp 1667941163
transform 1 0 43700 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1667941163
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1667941163
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_489
timestamp 1667941163
transform 1 0 46092 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_514
timestamp 1667941163
transform 1 0 48392 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_14
timestamp 1667941163
transform 1 0 2392 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_26
timestamp 1667941163
transform 1 0 3496 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_38
timestamp 1667941163
transform 1 0 4600 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_50
timestamp 1667941163
transform 1 0 5704 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1667941163
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1667941163
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1667941163
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1667941163
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1667941163
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_122
timestamp 1667941163
transform 1 0 12328 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_130
timestamp 1667941163
transform 1 0 13064 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_139
timestamp 1667941163
transform 1 0 13892 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_159
timestamp 1667941163
transform 1 0 15732 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1667941163
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_174
timestamp 1667941163
transform 1 0 17112 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_186
timestamp 1667941163
transform 1 0 18216 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_204
timestamp 1667941163
transform 1 0 19872 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_216
timestamp 1667941163
transform 1 0 20976 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_233
timestamp 1667941163
transform 1 0 22540 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_237
timestamp 1667941163
transform 1 0 22908 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_254
timestamp 1667941163
transform 1 0 24472 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_267
timestamp 1667941163
transform 1 0 25668 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_277
timestamp 1667941163
transform 1 0 26588 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1667941163
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1667941163
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_317
timestamp 1667941163
transform 1 0 30268 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_331
timestamp 1667941163
transform 1 0 31556 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1667941163
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_355
timestamp 1667941163
transform 1 0 33764 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_360
timestamp 1667941163
transform 1 0 34224 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_369
timestamp 1667941163
transform 1 0 35052 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_378
timestamp 1667941163
transform 1 0 35880 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_382
timestamp 1667941163
transform 1 0 36248 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_390
timestamp 1667941163
transform 1 0 36984 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_411
timestamp 1667941163
transform 1 0 38916 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_418
timestamp 1667941163
transform 1 0 39560 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_430
timestamp 1667941163
transform 1 0 40664 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_443
timestamp 1667941163
transform 1 0 41860 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1667941163
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_449
timestamp 1667941163
transform 1 0 42412 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_457
timestamp 1667941163
transform 1 0 43148 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_477
timestamp 1667941163
transform 1 0 44988 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_502
timestamp 1667941163
transform 1 0 47288 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_505
timestamp 1667941163
transform 1 0 47564 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_510
timestamp 1667941163
transform 1 0 48024 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_11
timestamp 1667941163
transform 1 0 2116 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1667941163
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1667941163
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1667941163
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1667941163
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1667941163
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1667941163
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1667941163
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1667941163
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_109
timestamp 1667941163
transform 1 0 11132 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_129
timestamp 1667941163
transform 1 0 12972 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp 1667941163
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_149
timestamp 1667941163
transform 1 0 14812 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_154
timestamp 1667941163
transform 1 0 15272 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_166
timestamp 1667941163
transform 1 0 16376 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_178
timestamp 1667941163
transform 1 0 17480 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_186
timestamp 1667941163
transform 1 0 18216 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1667941163
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_202
timestamp 1667941163
transform 1 0 19688 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_214
timestamp 1667941163
transform 1 0 20792 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_226
timestamp 1667941163
transform 1 0 21896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_238
timestamp 1667941163
transform 1 0 23000 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_248
timestamp 1667941163
transform 1 0 23920 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1667941163
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1667941163
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_289
timestamp 1667941163
transform 1 0 27692 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_297
timestamp 1667941163
transform 1 0 28428 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_305
timestamp 1667941163
transform 1 0 29164 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_321
timestamp 1667941163
transform 1 0 30636 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_331
timestamp 1667941163
transform 1 0 31556 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_343
timestamp 1667941163
transform 1 0 32660 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_355
timestamp 1667941163
transform 1 0 33764 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1667941163
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_371
timestamp 1667941163
transform 1 0 35236 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_380
timestamp 1667941163
transform 1 0 36064 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_386
timestamp 1667941163
transform 1 0 36616 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_394
timestamp 1667941163
transform 1 0 37352 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_418
timestamp 1667941163
transform 1 0 39560 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_421
timestamp 1667941163
transform 1 0 39836 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_429
timestamp 1667941163
transform 1 0 40572 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_435
timestamp 1667941163
transform 1 0 41124 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_445
timestamp 1667941163
transform 1 0 42044 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_462
timestamp 1667941163
transform 1 0 43608 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_471
timestamp 1667941163
transform 1 0 44436 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1667941163
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1667941163
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_489
timestamp 1667941163
transform 1 0 46092 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_514
timestamp 1667941163
transform 1 0 48392 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_9
timestamp 1667941163
transform 1 0 1932 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_31
timestamp 1667941163
transform 1 0 3956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_43
timestamp 1667941163
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1667941163
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1667941163
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1667941163
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1667941163
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1667941163
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1667941163
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_130
timestamp 1667941163
transform 1 0 13064 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_142
timestamp 1667941163
transform 1 0 14168 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_154
timestamp 1667941163
transform 1 0 15272 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1667941163
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_181
timestamp 1667941163
transform 1 0 17756 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_189
timestamp 1667941163
transform 1 0 18492 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_200
timestamp 1667941163
transform 1 0 19504 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_212
timestamp 1667941163
transform 1 0 20608 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_229
timestamp 1667941163
transform 1 0 22172 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_238
timestamp 1667941163
transform 1 0 23000 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_258
timestamp 1667941163
transform 1 0 24840 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_270
timestamp 1667941163
transform 1 0 25944 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_274
timestamp 1667941163
transform 1 0 26312 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1667941163
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_294
timestamp 1667941163
transform 1 0 28152 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_303
timestamp 1667941163
transform 1 0 28980 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_315
timestamp 1667941163
transform 1 0 30084 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 1667941163
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_343
timestamp 1667941163
transform 1 0 32660 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_351
timestamp 1667941163
transform 1 0 33396 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_360
timestamp 1667941163
transform 1 0 34224 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_372
timestamp 1667941163
transform 1 0 35328 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_388
timestamp 1667941163
transform 1 0 36800 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_401
timestamp 1667941163
transform 1 0 37996 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_405
timestamp 1667941163
transform 1 0 38364 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_414
timestamp 1667941163
transform 1 0 39192 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_426
timestamp 1667941163
transform 1 0 40296 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_443
timestamp 1667941163
transform 1 0 41860 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1667941163
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_449
timestamp 1667941163
transform 1 0 42412 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_456
timestamp 1667941163
transform 1 0 43056 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_465
timestamp 1667941163
transform 1 0 43884 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_473
timestamp 1667941163
transform 1 0 44620 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_492
timestamp 1667941163
transform 1 0 46368 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_499
timestamp 1667941163
transform 1 0 47012 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1667941163
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_505
timestamp 1667941163
transform 1 0 47564 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_510
timestamp 1667941163
transform 1 0 48024 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_9
timestamp 1667941163
transform 1 0 1932 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_13
timestamp 1667941163
transform 1 0 2300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_25
timestamp 1667941163
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1667941163
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1667941163
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1667941163
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1667941163
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1667941163
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1667941163
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_109
timestamp 1667941163
transform 1 0 11132 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_118
timestamp 1667941163
transform 1 0 11960 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_122
timestamp 1667941163
transform 1 0 12328 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_130
timestamp 1667941163
transform 1 0 13064 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1667941163
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_149
timestamp 1667941163
transform 1 0 14812 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_166
timestamp 1667941163
transform 1 0 16376 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_188
timestamp 1667941163
transform 1 0 18400 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1667941163
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_221
timestamp 1667941163
transform 1 0 21436 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_241
timestamp 1667941163
transform 1 0 23276 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_249
timestamp 1667941163
transform 1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_261
timestamp 1667941163
transform 1 0 25116 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_269
timestamp 1667941163
transform 1 0 25852 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_280
timestamp 1667941163
transform 1 0 26864 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_284
timestamp 1667941163
transform 1 0 27232 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_291
timestamp 1667941163
transform 1 0 27876 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1667941163
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1667941163
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_321
timestamp 1667941163
transform 1 0 30636 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_331
timestamp 1667941163
transform 1 0 31556 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_343
timestamp 1667941163
transform 1 0 32660 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_351
timestamp 1667941163
transform 1 0 33396 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_358
timestamp 1667941163
transform 1 0 34040 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_372
timestamp 1667941163
transform 1 0 35328 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_379
timestamp 1667941163
transform 1 0 35972 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_391
timestamp 1667941163
transform 1 0 37076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_403
timestamp 1667941163
transform 1 0 38180 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_407
timestamp 1667941163
transform 1 0 38548 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_414
timestamp 1667941163
transform 1 0 39192 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_421
timestamp 1667941163
transform 1 0 39836 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_429
timestamp 1667941163
transform 1 0 40572 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_436
timestamp 1667941163
transform 1 0 41216 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_448
timestamp 1667941163
transform 1 0 42320 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_458
timestamp 1667941163
transform 1 0 43240 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_466
timestamp 1667941163
transform 1 0 43976 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_474
timestamp 1667941163
transform 1 0 44712 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1667941163
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_489
timestamp 1667941163
transform 1 0 46092 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_514
timestamp 1667941163
transform 1 0 48392 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1667941163
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1667941163
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1667941163
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1667941163
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1667941163
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1667941163
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_93
timestamp 1667941163
transform 1 0 9660 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_101
timestamp 1667941163
transform 1 0 10396 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_109
timestamp 1667941163
transform 1 0 11132 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_131
timestamp 1667941163
transform 1 0 13156 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_144
timestamp 1667941163
transform 1 0 14352 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_155
timestamp 1667941163
transform 1 0 15364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1667941163
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_173
timestamp 1667941163
transform 1 0 17020 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_176
timestamp 1667941163
transform 1 0 17296 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_187
timestamp 1667941163
transform 1 0 18308 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_196
timestamp 1667941163
transform 1 0 19136 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_208
timestamp 1667941163
transform 1 0 20240 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1667941163
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_233
timestamp 1667941163
transform 1 0 22540 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_243
timestamp 1667941163
transform 1 0 23460 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_251
timestamp 1667941163
transform 1 0 24196 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_258
timestamp 1667941163
transform 1 0 24840 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1667941163
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_286
timestamp 1667941163
transform 1 0 27416 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_294
timestamp 1667941163
transform 1 0 28152 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_303
timestamp 1667941163
transform 1 0 28980 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_310
timestamp 1667941163
transform 1 0 29624 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_322
timestamp 1667941163
transform 1 0 30728 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_333
timestamp 1667941163
transform 1 0 31740 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_353
timestamp 1667941163
transform 1 0 33580 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_363
timestamp 1667941163
transform 1 0 34500 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_369
timestamp 1667941163
transform 1 0 35052 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_379
timestamp 1667941163
transform 1 0 35972 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_383
timestamp 1667941163
transform 1 0 36340 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_387
timestamp 1667941163
transform 1 0 36708 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1667941163
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_400
timestamp 1667941163
transform 1 0 37904 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_412
timestamp 1667941163
transform 1 0 39008 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_425
timestamp 1667941163
transform 1 0 40204 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_437
timestamp 1667941163
transform 1 0 41308 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_446
timestamp 1667941163
transform 1 0 42136 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_449
timestamp 1667941163
transform 1 0 42412 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_465
timestamp 1667941163
transform 1 0 43884 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_475
timestamp 1667941163
transform 1 0 44804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_487
timestamp 1667941163
transform 1 0 45908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_502
timestamp 1667941163
transform 1 0 47288 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_505
timestamp 1667941163
transform 1 0 47564 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_510
timestamp 1667941163
transform 1 0 48024 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1667941163
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1667941163
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_37
timestamp 1667941163
transform 1 0 4508 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_43
timestamp 1667941163
transform 1 0 5060 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_55
timestamp 1667941163
transform 1 0 6164 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_67
timestamp 1667941163
transform 1 0 7268 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_79
timestamp 1667941163
transform 1 0 8372 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1667941163
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_91
timestamp 1667941163
transform 1 0 9476 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_95
timestamp 1667941163
transform 1 0 9844 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_120
timestamp 1667941163
transform 1 0 12144 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_132
timestamp 1667941163
transform 1 0 13248 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_156
timestamp 1667941163
transform 1 0 15456 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_163
timestamp 1667941163
transform 1 0 16100 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_175
timestamp 1667941163
transform 1 0 17204 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1667941163
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_205
timestamp 1667941163
transform 1 0 19964 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_217
timestamp 1667941163
transform 1 0 21068 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_235
timestamp 1667941163
transform 1 0 22724 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_241
timestamp 1667941163
transform 1 0 23276 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_247
timestamp 1667941163
transform 1 0 23828 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1667941163
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_259
timestamp 1667941163
transform 1 0 24932 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_271
timestamp 1667941163
transform 1 0 26036 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_283
timestamp 1667941163
transform 1 0 27140 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1667941163
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1667941163
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_337
timestamp 1667941163
transform 1 0 32108 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_346
timestamp 1667941163
transform 1 0 32936 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_354
timestamp 1667941163
transform 1 0 33672 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_361
timestamp 1667941163
transform 1 0 34316 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_374
timestamp 1667941163
transform 1 0 35512 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_394
timestamp 1667941163
transform 1 0 37352 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_404
timestamp 1667941163
transform 1 0 38272 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_416
timestamp 1667941163
transform 1 0 39376 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_421
timestamp 1667941163
transform 1 0 39836 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_429
timestamp 1667941163
transform 1 0 40572 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_441
timestamp 1667941163
transform 1 0 41676 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_462
timestamp 1667941163
transform 1 0 43608 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_471
timestamp 1667941163
transform 1 0 44436 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1667941163
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1667941163
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_489
timestamp 1667941163
transform 1 0 46092 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_514
timestamp 1667941163
transform 1 0 48392 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1667941163
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_27
timestamp 1667941163
transform 1 0 3588 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1667941163
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1667941163
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1667941163
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_93
timestamp 1667941163
transform 1 0 9660 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_102
timestamp 1667941163
transform 1 0 10488 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1667941163
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_121
timestamp 1667941163
transform 1 0 12236 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_126
timestamp 1667941163
transform 1 0 12696 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_138
timestamp 1667941163
transform 1 0 13800 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_159
timestamp 1667941163
transform 1 0 15732 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1667941163
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_181
timestamp 1667941163
transform 1 0 17756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_185
timestamp 1667941163
transform 1 0 18124 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_189
timestamp 1667941163
transform 1 0 18492 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_197
timestamp 1667941163
transform 1 0 19228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_214
timestamp 1667941163
transform 1 0 20792 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1667941163
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_237
timestamp 1667941163
transform 1 0 22908 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_249
timestamp 1667941163
transform 1 0 24012 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_258
timestamp 1667941163
transform 1 0 24840 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_266
timestamp 1667941163
transform 1 0 25576 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1667941163
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_289
timestamp 1667941163
transform 1 0 27692 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_293
timestamp 1667941163
transform 1 0 28060 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_299
timestamp 1667941163
transform 1 0 28612 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_306
timestamp 1667941163
transform 1 0 29256 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_313
timestamp 1667941163
transform 1 0 29900 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_321
timestamp 1667941163
transform 1 0 30636 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1667941163
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1667941163
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_353
timestamp 1667941163
transform 1 0 33580 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_357
timestamp 1667941163
transform 1 0 33948 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_364
timestamp 1667941163
transform 1 0 34592 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_376
timestamp 1667941163
transform 1 0 35696 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_388
timestamp 1667941163
transform 1 0 36800 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_411
timestamp 1667941163
transform 1 0 38916 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_423
timestamp 1667941163
transform 1 0 40020 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_435
timestamp 1667941163
transform 1 0 41124 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1667941163
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1667941163
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1667941163
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1667941163
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_485
timestamp 1667941163
transform 1 0 45724 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_493
timestamp 1667941163
transform 1 0 46460 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_499
timestamp 1667941163
transform 1 0 47012 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1667941163
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_505
timestamp 1667941163
transform 1 0 47564 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_510
timestamp 1667941163
transform 1 0 48024 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_11
timestamp 1667941163
transform 1 0 2116 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1667941163
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1667941163
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_38
timestamp 1667941163
transform 1 0 4600 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_50
timestamp 1667941163
transform 1 0 5704 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_62
timestamp 1667941163
transform 1 0 6808 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_74
timestamp 1667941163
transform 1 0 7912 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1667941163
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_118
timestamp 1667941163
transform 1 0 11960 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_126
timestamp 1667941163
transform 1 0 12696 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1667941163
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_153
timestamp 1667941163
transform 1 0 15180 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_170
timestamp 1667941163
transform 1 0 16744 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_182
timestamp 1667941163
transform 1 0 17848 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1667941163
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_206
timestamp 1667941163
transform 1 0 20056 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_218
timestamp 1667941163
transform 1 0 21160 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_230
timestamp 1667941163
transform 1 0 22264 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_238
timestamp 1667941163
transform 1 0 23000 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1667941163
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_263
timestamp 1667941163
transform 1 0 25300 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_277
timestamp 1667941163
transform 1 0 26588 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_287
timestamp 1667941163
transform 1 0 27508 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_293
timestamp 1667941163
transform 1 0 28060 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_303
timestamp 1667941163
transform 1 0 28980 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1667941163
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1667941163
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_333
timestamp 1667941163
transform 1 0 31740 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_341
timestamp 1667941163
transform 1 0 32476 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_346
timestamp 1667941163
transform 1 0 32936 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_359
timestamp 1667941163
transform 1 0 34132 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_389
timestamp 1667941163
transform 1 0 36892 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_405
timestamp 1667941163
transform 1 0 38364 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_417
timestamp 1667941163
transform 1 0 39468 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_421
timestamp 1667941163
transform 1 0 39836 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_439
timestamp 1667941163
transform 1 0 41492 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_447
timestamp 1667941163
transform 1 0 42228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_454
timestamp 1667941163
transform 1 0 42872 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_463
timestamp 1667941163
transform 1 0 43700 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_467
timestamp 1667941163
transform 1 0 44068 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_473
timestamp 1667941163
transform 1 0 44620 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1667941163
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_489
timestamp 1667941163
transform 1 0 46092 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_514
timestamp 1667941163
transform 1 0 48392 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_9
timestamp 1667941163
transform 1 0 1932 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_31
timestamp 1667941163
transform 1 0 3956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_43
timestamp 1667941163
transform 1 0 5060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1667941163
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1667941163
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_81
timestamp 1667941163
transform 1 0 8556 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_89
timestamp 1667941163
transform 1 0 9292 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_97
timestamp 1667941163
transform 1 0 10028 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_104
timestamp 1667941163
transform 1 0 10672 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_133
timestamp 1667941163
transform 1 0 13340 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_148
timestamp 1667941163
transform 1 0 14720 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_156
timestamp 1667941163
transform 1 0 15456 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1667941163
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_184
timestamp 1667941163
transform 1 0 18032 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_196
timestamp 1667941163
transform 1 0 19136 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_204
timestamp 1667941163
transform 1 0 19872 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1667941163
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_237
timestamp 1667941163
transform 1 0 22908 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_243
timestamp 1667941163
transform 1 0 23460 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_263
timestamp 1667941163
transform 1 0 25300 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1667941163
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_299
timestamp 1667941163
transform 1 0 28612 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_319
timestamp 1667941163
transform 1 0 30452 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_332
timestamp 1667941163
transform 1 0 31648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_343
timestamp 1667941163
transform 1 0 32660 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_350
timestamp 1667941163
transform 1 0 33304 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_370
timestamp 1667941163
transform 1 0 35144 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_382
timestamp 1667941163
transform 1 0 36248 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_390
timestamp 1667941163
transform 1 0 36984 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_417
timestamp 1667941163
transform 1 0 39468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_426
timestamp 1667941163
transform 1 0 40296 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_430
timestamp 1667941163
transform 1 0 40664 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_434
timestamp 1667941163
transform 1 0 41032 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_446
timestamp 1667941163
transform 1 0 42136 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_449
timestamp 1667941163
transform 1 0 42412 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_459
timestamp 1667941163
transform 1 0 43332 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_466
timestamp 1667941163
transform 1 0 43976 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_486
timestamp 1667941163
transform 1 0 45816 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_498
timestamp 1667941163
transform 1 0 46920 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_502
timestamp 1667941163
transform 1 0 47288 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_505
timestamp 1667941163
transform 1 0 47564 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_510
timestamp 1667941163
transform 1 0 48024 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_9
timestamp 1667941163
transform 1 0 1932 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_13
timestamp 1667941163
transform 1 0 2300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_25
timestamp 1667941163
transform 1 0 3404 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1667941163
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1667941163
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1667941163
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1667941163
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1667941163
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1667941163
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_121
timestamp 1667941163
transform 1 0 12236 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_125
timestamp 1667941163
transform 1 0 12604 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1667941163
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_146
timestamp 1667941163
transform 1 0 14536 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_163
timestamp 1667941163
transform 1 0 16100 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_175
timestamp 1667941163
transform 1 0 17204 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1667941163
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_205
timestamp 1667941163
transform 1 0 19964 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_214
timestamp 1667941163
transform 1 0 20792 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_227
timestamp 1667941163
transform 1 0 21988 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_234
timestamp 1667941163
transform 1 0 22632 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_238
timestamp 1667941163
transform 1 0 23000 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_244
timestamp 1667941163
transform 1 0 23552 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_263
timestamp 1667941163
transform 1 0 25300 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_272
timestamp 1667941163
transform 1 0 26128 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1667941163
transform 1 0 26496 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_285
timestamp 1667941163
transform 1 0 27324 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_297
timestamp 1667941163
transform 1 0 28428 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_305
timestamp 1667941163
transform 1 0 29164 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_317
timestamp 1667941163
transform 1 0 30268 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_336
timestamp 1667941163
transform 1 0 32016 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_350
timestamp 1667941163
transform 1 0 33304 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_362
timestamp 1667941163
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_397
timestamp 1667941163
transform 1 0 37628 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_405
timestamp 1667941163
transform 1 0 38364 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_409
timestamp 1667941163
transform 1 0 38732 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_418
timestamp 1667941163
transform 1 0 39560 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_421
timestamp 1667941163
transform 1 0 39836 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_428
timestamp 1667941163
transform 1 0 40480 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_436
timestamp 1667941163
transform 1 0 41216 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_458
timestamp 1667941163
transform 1 0 43240 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_471
timestamp 1667941163
transform 1 0 44436 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1667941163
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_477
timestamp 1667941163
transform 1 0 44988 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_482
timestamp 1667941163
transform 1 0 45448 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_511
timestamp 1667941163
transform 1 0 48116 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_515
timestamp 1667941163
transform 1 0 48484 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1667941163
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1667941163
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1667941163
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1667941163
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1667941163
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1667941163
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_93
timestamp 1667941163
transform 1 0 9660 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_104
timestamp 1667941163
transform 1 0 10672 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_137
timestamp 1667941163
transform 1 0 13708 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_141
timestamp 1667941163
transform 1 0 14076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_158
timestamp 1667941163
transform 1 0 15640 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1667941163
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_177
timestamp 1667941163
transform 1 0 17388 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_190
timestamp 1667941163
transform 1 0 18584 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_202
timestamp 1667941163
transform 1 0 19688 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_206
timestamp 1667941163
transform 1 0 20056 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_216
timestamp 1667941163
transform 1 0 20976 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_234
timestamp 1667941163
transform 1 0 22632 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_242
timestamp 1667941163
transform 1 0 23368 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_250
timestamp 1667941163
transform 1 0 24104 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_257
timestamp 1667941163
transform 1 0 24748 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_269
timestamp 1667941163
transform 1 0 25852 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_277
timestamp 1667941163
transform 1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1667941163
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_321
timestamp 1667941163
transform 1 0 30636 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_329
timestamp 1667941163
transform 1 0 31372 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_334
timestamp 1667941163
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_344
timestamp 1667941163
transform 1 0 32752 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_352
timestamp 1667941163
transform 1 0 33488 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_359
timestamp 1667941163
transform 1 0 34132 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_371
timestamp 1667941163
transform 1 0 35236 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_386
timestamp 1667941163
transform 1 0 36616 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_405
timestamp 1667941163
transform 1 0 38364 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_411
timestamp 1667941163
transform 1 0 38916 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_422
timestamp 1667941163
transform 1 0 39928 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_431
timestamp 1667941163
transform 1 0 40756 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_440
timestamp 1667941163
transform 1 0 41584 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_449
timestamp 1667941163
transform 1 0 42412 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_453
timestamp 1667941163
transform 1 0 42780 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_459
timestamp 1667941163
transform 1 0 43332 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_479
timestamp 1667941163
transform 1 0 45172 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_487
timestamp 1667941163
transform 1 0 45908 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_491
timestamp 1667941163
transform 1 0 46276 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1667941163
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_505
timestamp 1667941163
transform 1 0 47564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_513
timestamp 1667941163
transform 1 0 48300 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1667941163
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1667941163
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1667941163
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1667941163
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1667941163
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_97
timestamp 1667941163
transform 1 0 10028 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_119
timestamp 1667941163
transform 1 0 12052 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_131
timestamp 1667941163
transform 1 0 13156 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1667941163
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_153
timestamp 1667941163
transform 1 0 15180 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_161
timestamp 1667941163
transform 1 0 15916 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_178
timestamp 1667941163
transform 1 0 17480 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_182
timestamp 1667941163
transform 1 0 17848 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_193
timestamp 1667941163
transform 1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_215
timestamp 1667941163
transform 1 0 20884 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_222
timestamp 1667941163
transform 1 0 21528 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_230
timestamp 1667941163
transform 1 0 22264 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_238
timestamp 1667941163
transform 1 0 23000 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1667941163
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_260
timestamp 1667941163
transform 1 0 25024 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_272
timestamp 1667941163
transform 1 0 26128 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_284
timestamp 1667941163
transform 1 0 27232 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_290
timestamp 1667941163
transform 1 0 27784 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_302
timestamp 1667941163
transform 1 0 28888 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_319
timestamp 1667941163
transform 1 0 30452 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_331
timestamp 1667941163
transform 1 0 31556 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_343
timestamp 1667941163
transform 1 0 32660 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_351
timestamp 1667941163
transform 1 0 33396 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_362
timestamp 1667941163
transform 1 0 34408 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_387
timestamp 1667941163
transform 1 0 36708 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_396
timestamp 1667941163
transform 1 0 37536 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_408
timestamp 1667941163
transform 1 0 38640 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_418
timestamp 1667941163
transform 1 0 39560 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_421
timestamp 1667941163
transform 1 0 39836 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_428
timestamp 1667941163
transform 1 0 40480 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_440
timestamp 1667941163
transform 1 0 41584 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_452
timestamp 1667941163
transform 1 0 42688 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_464
timestamp 1667941163
transform 1 0 43792 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_477
timestamp 1667941163
transform 1 0 44988 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_485
timestamp 1667941163
transform 1 0 45724 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_508
timestamp 1667941163
transform 1 0 47840 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1667941163
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1667941163
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1667941163
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1667941163
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1667941163
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1667941163
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1667941163
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1667941163
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1667941163
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1667941163
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_122
timestamp 1667941163
transform 1 0 12328 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_134
timestamp 1667941163
transform 1 0 13432 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_146
timestamp 1667941163
transform 1 0 14536 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_158
timestamp 1667941163
transform 1 0 15640 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1667941163
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_179
timestamp 1667941163
transform 1 0 17572 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_194
timestamp 1667941163
transform 1 0 18952 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_202
timestamp 1667941163
transform 1 0 19688 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_208
timestamp 1667941163
transform 1 0 20240 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1667941163
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_231
timestamp 1667941163
transform 1 0 22356 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_236
timestamp 1667941163
transform 1 0 22816 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_252
timestamp 1667941163
transform 1 0 24288 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_262
timestamp 1667941163
transform 1 0 25208 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_269
timestamp 1667941163
transform 1 0 25852 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_277
timestamp 1667941163
transform 1 0 26588 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_295
timestamp 1667941163
transform 1 0 28244 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_313
timestamp 1667941163
transform 1 0 29900 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_325
timestamp 1667941163
transform 1 0 31004 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_333
timestamp 1667941163
transform 1 0 31740 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_341
timestamp 1667941163
transform 1 0 32476 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_348
timestamp 1667941163
transform 1 0 33120 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_354
timestamp 1667941163
transform 1 0 33672 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_371
timestamp 1667941163
transform 1 0 35236 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_383
timestamp 1667941163
transform 1 0 36340 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_387
timestamp 1667941163
transform 1 0 36708 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1667941163
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_405
timestamp 1667941163
transform 1 0 38364 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_413
timestamp 1667941163
transform 1 0 39100 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_425
timestamp 1667941163
transform 1 0 40204 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_436
timestamp 1667941163
transform 1 0 41216 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1667941163
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1667941163
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1667941163
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_485
timestamp 1667941163
transform 1 0 45724 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_494
timestamp 1667941163
transform 1 0 46552 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_502
timestamp 1667941163
transform 1 0 47288 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_505
timestamp 1667941163
transform 1 0 47564 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_513
timestamp 1667941163
transform 1 0 48300 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1667941163
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1667941163
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1667941163
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1667941163
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1667941163
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1667941163
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1667941163
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1667941163
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1667941163
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1667941163
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_150
timestamp 1667941163
transform 1 0 14904 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_162
timestamp 1667941163
transform 1 0 16008 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_170
timestamp 1667941163
transform 1 0 16744 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_175
timestamp 1667941163
transform 1 0 17204 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_183
timestamp 1667941163
transform 1 0 17940 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_190
timestamp 1667941163
transform 1 0 18584 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_209
timestamp 1667941163
transform 1 0 20332 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_228
timestamp 1667941163
transform 1 0 22080 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_236
timestamp 1667941163
transform 1 0 22816 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_246
timestamp 1667941163
transform 1 0 23736 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_264
timestamp 1667941163
transform 1 0 25392 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_272
timestamp 1667941163
transform 1 0 26128 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_280
timestamp 1667941163
transform 1 0 26864 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_298
timestamp 1667941163
transform 1 0 28520 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_306
timestamp 1667941163
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_320
timestamp 1667941163
transform 1 0 30544 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_332
timestamp 1667941163
transform 1 0 31648 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_338
timestamp 1667941163
transform 1 0 32200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_355
timestamp 1667941163
transform 1 0 33764 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1667941163
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_381
timestamp 1667941163
transform 1 0 36156 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_387
timestamp 1667941163
transform 1 0 36708 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_399
timestamp 1667941163
transform 1 0 37812 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_411
timestamp 1667941163
transform 1 0 38916 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_418
timestamp 1667941163
transform 1 0 39560 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_421
timestamp 1667941163
transform 1 0 39836 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_439
timestamp 1667941163
transform 1 0 41492 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_451
timestamp 1667941163
transform 1 0 42596 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_463
timestamp 1667941163
transform 1 0 43700 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1667941163
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1667941163
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1667941163
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1667941163
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_513
timestamp 1667941163
transform 1 0 48300 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_9
timestamp 1667941163
transform 1 0 1932 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_13
timestamp 1667941163
transform 1 0 2300 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_25
timestamp 1667941163
transform 1 0 3404 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_37
timestamp 1667941163
transform 1 0 4508 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_49
timestamp 1667941163
transform 1 0 5612 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1667941163
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1667941163
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1667941163
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1667941163
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1667941163
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_121
timestamp 1667941163
transform 1 0 12236 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_128
timestamp 1667941163
transform 1 0 12880 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_136
timestamp 1667941163
transform 1 0 13616 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_154
timestamp 1667941163
transform 1 0 15272 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1667941163
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_181
timestamp 1667941163
transform 1 0 17756 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_201
timestamp 1667941163
transform 1 0 19596 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_213
timestamp 1667941163
transform 1 0 20700 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_217
timestamp 1667941163
transform 1 0 21068 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1667941163
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_233
timestamp 1667941163
transform 1 0 22540 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_247
timestamp 1667941163
transform 1 0 23828 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_251
timestamp 1667941163
transform 1 0 24196 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_257
timestamp 1667941163
transform 1 0 24748 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_277
timestamp 1667941163
transform 1 0 26588 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_289
timestamp 1667941163
transform 1 0 27692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_301
timestamp 1667941163
transform 1 0 28796 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_307
timestamp 1667941163
transform 1 0 29348 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_324
timestamp 1667941163
transform 1 0 30912 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_334
timestamp 1667941163
transform 1 0 31832 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_347
timestamp 1667941163
transform 1 0 33028 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_359
timestamp 1667941163
transform 1 0 34132 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_371
timestamp 1667941163
transform 1 0 35236 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_383
timestamp 1667941163
transform 1 0 36340 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_390
timestamp 1667941163
transform 1 0 36984 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_407
timestamp 1667941163
transform 1 0 38548 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_419
timestamp 1667941163
transform 1 0 39652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_431
timestamp 1667941163
transform 1 0 40756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_443
timestamp 1667941163
transform 1 0 41860 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1667941163
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1667941163
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1667941163
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1667941163
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1667941163
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_497
timestamp 1667941163
transform 1 0 46828 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_502
timestamp 1667941163
transform 1 0 47288 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_505
timestamp 1667941163
transform 1 0 47564 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_509
timestamp 1667941163
transform 1 0 47932 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_514
timestamp 1667941163
transform 1 0 48392 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_26
timestamp 1667941163
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1667941163
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1667941163
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1667941163
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1667941163
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_109
timestamp 1667941163
transform 1 0 11132 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_117
timestamp 1667941163
transform 1 0 11868 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_135
timestamp 1667941163
transform 1 0 13524 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1667941163
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_165
timestamp 1667941163
transform 1 0 16284 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_175
timestamp 1667941163
transform 1 0 17204 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_187
timestamp 1667941163
transform 1 0 18308 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1667941163
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_207
timestamp 1667941163
transform 1 0 20148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_219
timestamp 1667941163
transform 1 0 21252 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_225
timestamp 1667941163
transform 1 0 21804 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_237
timestamp 1667941163
transform 1 0 22908 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_247
timestamp 1667941163
transform 1 0 23828 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1667941163
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_261
timestamp 1667941163
transform 1 0 25116 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_269
timestamp 1667941163
transform 1 0 25852 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_281
timestamp 1667941163
transform 1 0 26956 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_293
timestamp 1667941163
transform 1 0 28060 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_305
timestamp 1667941163
transform 1 0 29164 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_319
timestamp 1667941163
transform 1 0 30452 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_325
timestamp 1667941163
transform 1 0 31004 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_342
timestamp 1667941163
transform 1 0 32568 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_354
timestamp 1667941163
transform 1 0 33672 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_362
timestamp 1667941163
transform 1 0 34408 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_371
timestamp 1667941163
transform 1 0 35236 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_393
timestamp 1667941163
transform 1 0 37260 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1667941163
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1667941163
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1667941163
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1667941163
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1667941163
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1667941163
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1667941163
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1667941163
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1667941163
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_489
timestamp 1667941163
transform 1 0 46092 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_514
timestamp 1667941163
transform 1 0 48392 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_11
timestamp 1667941163
transform 1 0 2116 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1667941163
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1667941163
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1667941163
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1667941163
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1667941163
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_61
timestamp 1667941163
transform 1 0 6716 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_68
timestamp 1667941163
transform 1 0 7360 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_75
timestamp 1667941163
transform 1 0 8004 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_87
timestamp 1667941163
transform 1 0 9108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_99
timestamp 1667941163
transform 1 0 10212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1667941163
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_121
timestamp 1667941163
transform 1 0 12236 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_132
timestamp 1667941163
transform 1 0 13248 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_144
timestamp 1667941163
transform 1 0 14352 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1667941163
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_181
timestamp 1667941163
transform 1 0 17756 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_188
timestamp 1667941163
transform 1 0 18400 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_200
timestamp 1667941163
transform 1 0 19504 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_208
timestamp 1667941163
transform 1 0 20240 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_219
timestamp 1667941163
transform 1 0 21252 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1667941163
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_231
timestamp 1667941163
transform 1 0 22356 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_240
timestamp 1667941163
transform 1 0 23184 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_252
timestamp 1667941163
transform 1 0 24288 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_264
timestamp 1667941163
transform 1 0 25392 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_272
timestamp 1667941163
transform 1 0 26128 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_289
timestamp 1667941163
transform 1 0 27692 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_299
timestamp 1667941163
transform 1 0 28612 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_311
timestamp 1667941163
transform 1 0 29716 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_319
timestamp 1667941163
transform 1 0 30452 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_327
timestamp 1667941163
transform 1 0 31188 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_334
timestamp 1667941163
transform 1 0 31832 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_343
timestamp 1667941163
transform 1 0 32660 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_351
timestamp 1667941163
transform 1 0 33396 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_361
timestamp 1667941163
transform 1 0 34316 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_374
timestamp 1667941163
transform 1 0 35512 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_378
timestamp 1667941163
transform 1 0 35880 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_384
timestamp 1667941163
transform 1 0 36432 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_401
timestamp 1667941163
transform 1 0 37996 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_410
timestamp 1667941163
transform 1 0 38824 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_414
timestamp 1667941163
transform 1 0 39192 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_431
timestamp 1667941163
transform 1 0 40756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_443
timestamp 1667941163
transform 1 0 41860 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1667941163
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1667941163
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1667941163
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1667941163
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1667941163
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_497
timestamp 1667941163
transform 1 0 46828 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_502
timestamp 1667941163
transform 1 0 47288 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_505
timestamp 1667941163
transform 1 0 47564 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_510
timestamp 1667941163
transform 1 0 48024 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1667941163
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1667941163
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_61
timestamp 1667941163
transform 1 0 6716 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_81
timestamp 1667941163
transform 1 0 8556 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1667941163
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1667941163
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1667941163
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_133
timestamp 1667941163
transform 1 0 13340 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_137
timestamp 1667941163
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1667941163
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_165
timestamp 1667941163
transform 1 0 16284 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_184
timestamp 1667941163
transform 1 0 18032 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_192
timestamp 1667941163
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_201
timestamp 1667941163
transform 1 0 19596 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_218
timestamp 1667941163
transform 1 0 21160 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_226
timestamp 1667941163
transform 1 0 21896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_243
timestamp 1667941163
transform 1 0 23460 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1667941163
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_261
timestamp 1667941163
transform 1 0 25116 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_269
timestamp 1667941163
transform 1 0 25852 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_279
timestamp 1667941163
transform 1 0 26772 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_291
timestamp 1667941163
transform 1 0 27876 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_297
timestamp 1667941163
transform 1 0 28428 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_306
timestamp 1667941163
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_331
timestamp 1667941163
transform 1 0 31556 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_346
timestamp 1667941163
transform 1 0 32936 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_361
timestamp 1667941163
transform 1 0 34316 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_374
timestamp 1667941163
transform 1 0 35512 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_382
timestamp 1667941163
transform 1 0 36248 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_388
timestamp 1667941163
transform 1 0 36800 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_408
timestamp 1667941163
transform 1 0 38640 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_418
timestamp 1667941163
transform 1 0 39560 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1667941163
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1667941163
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1667941163
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1667941163
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1667941163
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1667941163
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1667941163
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_489
timestamp 1667941163
transform 1 0 46092 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_514
timestamp 1667941163
transform 1 0 48392 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1667941163
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_27
timestamp 1667941163
transform 1 0 3588 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1667941163
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1667941163
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_62
timestamp 1667941163
transform 1 0 6808 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_71
timestamp 1667941163
transform 1 0 7636 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_91
timestamp 1667941163
transform 1 0 9476 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_103
timestamp 1667941163
transform 1 0 10580 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1667941163
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_121
timestamp 1667941163
transform 1 0 12236 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_127
timestamp 1667941163
transform 1 0 12788 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_133
timestamp 1667941163
transform 1 0 13340 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_138
timestamp 1667941163
transform 1 0 13800 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_147
timestamp 1667941163
transform 1 0 14628 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_159
timestamp 1667941163
transform 1 0 15732 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_164
timestamp 1667941163
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_178
timestamp 1667941163
transform 1 0 17480 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_190
timestamp 1667941163
transform 1 0 18584 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_202
timestamp 1667941163
transform 1 0 19688 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_208
timestamp 1667941163
transform 1 0 20240 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_215
timestamp 1667941163
transform 1 0 20884 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1667941163
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_229
timestamp 1667941163
transform 1 0 22172 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_236
timestamp 1667941163
transform 1 0 22816 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_248
timestamp 1667941163
transform 1 0 23920 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_252
timestamp 1667941163
transform 1 0 24288 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_261
timestamp 1667941163
transform 1 0 25116 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_278
timestamp 1667941163
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_299
timestamp 1667941163
transform 1 0 28612 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_319
timestamp 1667941163
transform 1 0 30452 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_325
timestamp 1667941163
transform 1 0 31004 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_334
timestamp 1667941163
transform 1 0 31832 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_365
timestamp 1667941163
transform 1 0 34684 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_374
timestamp 1667941163
transform 1 0 35512 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_381
timestamp 1667941163
transform 1 0 36156 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_389
timestamp 1667941163
transform 1 0 36892 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_403
timestamp 1667941163
transform 1 0 38180 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_413
timestamp 1667941163
transform 1 0 39100 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_425
timestamp 1667941163
transform 1 0 40204 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_437
timestamp 1667941163
transform 1 0 41308 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_445
timestamp 1667941163
transform 1 0 42044 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1667941163
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1667941163
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1667941163
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1667941163
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1667941163
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1667941163
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_505
timestamp 1667941163
transform 1 0 47564 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_510
timestamp 1667941163
transform 1 0 48024 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1667941163
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1667941163
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_43
timestamp 1667941163
transform 1 0 5060 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_53
timestamp 1667941163
transform 1 0 5980 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_60
timestamp 1667941163
transform 1 0 6624 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_72
timestamp 1667941163
transform 1 0 7728 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1667941163
transform 1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1667941163
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_109
timestamp 1667941163
transform 1 0 11132 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_117
timestamp 1667941163
transform 1 0 11868 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_135
timestamp 1667941163
transform 1 0 13524 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1667941163
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_151
timestamp 1667941163
transform 1 0 14996 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_162
timestamp 1667941163
transform 1 0 16008 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_173
timestamp 1667941163
transform 1 0 17020 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_180
timestamp 1667941163
transform 1 0 17664 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_187
timestamp 1667941163
transform 1 0 18308 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1667941163
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_208
timestamp 1667941163
transform 1 0 20240 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_214
timestamp 1667941163
transform 1 0 20792 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_218
timestamp 1667941163
transform 1 0 21160 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_230
timestamp 1667941163
transform 1 0 22264 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_242
timestamp 1667941163
transform 1 0 23368 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_250
timestamp 1667941163
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_271
timestamp 1667941163
transform 1 0 26036 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_279
timestamp 1667941163
transform 1 0 26772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_291
timestamp 1667941163
transform 1 0 27876 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_299
timestamp 1667941163
transform 1 0 28612 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_306
timestamp 1667941163
transform 1 0 29256 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_321
timestamp 1667941163
transform 1 0 30636 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_343
timestamp 1667941163
transform 1 0 32660 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_354
timestamp 1667941163
transform 1 0 33672 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_362
timestamp 1667941163
transform 1 0 34408 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_372
timestamp 1667941163
transform 1 0 35328 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_379
timestamp 1667941163
transform 1 0 35972 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_391
timestamp 1667941163
transform 1 0 37076 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_399
timestamp 1667941163
transform 1 0 37812 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_418
timestamp 1667941163
transform 1 0 39560 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1667941163
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1667941163
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1667941163
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1667941163
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1667941163
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1667941163
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1667941163
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_489
timestamp 1667941163
transform 1 0 46092 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_514
timestamp 1667941163
transform 1 0 48392 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1667941163
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_27
timestamp 1667941163
transform 1 0 3588 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1667941163
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1667941163
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_69
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_79
timestamp 1667941163
transform 1 0 8372 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_90
timestamp 1667941163
transform 1 0 9384 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_102
timestamp 1667941163
transform 1 0 10488 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_110
timestamp 1667941163
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_125
timestamp 1667941163
transform 1 0 12604 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_138
timestamp 1667941163
transform 1 0 13800 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_150
timestamp 1667941163
transform 1 0 14904 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_162
timestamp 1667941163
transform 1 0 16008 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_180
timestamp 1667941163
transform 1 0 17664 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_194
timestamp 1667941163
transform 1 0 18952 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_198
timestamp 1667941163
transform 1 0 19320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_215
timestamp 1667941163
transform 1 0 20884 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1667941163
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_235
timestamp 1667941163
transform 1 0 22724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_247
timestamp 1667941163
transform 1 0 23828 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_259
timestamp 1667941163
transform 1 0 24932 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_271
timestamp 1667941163
transform 1 0 26036 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1667941163
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1667941163
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_317
timestamp 1667941163
transform 1 0 30268 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1667941163
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1667941163
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1667941163
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1667941163
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1667941163
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1667941163
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1667941163
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1667941163
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1667941163
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1667941163
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1667941163
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1667941163
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1667941163
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1667941163
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_497
timestamp 1667941163
transform 1 0 46828 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_502
timestamp 1667941163
transform 1 0 47288 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_505
timestamp 1667941163
transform 1 0 47564 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_510
timestamp 1667941163
transform 1 0 48024 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1667941163
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_45
timestamp 1667941163
transform 1 0 5244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_57
timestamp 1667941163
transform 1 0 6348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_69
timestamp 1667941163
transform 1 0 7452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_81
timestamp 1667941163
transform 1 0 8556 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_90
timestamp 1667941163
transform 1 0 9384 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_102
timestamp 1667941163
transform 1 0 10488 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_114
timestamp 1667941163
transform 1 0 11592 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_126
timestamp 1667941163
transform 1 0 12696 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_137
timestamp 1667941163
transform 1 0 13708 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_160
timestamp 1667941163
transform 1 0 15824 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_170
timestamp 1667941163
transform 1 0 16744 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1667941163
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_209
timestamp 1667941163
transform 1 0 20332 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_219
timestamp 1667941163
transform 1 0 21252 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_227
timestamp 1667941163
transform 1 0 21988 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_232
timestamp 1667941163
transform 1 0 22448 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_240
timestamp 1667941163
transform 1 0 23184 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_48_246
timestamp 1667941163
transform 1 0 23736 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1667941163
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_277
timestamp 1667941163
transform 1 0 26588 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_285
timestamp 1667941163
transform 1 0 27324 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_290
timestamp 1667941163
transform 1 0 27784 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_48_299
timestamp 1667941163
transform 1 0 28612 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1667941163
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_338
timestamp 1667941163
transform 1 0 32200 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_350
timestamp 1667941163
transform 1 0 33304 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_362
timestamp 1667941163
transform 1 0 34408 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_396
timestamp 1667941163
transform 1 0 37536 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_408
timestamp 1667941163
transform 1 0 38640 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1667941163
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1667941163
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1667941163
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1667941163
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1667941163
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1667941163
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1667941163
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_489
timestamp 1667941163
transform 1 0 46092 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_514
timestamp 1667941163
transform 1 0 48392 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1667941163
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1667941163
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_39
timestamp 1667941163
transform 1 0 4692 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_43
timestamp 1667941163
transform 1 0 5060 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_50
timestamp 1667941163
transform 1 0 5704 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_65
timestamp 1667941163
transform 1 0 7084 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_73
timestamp 1667941163
transform 1 0 7820 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_83
timestamp 1667941163
transform 1 0 8740 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_95
timestamp 1667941163
transform 1 0 9844 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_107
timestamp 1667941163
transform 1 0 10948 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1667941163
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1667941163
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1667941163
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_149
timestamp 1667941163
transform 1 0 14812 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_157
timestamp 1667941163
transform 1 0 15548 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_165
timestamp 1667941163
transform 1 0 16284 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_176
timestamp 1667941163
transform 1 0 17296 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_188
timestamp 1667941163
transform 1 0 18400 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_200
timestamp 1667941163
transform 1 0 19504 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_212
timestamp 1667941163
transform 1 0 20608 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1667941163
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_236
timestamp 1667941163
transform 1 0 22816 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_248
timestamp 1667941163
transform 1 0 23920 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_268
timestamp 1667941163
transform 1 0 25760 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_278
timestamp 1667941163
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_287
timestamp 1667941163
transform 1 0 27508 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_297
timestamp 1667941163
transform 1 0 28428 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_310
timestamp 1667941163
transform 1 0 29624 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_318
timestamp 1667941163
transform 1 0 30360 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_327
timestamp 1667941163
transform 1 0 31188 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1667941163
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1667941163
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1667941163
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1667941163
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1667941163
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1667941163
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1667941163
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1667941163
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1667941163
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1667941163
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1667941163
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_497
timestamp 1667941163
transform 1 0 46828 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_502
timestamp 1667941163
transform 1 0 47288 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_505
timestamp 1667941163
transform 1 0 47564 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_510
timestamp 1667941163
transform 1 0 48024 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1667941163
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1667941163
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_51
timestamp 1667941163
transform 1 0 5796 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_79
timestamp 1667941163
transform 1 0 8372 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1667941163
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1667941163
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1667941163
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_121
timestamp 1667941163
transform 1 0 12236 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_131
timestamp 1667941163
transform 1 0 13156 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1667941163
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_153
timestamp 1667941163
transform 1 0 15180 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1667941163
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1667941163
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1667941163
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1667941163
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_216
timestamp 1667941163
transform 1 0 20976 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_229
timestamp 1667941163
transform 1 0 22172 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_242
timestamp 1667941163
transform 1 0 23368 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_246
timestamp 1667941163
transform 1 0 23736 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_250
timestamp 1667941163
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_260
timestamp 1667941163
transform 1 0 25024 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_280
timestamp 1667941163
transform 1 0 26864 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_284
timestamp 1667941163
transform 1 0 27232 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1667941163
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1667941163
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_316
timestamp 1667941163
transform 1 0 30176 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_328
timestamp 1667941163
transform 1 0 31280 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_340
timestamp 1667941163
transform 1 0 32384 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_352
timestamp 1667941163
transform 1 0 33488 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1667941163
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1667941163
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1667941163
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1667941163
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1667941163
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1667941163
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1667941163
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1667941163
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1667941163
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1667941163
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1667941163
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1667941163
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_489
timestamp 1667941163
transform 1 0 46092 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_514
timestamp 1667941163
transform 1 0 48392 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1667941163
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1667941163
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_39
timestamp 1667941163
transform 1 0 4692 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_44
timestamp 1667941163
transform 1 0 5152 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_54
timestamp 1667941163
transform 1 0 6072 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_63
timestamp 1667941163
transform 1 0 6900 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_51_73
timestamp 1667941163
transform 1 0 7820 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_87
timestamp 1667941163
transform 1 0 9108 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_94
timestamp 1667941163
transform 1 0 9752 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_106
timestamp 1667941163
transform 1 0 10856 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_117
timestamp 1667941163
transform 1 0 11868 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_134
timestamp 1667941163
transform 1 0 13432 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_146
timestamp 1667941163
transform 1 0 14536 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_152
timestamp 1667941163
transform 1 0 15088 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_160
timestamp 1667941163
transform 1 0 15824 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_176
timestamp 1667941163
transform 1 0 17296 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_183
timestamp 1667941163
transform 1 0 17940 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_189
timestamp 1667941163
transform 1 0 18492 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_198
timestamp 1667941163
transform 1 0 19320 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_210
timestamp 1667941163
transform 1 0 20424 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1667941163
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_233
timestamp 1667941163
transform 1 0 22540 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_242
timestamp 1667941163
transform 1 0 23368 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_250
timestamp 1667941163
transform 1 0 24104 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_257
timestamp 1667941163
transform 1 0 24748 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_277
timestamp 1667941163
transform 1 0 26588 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_289
timestamp 1667941163
transform 1 0 27692 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_297
timestamp 1667941163
transform 1 0 28428 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_308
timestamp 1667941163
transform 1 0 29440 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_322
timestamp 1667941163
transform 1 0 30728 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_334
timestamp 1667941163
transform 1 0 31832 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1667941163
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1667941163
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1667941163
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1667941163
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1667941163
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1667941163
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1667941163
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1667941163
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1667941163
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1667941163
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1667941163
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1667941163
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1667941163
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_497
timestamp 1667941163
transform 1 0 46828 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_502
timestamp 1667941163
transform 1 0 47288 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_505
timestamp 1667941163
transform 1 0 47564 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_510
timestamp 1667941163
transform 1 0 48024 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1667941163
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1667941163
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_41
timestamp 1667941163
transform 1 0 4876 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_49
timestamp 1667941163
transform 1 0 5612 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_56
timestamp 1667941163
transform 1 0 6256 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_64
timestamp 1667941163
transform 1 0 6992 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 1667941163
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_103
timestamp 1667941163
transform 1 0 10580 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_115
timestamp 1667941163
transform 1 0 11684 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_119
timestamp 1667941163
transform 1 0 12052 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_126
timestamp 1667941163
transform 1 0 12696 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_134
timestamp 1667941163
transform 1 0 13432 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1667941163
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_146
timestamp 1667941163
transform 1 0 14536 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_158
timestamp 1667941163
transform 1 0 15640 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_168
timestamp 1667941163
transform 1 0 16560 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_176
timestamp 1667941163
transform 1 0 17296 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_187
timestamp 1667941163
transform 1 0 18308 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1667941163
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_215
timestamp 1667941163
transform 1 0 20884 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_227
timestamp 1667941163
transform 1 0 21988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_239
timestamp 1667941163
transform 1 0 23092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1667941163
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1667941163
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_289
timestamp 1667941163
transform 1 0 27692 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_297
timestamp 1667941163
transform 1 0 28428 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_302
timestamp 1667941163
transform 1 0 28888 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_317
timestamp 1667941163
transform 1 0 30268 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_326
timestamp 1667941163
transform 1 0 31096 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_334
timestamp 1667941163
transform 1 0 31832 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_341
timestamp 1667941163
transform 1 0 32476 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_353
timestamp 1667941163
transform 1 0 33580 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_361
timestamp 1667941163
transform 1 0 34316 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1667941163
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1667941163
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1667941163
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1667941163
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1667941163
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1667941163
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1667941163
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1667941163
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1667941163
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1667941163
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1667941163
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1667941163
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1667941163
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_513
timestamp 1667941163
transform 1 0 48300 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_27
timestamp 1667941163
transform 1 0 3588 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1667941163
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1667941163
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_53_80
timestamp 1667941163
transform 1 0 8464 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_92
timestamp 1667941163
transform 1 0 9568 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_104
timestamp 1667941163
transform 1 0 10672 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_117
timestamp 1667941163
transform 1 0 11868 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_134
timestamp 1667941163
transform 1 0 13432 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_147
timestamp 1667941163
transform 1 0 14628 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_153
timestamp 1667941163
transform 1 0 15180 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1667941163
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1667941163
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_174
timestamp 1667941163
transform 1 0 17112 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_178
timestamp 1667941163
transform 1 0 17480 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_182
timestamp 1667941163
transform 1 0 17848 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_194
timestamp 1667941163
transform 1 0 18952 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_206
timestamp 1667941163
transform 1 0 20056 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_214
timestamp 1667941163
transform 1 0 20792 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1667941163
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_234
timestamp 1667941163
transform 1 0 22632 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_246
timestamp 1667941163
transform 1 0 23736 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_254
timestamp 1667941163
transform 1 0 24472 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_264
timestamp 1667941163
transform 1 0 25392 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_276
timestamp 1667941163
transform 1 0 26496 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_289
timestamp 1667941163
transform 1 0 27692 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_301
timestamp 1667941163
transform 1 0 28796 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1667941163
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1667941163
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_346
timestamp 1667941163
transform 1 0 32936 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_358
timestamp 1667941163
transform 1 0 34040 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_370
timestamp 1667941163
transform 1 0 35144 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_382
timestamp 1667941163
transform 1 0 36248 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_390
timestamp 1667941163
transform 1 0 36984 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1667941163
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1667941163
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1667941163
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1667941163
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1667941163
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1667941163
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1667941163
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1667941163
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1667941163
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1667941163
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1667941163
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1667941163
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_513
timestamp 1667941163
transform 1 0 48300 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1667941163
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1667941163
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1667941163
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1667941163
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1667941163
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1667941163
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1667941163
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_121
timestamp 1667941163
transform 1 0 12236 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_126
timestamp 1667941163
transform 1 0 12696 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_138
timestamp 1667941163
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_168
timestamp 1667941163
transform 1 0 16560 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_180
timestamp 1667941163
transform 1 0 17664 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_192
timestamp 1667941163
transform 1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_209
timestamp 1667941163
transform 1 0 20332 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_227
timestamp 1667941163
transform 1 0 21988 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_231
timestamp 1667941163
transform 1 0 22356 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_240
timestamp 1667941163
transform 1 0 23184 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_250
timestamp 1667941163
transform 1 0 24104 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_271
timestamp 1667941163
transform 1 0 26036 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_287
timestamp 1667941163
transform 1 0 27508 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_295
timestamp 1667941163
transform 1 0 28244 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_306
timestamp 1667941163
transform 1 0 29256 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_329
timestamp 1667941163
transform 1 0 31372 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_338
timestamp 1667941163
transform 1 0 32200 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_346
timestamp 1667941163
transform 1 0 32936 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_358
timestamp 1667941163
transform 1 0 34040 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1667941163
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1667941163
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1667941163
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1667941163
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1667941163
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1667941163
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1667941163
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1667941163
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1667941163
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1667941163
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1667941163
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1667941163
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1667941163
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_513
timestamp 1667941163
transform 1 0 48300 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_32
timestamp 1667941163
transform 1 0 4048 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_44
timestamp 1667941163
transform 1 0 5152 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1667941163
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1667941163
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1667941163
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1667941163
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1667941163
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1667941163
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1667941163
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_149
timestamp 1667941163
transform 1 0 14812 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_164
timestamp 1667941163
transform 1 0 16192 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_185
timestamp 1667941163
transform 1 0 18124 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_194
timestamp 1667941163
transform 1 0 18952 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_206
timestamp 1667941163
transform 1 0 20056 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_218
timestamp 1667941163
transform 1 0 21160 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_243
timestamp 1667941163
transform 1 0 23460 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_247
timestamp 1667941163
transform 1 0 23828 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_254
timestamp 1667941163
transform 1 0 24472 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_266
timestamp 1667941163
transform 1 0 25576 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_278
timestamp 1667941163
transform 1 0 26680 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_299
timestamp 1667941163
transform 1 0 28612 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_319
timestamp 1667941163
transform 1 0 30452 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_325
timestamp 1667941163
transform 1 0 31004 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_334
timestamp 1667941163
transform 1 0 31832 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_355
timestamp 1667941163
transform 1 0 33764 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_367
timestamp 1667941163
transform 1 0 34868 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_379
timestamp 1667941163
transform 1 0 35972 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1667941163
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1667941163
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1667941163
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1667941163
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1667941163
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1667941163
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1667941163
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1667941163
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1667941163
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1667941163
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1667941163
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1667941163
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_505
timestamp 1667941163
transform 1 0 47564 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_510
timestamp 1667941163
transform 1 0 48024 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_7
timestamp 1667941163
transform 1 0 1748 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_11
timestamp 1667941163
transform 1 0 2116 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_18
timestamp 1667941163
transform 1 0 2760 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_26
timestamp 1667941163
transform 1 0 3496 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1667941163
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1667941163
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1667941163
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1667941163
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1667941163
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_121
timestamp 1667941163
transform 1 0 12236 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_130
timestamp 1667941163
transform 1 0 13064 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_138
timestamp 1667941163
transform 1 0 13800 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_149
timestamp 1667941163
transform 1 0 14812 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_161
timestamp 1667941163
transform 1 0 15916 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_165
timestamp 1667941163
transform 1 0 16284 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_174
timestamp 1667941163
transform 1 0 17112 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_194
timestamp 1667941163
transform 1 0 18952 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_218
timestamp 1667941163
transform 1 0 21160 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_222
timestamp 1667941163
transform 1 0 21528 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_231
timestamp 1667941163
transform 1 0 22356 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_241
timestamp 1667941163
transform 1 0 23276 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_249
timestamp 1667941163
transform 1 0 24012 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_271
timestamp 1667941163
transform 1 0 26036 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_283
timestamp 1667941163
transform 1 0 27140 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_295
timestamp 1667941163
transform 1 0 28244 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_303
timestamp 1667941163
transform 1 0 28980 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1667941163
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_330
timestamp 1667941163
transform 1 0 31464 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_338
timestamp 1667941163
transform 1 0 32200 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_350
timestamp 1667941163
transform 1 0 33304 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_362
timestamp 1667941163
transform 1 0 34408 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1667941163
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1667941163
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1667941163
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1667941163
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1667941163
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1667941163
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1667941163
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1667941163
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1667941163
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1667941163
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1667941163
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_489
timestamp 1667941163
transform 1 0 46092 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_514
timestamp 1667941163
transform 1 0 48392 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1667941163
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1667941163
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1667941163
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1667941163
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1667941163
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1667941163
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1667941163
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1667941163
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1667941163
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_117
timestamp 1667941163
transform 1 0 11868 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_124
timestamp 1667941163
transform 1 0 12512 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_144
timestamp 1667941163
transform 1 0 14352 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_156
timestamp 1667941163
transform 1 0 15456 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_177
timestamp 1667941163
transform 1 0 17388 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_183
timestamp 1667941163
transform 1 0 17940 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_190
timestamp 1667941163
transform 1 0 18584 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_198
timestamp 1667941163
transform 1 0 19320 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_216
timestamp 1667941163
transform 1 0 20976 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1667941163
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1667941163
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1667941163
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1667941163
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_317
timestamp 1667941163
transform 1 0 30268 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_325
timestamp 1667941163
transform 1 0 31004 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_332
timestamp 1667941163
transform 1 0 31648 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_377
timestamp 1667941163
transform 1 0 35788 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_389
timestamp 1667941163
transform 1 0 36892 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1667941163
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1667941163
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1667941163
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1667941163
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1667941163
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1667941163
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1667941163
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1667941163
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1667941163
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1667941163
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_505
timestamp 1667941163
transform 1 0 47564 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_510
timestamp 1667941163
transform 1 0 48024 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1667941163
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1667941163
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1667941163
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1667941163
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_109
timestamp 1667941163
transform 1 0 11132 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_115
timestamp 1667941163
transform 1 0 11684 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_132
timestamp 1667941163
transform 1 0 13248 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_155
timestamp 1667941163
transform 1 0 15364 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_175
timestamp 1667941163
transform 1 0 17204 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_187
timestamp 1667941163
transform 1 0 18308 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1667941163
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_211
timestamp 1667941163
transform 1 0 20516 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_223
timestamp 1667941163
transform 1 0 21620 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_228
timestamp 1667941163
transform 1 0 22080 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_232
timestamp 1667941163
transform 1 0 22448 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_236
timestamp 1667941163
transform 1 0 22816 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_248
timestamp 1667941163
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_277
timestamp 1667941163
transform 1 0 26588 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1667941163
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1667941163
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1667941163
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_320
timestamp 1667941163
transform 1 0 30544 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_331
timestamp 1667941163
transform 1 0 31556 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_343
timestamp 1667941163
transform 1 0 32660 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_355
timestamp 1667941163
transform 1 0 33764 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1667941163
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1667941163
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1667941163
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1667941163
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1667941163
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1667941163
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1667941163
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1667941163
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1667941163
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1667941163
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1667941163
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1667941163
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1667941163
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_513
timestamp 1667941163
transform 1 0 48300 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_9
timestamp 1667941163
transform 1 0 1932 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_21
timestamp 1667941163
transform 1 0 3036 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_33
timestamp 1667941163
transform 1 0 4140 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_45
timestamp 1667941163
transform 1 0 5244 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_53
timestamp 1667941163
transform 1 0 5980 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1667941163
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1667941163
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1667941163
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1667941163
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_145
timestamp 1667941163
transform 1 0 14444 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_149
timestamp 1667941163
transform 1 0 14812 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1667941163
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1667941163
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1667941163
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1667941163
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1667941163
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1667941163
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1667941163
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_234
timestamp 1667941163
transform 1 0 22632 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_243
timestamp 1667941163
transform 1 0 23460 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_251
timestamp 1667941163
transform 1 0 24196 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_256
timestamp 1667941163
transform 1 0 24656 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_265
timestamp 1667941163
transform 1 0 25484 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_275
timestamp 1667941163
transform 1 0 26404 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1667941163
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_299
timestamp 1667941163
transform 1 0 28612 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_309
timestamp 1667941163
transform 1 0 29532 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_333
timestamp 1667941163
transform 1 0 31740 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1667941163
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1667941163
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1667941163
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1667941163
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1667941163
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1667941163
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1667941163
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1667941163
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1667941163
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1667941163
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1667941163
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1667941163
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1667941163
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_505
timestamp 1667941163
transform 1 0 47564 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_513
timestamp 1667941163
transform 1 0 48300 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1667941163
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1667941163
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1667941163
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1667941163
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1667941163
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1667941163
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1667941163
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_133
timestamp 1667941163
transform 1 0 13340 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_138
timestamp 1667941163
transform 1 0 13800 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_145
timestamp 1667941163
transform 1 0 14444 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_149
timestamp 1667941163
transform 1 0 14812 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_60_162
timestamp 1667941163
transform 1 0 16008 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_170
timestamp 1667941163
transform 1 0 16744 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_181
timestamp 1667941163
transform 1 0 17756 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_192
timestamp 1667941163
transform 1 0 18768 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_203
timestamp 1667941163
transform 1 0 19780 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_215
timestamp 1667941163
transform 1 0 20884 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_219
timestamp 1667941163
transform 1 0 21252 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_226
timestamp 1667941163
transform 1 0 21896 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_237
timestamp 1667941163
transform 1 0 22908 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_246
timestamp 1667941163
transform 1 0 23736 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_271
timestamp 1667941163
transform 1 0 26036 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_279
timestamp 1667941163
transform 1 0 26772 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_287
timestamp 1667941163
transform 1 0 27508 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_295
timestamp 1667941163
transform 1 0 28244 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_306
timestamp 1667941163
transform 1 0 29256 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_317
timestamp 1667941163
transform 1 0 30268 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_326
timestamp 1667941163
transform 1 0 31096 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_338
timestamp 1667941163
transform 1 0 32200 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_350
timestamp 1667941163
transform 1 0 33304 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_362
timestamp 1667941163
transform 1 0 34408 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1667941163
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1667941163
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1667941163
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1667941163
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1667941163
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1667941163
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1667941163
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1667941163
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1667941163
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1667941163
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1667941163
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1667941163
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1667941163
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_513
timestamp 1667941163
transform 1 0 48300 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1667941163
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1667941163
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1667941163
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1667941163
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1667941163
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_125
timestamp 1667941163
transform 1 0 12604 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_130
timestamp 1667941163
transform 1 0 13064 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_143
timestamp 1667941163
transform 1 0 14260 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_152
timestamp 1667941163
transform 1 0 15088 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_61_166
timestamp 1667941163
transform 1 0 16376 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_174
timestamp 1667941163
transform 1 0 17112 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_61_184
timestamp 1667941163
transform 1 0 18032 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_200
timestamp 1667941163
transform 1 0 19504 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_209
timestamp 1667941163
transform 1 0 20332 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_221
timestamp 1667941163
transform 1 0 21436 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_243
timestamp 1667941163
transform 1 0 23460 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_255
timestamp 1667941163
transform 1 0 24564 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_265
timestamp 1667941163
transform 1 0 25484 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_274
timestamp 1667941163
transform 1 0 26312 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_293
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_312
timestamp 1667941163
transform 1 0 29808 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_322
timestamp 1667941163
transform 1 0 30728 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_334
timestamp 1667941163
transform 1 0 31832 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_346
timestamp 1667941163
transform 1 0 32936 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_354
timestamp 1667941163
transform 1 0 33672 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_366
timestamp 1667941163
transform 1 0 34776 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_378
timestamp 1667941163
transform 1 0 35880 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_390
timestamp 1667941163
transform 1 0 36984 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1667941163
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1667941163
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1667941163
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1667941163
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1667941163
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1667941163
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1667941163
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1667941163
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1667941163
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1667941163
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_505
timestamp 1667941163
transform 1 0 47564 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_510
timestamp 1667941163
transform 1 0 48024 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1667941163
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1667941163
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1667941163
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1667941163
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1667941163
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1667941163
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1667941163
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1667941163
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_121
timestamp 1667941163
transform 1 0 12236 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_138
timestamp 1667941163
transform 1 0 13800 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_158
timestamp 1667941163
transform 1 0 15640 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_162
timestamp 1667941163
transform 1 0 16008 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_170
timestamp 1667941163
transform 1 0 16744 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_182
timestamp 1667941163
transform 1 0 17848 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_194
timestamp 1667941163
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_202
timestamp 1667941163
transform 1 0 19688 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_206
timestamp 1667941163
transform 1 0 20056 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_213
timestamp 1667941163
transform 1 0 20700 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_225
timestamp 1667941163
transform 1 0 21804 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_232
timestamp 1667941163
transform 1 0 22448 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_244
timestamp 1667941163
transform 1 0 23552 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_258
timestamp 1667941163
transform 1 0 24840 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_269
timestamp 1667941163
transform 1 0 25852 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_276
timestamp 1667941163
transform 1 0 26496 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_283
timestamp 1667941163
transform 1 0 27140 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1667941163
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1667941163
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_340
timestamp 1667941163
transform 1 0 32384 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_352
timestamp 1667941163
transform 1 0 33488 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_359
timestamp 1667941163
transform 1 0 34132 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1667941163
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1667941163
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1667941163
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1667941163
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1667941163
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1667941163
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1667941163
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1667941163
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1667941163
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1667941163
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1667941163
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_489
timestamp 1667941163
transform 1 0 46092 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_514
timestamp 1667941163
transform 1 0 48392 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1667941163
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1667941163
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1667941163
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1667941163
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1667941163
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1667941163
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1667941163
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1667941163
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1667941163
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1667941163
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_125
timestamp 1667941163
transform 1 0 12604 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_131
timestamp 1667941163
transform 1 0 13156 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_141
timestamp 1667941163
transform 1 0 14076 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_153
timestamp 1667941163
transform 1 0 15180 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_166
timestamp 1667941163
transform 1 0 16376 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_181
timestamp 1667941163
transform 1 0 17756 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_203
timestamp 1667941163
transform 1 0 19780 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_215
timestamp 1667941163
transform 1 0 20884 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1667941163
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_236
timestamp 1667941163
transform 1 0 22816 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_248
timestamp 1667941163
transform 1 0 23920 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_254
timestamp 1667941163
transform 1 0 24472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_266
timestamp 1667941163
transform 1 0 25576 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_274
timestamp 1667941163
transform 1 0 26312 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_293
timestamp 1667941163
transform 1 0 28060 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_297
timestamp 1667941163
transform 1 0 28428 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_315
timestamp 1667941163
transform 1 0 30084 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_327
timestamp 1667941163
transform 1 0 31188 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1667941163
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_347
timestamp 1667941163
transform 1 0 33028 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_354
timestamp 1667941163
transform 1 0 33672 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_366
timestamp 1667941163
transform 1 0 34776 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_378
timestamp 1667941163
transform 1 0 35880 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_390
timestamp 1667941163
transform 1 0 36984 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1667941163
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1667941163
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1667941163
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1667941163
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1667941163
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1667941163
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1667941163
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1667941163
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1667941163
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1667941163
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1667941163
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_505
timestamp 1667941163
transform 1 0 47564 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_510
timestamp 1667941163
transform 1 0 48024 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_9
timestamp 1667941163
transform 1 0 1932 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_21
timestamp 1667941163
transform 1 0 3036 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1667941163
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1667941163
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1667941163
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1667941163
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1667941163
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1667941163
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1667941163
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1667941163
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_121
timestamp 1667941163
transform 1 0 12236 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_138
timestamp 1667941163
transform 1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1667941163
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_165
timestamp 1667941163
transform 1 0 16284 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_171
timestamp 1667941163
transform 1 0 16836 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_177
timestamp 1667941163
transform 1 0 17388 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_181
timestamp 1667941163
transform 1 0 17756 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_187
timestamp 1667941163
transform 1 0 18308 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_194
timestamp 1667941163
transform 1 0 18952 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_210
timestamp 1667941163
transform 1 0 20424 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_216
timestamp 1667941163
transform 1 0 20976 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_233
timestamp 1667941163
transform 1 0 22540 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_238
timestamp 1667941163
transform 1 0 23000 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1667941163
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1667941163
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_257
timestamp 1667941163
transform 1 0 24748 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_263
timestamp 1667941163
transform 1 0 25300 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_274
timestamp 1667941163
transform 1 0 26312 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_283
timestamp 1667941163
transform 1 0 27140 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_292
timestamp 1667941163
transform 1 0 27968 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_304
timestamp 1667941163
transform 1 0 29072 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1667941163
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1667941163
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_350
timestamp 1667941163
transform 1 0 33304 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1667941163
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1667941163
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_383
timestamp 1667941163
transform 1 0 36340 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_395
timestamp 1667941163
transform 1 0 37444 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_407
timestamp 1667941163
transform 1 0 38548 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1667941163
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1667941163
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1667941163
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1667941163
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1667941163
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1667941163
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1667941163
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1667941163
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_489
timestamp 1667941163
transform 1 0 46092 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_514
timestamp 1667941163
transform 1 0 48392 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1667941163
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1667941163
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1667941163
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1667941163
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1667941163
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1667941163
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1667941163
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1667941163
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1667941163
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1667941163
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1667941163
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1667941163
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1667941163
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_125
timestamp 1667941163
transform 1 0 12604 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_129
timestamp 1667941163
transform 1 0 12972 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_141
timestamp 1667941163
transform 1 0 14076 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_159
timestamp 1667941163
transform 1 0 15732 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1667941163
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_169
timestamp 1667941163
transform 1 0 16652 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_177
timestamp 1667941163
transform 1 0 17388 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_184
timestamp 1667941163
transform 1 0 18032 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_202
timestamp 1667941163
transform 1 0 19688 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_222
timestamp 1667941163
transform 1 0 21528 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_225
timestamp 1667941163
transform 1 0 21804 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_236
timestamp 1667941163
transform 1 0 22816 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_242
timestamp 1667941163
transform 1 0 23368 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_250
timestamp 1667941163
transform 1 0 24104 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_262
timestamp 1667941163
transform 1 0 25208 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_271
timestamp 1667941163
transform 1 0 26036 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_278
timestamp 1667941163
transform 1 0 26680 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_281
timestamp 1667941163
transform 1 0 26956 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_299
timestamp 1667941163
transform 1 0 28612 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_311
timestamp 1667941163
transform 1 0 29716 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_317
timestamp 1667941163
transform 1 0 30268 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_321
timestamp 1667941163
transform 1 0 30636 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_333
timestamp 1667941163
transform 1 0 31740 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_337
timestamp 1667941163
transform 1 0 32108 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_347
timestamp 1667941163
transform 1 0 33028 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_355
timestamp 1667941163
transform 1 0 33764 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_363
timestamp 1667941163
transform 1 0 34500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_375
timestamp 1667941163
transform 1 0 35604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_387
timestamp 1667941163
transform 1 0 36708 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1667941163
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1667941163
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1667941163
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1667941163
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1667941163
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1667941163
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1667941163
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1667941163
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1667941163
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1667941163
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1667941163
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1667941163
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1667941163
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_505
timestamp 1667941163
transform 1 0 47564 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_510
timestamp 1667941163
transform 1 0 48024 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1667941163
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1667941163
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1667941163
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1667941163
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1667941163
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1667941163
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1667941163
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1667941163
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1667941163
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1667941163
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1667941163
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1667941163
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1667941163
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1667941163
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1667941163
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_66_141
timestamp 1667941163
transform 1 0 14076 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_152
timestamp 1667941163
transform 1 0 15088 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_164
timestamp 1667941163
transform 1 0 16192 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_170
timestamp 1667941163
transform 1 0 16744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_177
timestamp 1667941163
transform 1 0 17388 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1667941163
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1667941163
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_197
timestamp 1667941163
transform 1 0 19228 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_203
timestamp 1667941163
transform 1 0 19780 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_210
timestamp 1667941163
transform 1 0 20424 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_230
timestamp 1667941163
transform 1 0 22264 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_239
timestamp 1667941163
transform 1 0 23092 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_250
timestamp 1667941163
transform 1 0 24104 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_253
timestamp 1667941163
transform 1 0 24380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_66_261
timestamp 1667941163
transform 1 0 25116 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_278
timestamp 1667941163
transform 1 0 26680 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_289
timestamp 1667941163
transform 1 0 27692 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_296
timestamp 1667941163
transform 1 0 28336 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_309
timestamp 1667941163
transform 1 0 29532 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_319
timestamp 1667941163
transform 1 0 30452 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_328
timestamp 1667941163
transform 1 0 31280 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_336
timestamp 1667941163
transform 1 0 32016 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_345
timestamp 1667941163
transform 1 0 32844 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_354
timestamp 1667941163
transform 1 0 33672 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_362
timestamp 1667941163
transform 1 0 34408 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_365
timestamp 1667941163
transform 1 0 34684 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_374
timestamp 1667941163
transform 1 0 35512 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_386
timestamp 1667941163
transform 1 0 36616 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_398
timestamp 1667941163
transform 1 0 37720 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_410
timestamp 1667941163
transform 1 0 38824 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_418
timestamp 1667941163
transform 1 0 39560 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1667941163
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1667941163
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1667941163
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1667941163
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1667941163
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1667941163
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1667941163
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1667941163
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_501
timestamp 1667941163
transform 1 0 47196 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_507
timestamp 1667941163
transform 1 0 47748 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_515
timestamp 1667941163
transform 1 0 48484 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_3
timestamp 1667941163
transform 1 0 1380 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_9
timestamp 1667941163
transform 1 0 1932 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_21
timestamp 1667941163
transform 1 0 3036 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_33
timestamp 1667941163
transform 1 0 4140 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_45
timestamp 1667941163
transform 1 0 5244 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_53
timestamp 1667941163
transform 1 0 5980 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1667941163
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1667941163
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1667941163
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1667941163
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1667941163
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1667941163
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1667941163
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1667941163
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_137
timestamp 1667941163
transform 1 0 13708 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_145
timestamp 1667941163
transform 1 0 14444 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_165
timestamp 1667941163
transform 1 0 16284 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_67_169
timestamp 1667941163
transform 1 0 16652 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_67_191
timestamp 1667941163
transform 1 0 18676 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_67_204
timestamp 1667941163
transform 1 0 19872 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_212
timestamp 1667941163
transform 1 0 20608 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_225
timestamp 1667941163
transform 1 0 21804 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_236
timestamp 1667941163
transform 1 0 22816 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_246
timestamp 1667941163
transform 1 0 23736 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_267
timestamp 1667941163
transform 1 0 25668 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_276
timestamp 1667941163
transform 1 0 26496 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1667941163
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_293
timestamp 1667941163
transform 1 0 28060 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_301
timestamp 1667941163
transform 1 0 28796 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_319
timestamp 1667941163
transform 1 0 30452 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1667941163
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1667941163
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_337
timestamp 1667941163
transform 1 0 32108 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_348
timestamp 1667941163
transform 1 0 33120 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_67_363
timestamp 1667941163
transform 1 0 34500 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1667941163
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1667941163
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1667941163
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1667941163
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1667941163
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1667941163
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1667941163
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1667941163
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1667941163
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1667941163
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1667941163
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1667941163
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1667941163
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1667941163
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_505
timestamp 1667941163
transform 1 0 47564 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_67_510
timestamp 1667941163
transform 1 0 48024 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1667941163
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1667941163
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1667941163
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1667941163
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1667941163
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1667941163
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1667941163
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1667941163
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1667941163
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1667941163
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1667941163
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1667941163
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1667941163
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1667941163
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1667941163
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_141
timestamp 1667941163
transform 1 0 14076 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_159
timestamp 1667941163
transform 1 0 15732 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_171
timestamp 1667941163
transform 1 0 16836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_183
timestamp 1667941163
transform 1 0 17940 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1667941163
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_197
timestamp 1667941163
transform 1 0 19228 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_210
timestamp 1667941163
transform 1 0 20424 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_222
timestamp 1667941163
transform 1 0 21528 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_234
timestamp 1667941163
transform 1 0 22632 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_246
timestamp 1667941163
transform 1 0 23736 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1667941163
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1667941163
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_277
timestamp 1667941163
transform 1 0 26588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_284
timestamp 1667941163
transform 1 0 27232 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_293
timestamp 1667941163
transform 1 0 28060 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_305
timestamp 1667941163
transform 1 0 29164 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_68_309
timestamp 1667941163
transform 1 0 29532 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_315
timestamp 1667941163
transform 1 0 30084 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_325
timestamp 1667941163
transform 1 0 31004 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_332
timestamp 1667941163
transform 1 0 31648 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_341
timestamp 1667941163
transform 1 0 32476 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_68_354
timestamp 1667941163
transform 1 0 33672 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_362
timestamp 1667941163
transform 1 0 34408 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1667941163
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1667941163
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1667941163
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1667941163
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1667941163
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1667941163
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1667941163
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1667941163
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1667941163
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1667941163
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1667941163
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1667941163
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1667941163
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_489
timestamp 1667941163
transform 1 0 46092 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_514
timestamp 1667941163
transform 1 0 48392 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1667941163
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1667941163
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1667941163
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1667941163
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1667941163
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1667941163
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1667941163
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1667941163
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1667941163
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1667941163
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1667941163
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1667941163
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1667941163
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1667941163
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1667941163
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1667941163
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1667941163
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1667941163
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1667941163
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_181
timestamp 1667941163
transform 1 0 17756 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_187
timestamp 1667941163
transform 1 0 18308 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_204
timestamp 1667941163
transform 1 0 19872 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_216
timestamp 1667941163
transform 1 0 20976 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_69_225
timestamp 1667941163
transform 1 0 21804 0 -1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_69_236
timestamp 1667941163
transform 1 0 22816 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_248
timestamp 1667941163
transform 1 0 23920 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_260
timestamp 1667941163
transform 1 0 25024 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_272
timestamp 1667941163
transform 1 0 26128 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_281
timestamp 1667941163
transform 1 0 26956 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_290
timestamp 1667941163
transform 1 0 27784 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_300
timestamp 1667941163
transform 1 0 28704 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_312
timestamp 1667941163
transform 1 0 29808 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_318
timestamp 1667941163
transform 1 0 30360 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_324
timestamp 1667941163
transform 1 0 30912 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_337
timestamp 1667941163
transform 1 0 32108 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_344
timestamp 1667941163
transform 1 0 32752 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_356
timestamp 1667941163
transform 1 0 33856 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_368
timestamp 1667941163
transform 1 0 34960 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_380
timestamp 1667941163
transform 1 0 36064 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1667941163
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1667941163
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1667941163
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1667941163
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1667941163
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1667941163
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1667941163
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1667941163
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1667941163
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1667941163
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_497
timestamp 1667941163
transform 1 0 46828 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_502
timestamp 1667941163
transform 1 0 47288 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_505
timestamp 1667941163
transform 1 0 47564 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_510
timestamp 1667941163
transform 1 0 48024 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_70_3
timestamp 1667941163
transform 1 0 1380 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_11
timestamp 1667941163
transform 1 0 2116 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1667941163
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1667941163
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1667941163
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1667941163
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1667941163
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1667941163
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1667941163
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1667941163
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1667941163
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1667941163
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1667941163
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1667941163
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1667941163
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1667941163
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1667941163
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_153
timestamp 1667941163
transform 1 0 15180 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_70_164
timestamp 1667941163
transform 1 0 16192 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_170
timestamp 1667941163
transform 1 0 16744 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_176
timestamp 1667941163
transform 1 0 17296 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_188
timestamp 1667941163
transform 1 0 18400 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_197
timestamp 1667941163
transform 1 0 19228 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_207
timestamp 1667941163
transform 1 0 20148 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_211
timestamp 1667941163
transform 1 0 20516 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_228
timestamp 1667941163
transform 1 0 22080 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_240
timestamp 1667941163
transform 1 0 23184 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_247
timestamp 1667941163
transform 1 0 23828 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1667941163
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_253
timestamp 1667941163
transform 1 0 24380 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_261
timestamp 1667941163
transform 1 0 25116 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_272
timestamp 1667941163
transform 1 0 26128 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_279
timestamp 1667941163
transform 1 0 26772 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_299
timestamp 1667941163
transform 1 0 28612 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1667941163
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1667941163
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_321
timestamp 1667941163
transform 1 0 30636 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_328
timestamp 1667941163
transform 1 0 31280 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_336
timestamp 1667941163
transform 1 0 32016 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_341
timestamp 1667941163
transform 1 0 32476 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_353
timestamp 1667941163
transform 1 0 33580 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_358
timestamp 1667941163
transform 1 0 34040 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1667941163
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1667941163
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1667941163
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1667941163
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1667941163
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1667941163
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1667941163
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1667941163
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1667941163
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1667941163
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1667941163
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1667941163
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_477
timestamp 1667941163
transform 1 0 44988 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_485
timestamp 1667941163
transform 1 0 45724 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_489
timestamp 1667941163
transform 1 0 46092 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_514
timestamp 1667941163
transform 1 0 48392 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_3
timestamp 1667941163
transform 1 0 1380 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_9
timestamp 1667941163
transform 1 0 1932 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_31
timestamp 1667941163
transform 1 0 3956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_43
timestamp 1667941163
transform 1 0 5060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1667941163
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1667941163
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1667941163
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1667941163
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1667941163
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1667941163
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1667941163
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1667941163
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1667941163
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_137
timestamp 1667941163
transform 1 0 13708 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_157
timestamp 1667941163
transform 1 0 15548 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_166
timestamp 1667941163
transform 1 0 16376 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_169
timestamp 1667941163
transform 1 0 16652 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_177
timestamp 1667941163
transform 1 0 17388 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_189
timestamp 1667941163
transform 1 0 18492 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_71_204
timestamp 1667941163
transform 1 0 19872 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_214
timestamp 1667941163
transform 1 0 20792 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_222
timestamp 1667941163
transform 1 0 21528 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_225
timestamp 1667941163
transform 1 0 21804 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_236
timestamp 1667941163
transform 1 0 22816 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_246
timestamp 1667941163
transform 1 0 23736 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_254
timestamp 1667941163
transform 1 0 24472 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_266
timestamp 1667941163
transform 1 0 25576 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_278
timestamp 1667941163
transform 1 0 26680 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_281
timestamp 1667941163
transform 1 0 26956 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_291
timestamp 1667941163
transform 1 0 27876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_303
timestamp 1667941163
transform 1 0 28980 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_310
timestamp 1667941163
transform 1 0 29624 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_322
timestamp 1667941163
transform 1 0 30728 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_334
timestamp 1667941163
transform 1 0 31832 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_337
timestamp 1667941163
transform 1 0 32108 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_345
timestamp 1667941163
transform 1 0 32844 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_352
timestamp 1667941163
transform 1 0 33488 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_364
timestamp 1667941163
transform 1 0 34592 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_384
timestamp 1667941163
transform 1 0 36432 0 -1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1667941163
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1667941163
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1667941163
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1667941163
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1667941163
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1667941163
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1667941163
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1667941163
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_473
timestamp 1667941163
transform 1 0 44620 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_502
timestamp 1667941163
transform 1 0 47288 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_505
timestamp 1667941163
transform 1 0 47564 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_510
timestamp 1667941163
transform 1 0 48024 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_72_3
timestamp 1667941163
transform 1 0 1380 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_9
timestamp 1667941163
transform 1 0 1932 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_13
timestamp 1667941163
transform 1 0 2300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_25
timestamp 1667941163
transform 1 0 3404 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1667941163
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1667941163
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1667941163
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1667941163
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1667941163
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1667941163
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1667941163
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1667941163
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1667941163
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1667941163
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1667941163
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1667941163
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_141
timestamp 1667941163
transform 1 0 14076 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_147
timestamp 1667941163
transform 1 0 14628 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_151
timestamp 1667941163
transform 1 0 14996 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_155
timestamp 1667941163
transform 1 0 15364 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_172
timestamp 1667941163
transform 1 0 16928 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_181
timestamp 1667941163
transform 1 0 17756 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_193
timestamp 1667941163
transform 1 0 18860 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_72_197
timestamp 1667941163
transform 1 0 19228 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_207
timestamp 1667941163
transform 1 0 20148 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_218
timestamp 1667941163
transform 1 0 21160 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_224
timestamp 1667941163
transform 1 0 21712 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_229
timestamp 1667941163
transform 1 0 22172 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_250
timestamp 1667941163
transform 1 0 24104 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_253
timestamp 1667941163
transform 1 0 24380 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_260
timestamp 1667941163
transform 1 0 25024 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_271
timestamp 1667941163
transform 1 0 26036 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_284
timestamp 1667941163
transform 1 0 27232 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_296
timestamp 1667941163
transform 1 0 28336 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1667941163
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_321
timestamp 1667941163
transform 1 0 30636 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_331
timestamp 1667941163
transform 1 0 31556 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_343
timestamp 1667941163
transform 1 0 32660 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_349
timestamp 1667941163
transform 1 0 33212 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_356
timestamp 1667941163
transform 1 0 33856 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_365
timestamp 1667941163
transform 1 0 34684 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_372
timestamp 1667941163
transform 1 0 35328 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_384
timestamp 1667941163
transform 1 0 36432 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_396
timestamp 1667941163
transform 1 0 37536 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_408
timestamp 1667941163
transform 1 0 38640 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1667941163
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1667941163
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1667941163
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1667941163
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1667941163
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1667941163
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_477
timestamp 1667941163
transform 1 0 44988 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_485
timestamp 1667941163
transform 1 0 45724 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_489
timestamp 1667941163
transform 1 0 46092 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_514
timestamp 1667941163
transform 1 0 48392 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1667941163
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1667941163
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1667941163
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_39
timestamp 1667941163
transform 1 0 4692 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_45
timestamp 1667941163
transform 1 0 5244 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_53
timestamp 1667941163
transform 1 0 5980 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1667941163
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1667941163
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1667941163
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1667941163
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1667941163
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1667941163
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1667941163
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1667941163
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1667941163
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_149
timestamp 1667941163
transform 1 0 14812 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_166
timestamp 1667941163
transform 1 0 16376 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_169
timestamp 1667941163
transform 1 0 16652 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_178
timestamp 1667941163
transform 1 0 17480 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_190
timestamp 1667941163
transform 1 0 18584 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_208
timestamp 1667941163
transform 1 0 20240 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_220
timestamp 1667941163
transform 1 0 21344 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_225
timestamp 1667941163
transform 1 0 21804 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_229
timestamp 1667941163
transform 1 0 22172 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_237
timestamp 1667941163
transform 1 0 22908 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_247
timestamp 1667941163
transform 1 0 23828 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_255
timestamp 1667941163
transform 1 0 24564 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_267
timestamp 1667941163
transform 1 0 25668 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_278
timestamp 1667941163
transform 1 0 26680 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_281
timestamp 1667941163
transform 1 0 26956 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_286
timestamp 1667941163
transform 1 0 27416 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_298
timestamp 1667941163
transform 1 0 28520 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_73_322
timestamp 1667941163
transform 1 0 30728 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_331
timestamp 1667941163
transform 1 0 31556 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1667941163
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_337
timestamp 1667941163
transform 1 0 32108 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_73_346
timestamp 1667941163
transform 1 0 32936 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_352
timestamp 1667941163
transform 1 0 33488 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_358
timestamp 1667941163
transform 1 0 34040 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_370
timestamp 1667941163
transform 1 0 35144 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_377
timestamp 1667941163
transform 1 0 35788 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_389
timestamp 1667941163
transform 1 0 36892 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1667941163
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1667941163
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1667941163
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1667941163
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1667941163
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1667941163
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1667941163
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1667941163
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1667941163
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1667941163
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_497
timestamp 1667941163
transform 1 0 46828 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_502
timestamp 1667941163
transform 1 0 47288 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_505
timestamp 1667941163
transform 1 0 47564 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_73_510
timestamp 1667941163
transform 1 0 48024 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_74_3
timestamp 1667941163
transform 1 0 1380 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_8
timestamp 1667941163
transform 1 0 1840 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_15
timestamp 1667941163
transform 1 0 2484 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_22
timestamp 1667941163
transform 1 0 3128 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1667941163
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_62
timestamp 1667941163
transform 1 0 6808 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_74
timestamp 1667941163
transform 1 0 7912 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_82
timestamp 1667941163
transform 1 0 8648 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1667941163
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1667941163
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1667941163
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1667941163
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1667941163
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1667941163
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1667941163
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1667941163
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_165
timestamp 1667941163
transform 1 0 16284 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_173
timestamp 1667941163
transform 1 0 17020 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_179
timestamp 1667941163
transform 1 0 17572 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_191
timestamp 1667941163
transform 1 0 18676 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1667941163
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_197
timestamp 1667941163
transform 1 0 19228 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_203
timestamp 1667941163
transform 1 0 19780 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_211
timestamp 1667941163
transform 1 0 20516 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_230
timestamp 1667941163
transform 1 0 22264 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_242
timestamp 1667941163
transform 1 0 23368 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_250
timestamp 1667941163
transform 1 0 24104 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_253
timestamp 1667941163
transform 1 0 24380 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_261
timestamp 1667941163
transform 1 0 25116 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_278
timestamp 1667941163
transform 1 0 26680 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_285
timestamp 1667941163
transform 1 0 27324 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_289
timestamp 1667941163
transform 1 0 27692 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_306
timestamp 1667941163
transform 1 0 29256 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_309
timestamp 1667941163
transform 1 0 29532 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_319
timestamp 1667941163
transform 1 0 30452 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_331
timestamp 1667941163
transform 1 0 31556 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_343
timestamp 1667941163
transform 1 0 32660 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_351
timestamp 1667941163
transform 1 0 33396 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_359
timestamp 1667941163
transform 1 0 34132 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1667941163
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_365
timestamp 1667941163
transform 1 0 34684 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_385
timestamp 1667941163
transform 1 0 36524 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_397
timestamp 1667941163
transform 1 0 37628 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_409
timestamp 1667941163
transform 1 0 38732 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_417
timestamp 1667941163
transform 1 0 39468 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1667941163
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1667941163
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1667941163
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1667941163
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1667941163
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1667941163
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1667941163
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_489
timestamp 1667941163
transform 1 0 46092 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_514
timestamp 1667941163
transform 1 0 48392 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_75_3
timestamp 1667941163
transform 1 0 1380 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_9
timestamp 1667941163
transform 1 0 1932 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_16
timestamp 1667941163
transform 1 0 2576 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_24
timestamp 1667941163
transform 1 0 3312 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_38
timestamp 1667941163
transform 1 0 4600 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_50
timestamp 1667941163
transform 1 0 5704 0 -1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1667941163
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1667941163
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1667941163
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1667941163
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1667941163
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1667941163
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1667941163
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1667941163
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1667941163
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1667941163
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1667941163
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1667941163
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_169
timestamp 1667941163
transform 1 0 16652 0 -1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_75_196
timestamp 1667941163
transform 1 0 19136 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_208
timestamp 1667941163
transform 1 0 20240 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_220
timestamp 1667941163
transform 1 0 21344 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1667941163
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1667941163
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1667941163
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_261
timestamp 1667941163
transform 1 0 25116 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_272
timestamp 1667941163
transform 1 0 26128 0 -1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1667941163
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_293
timestamp 1667941163
transform 1 0 28060 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_75_308
timestamp 1667941163
transform 1 0 29440 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_319
timestamp 1667941163
transform 1 0 30452 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_323
timestamp 1667941163
transform 1 0 30820 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1667941163
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1667941163
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_337
timestamp 1667941163
transform 1 0 32108 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_75_345
timestamp 1667941163
transform 1 0 32844 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_351
timestamp 1667941163
transform 1 0 33396 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_359
timestamp 1667941163
transform 1 0 34132 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_367
timestamp 1667941163
transform 1 0 34868 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_379
timestamp 1667941163
transform 1 0 35972 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1667941163
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1667941163
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1667941163
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1667941163
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1667941163
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1667941163
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1667941163
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1667941163
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1667941163
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1667941163
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1667941163
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_497
timestamp 1667941163
transform 1 0 46828 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_502
timestamp 1667941163
transform 1 0 47288 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_505
timestamp 1667941163
transform 1 0 47564 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_75_510
timestamp 1667941163
transform 1 0 48024 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_76_3
timestamp 1667941163
transform 1 0 1380 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_26
timestamp 1667941163
transform 1 0 3496 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_76_29
timestamp 1667941163
transform 1 0 3772 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_35
timestamp 1667941163
transform 1 0 4324 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_48
timestamp 1667941163
transform 1 0 5520 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_60
timestamp 1667941163
transform 1 0 6624 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_72
timestamp 1667941163
transform 1 0 7728 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1667941163
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1667941163
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1667941163
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1667941163
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1667941163
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1667941163
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1667941163
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1667941163
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1667941163
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1667941163
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1667941163
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1667941163
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1667941163
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_230
timestamp 1667941163
transform 1 0 22264 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_242
timestamp 1667941163
transform 1 0 23368 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_250
timestamp 1667941163
transform 1 0 24104 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1667941163
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1667941163
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1667941163
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_289
timestamp 1667941163
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1667941163
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1667941163
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_309
timestamp 1667941163
transform 1 0 29532 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_315
timestamp 1667941163
transform 1 0 30084 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_322
timestamp 1667941163
transform 1 0 30728 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_334
timestamp 1667941163
transform 1 0 31832 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_346
timestamp 1667941163
transform 1 0 32936 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_358
timestamp 1667941163
transform 1 0 34040 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1667941163
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1667941163
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1667941163
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1667941163
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1667941163
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1667941163
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1667941163
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1667941163
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1667941163
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1667941163
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1667941163
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1667941163
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1667941163
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1667941163
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1667941163
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_513
timestamp 1667941163
transform 1 0 48300 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_77_3
timestamp 1667941163
transform 1 0 1380 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_9
timestamp 1667941163
transform 1 0 1932 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_31
timestamp 1667941163
transform 1 0 3956 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1667941163
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1667941163
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1667941163
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1667941163
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1667941163
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_93
timestamp 1667941163
transform 1 0 9660 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_101
timestamp 1667941163
transform 1 0 10396 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1667941163
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1667941163
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1667941163
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1667941163
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1667941163
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1667941163
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1667941163
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1667941163
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1667941163
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1667941163
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1667941163
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_205
timestamp 1667941163
transform 1 0 19964 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_212
timestamp 1667941163
transform 1 0 20608 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1667941163
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1667941163
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1667941163
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1667941163
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1667941163
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1667941163
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1667941163
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1667941163
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1667941163
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1667941163
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1667941163
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1667941163
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1667941163
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1667941163
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1667941163
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1667941163
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1667941163
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1667941163
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1667941163
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1667941163
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1667941163
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1667941163
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1667941163
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1667941163
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1667941163
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1667941163
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1667941163
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1667941163
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1667941163
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1667941163
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_505
timestamp 1667941163
transform 1 0 47564 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_77_510
timestamp 1667941163
transform 1 0 48024 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_78_3
timestamp 1667941163
transform 1 0 1380 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_9
timestamp 1667941163
transform 1 0 1932 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_13
timestamp 1667941163
transform 1 0 2300 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_26
timestamp 1667941163
transform 1 0 3496 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_29
timestamp 1667941163
transform 1 0 3772 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_51
timestamp 1667941163
transform 1 0 5796 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_67
timestamp 1667941163
transform 1 0 7268 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_79
timestamp 1667941163
transform 1 0 8372 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1667941163
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1667941163
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_97
timestamp 1667941163
transform 1 0 10028 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_101
timestamp 1667941163
transform 1 0 10396 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_123
timestamp 1667941163
transform 1 0 12420 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_135
timestamp 1667941163
transform 1 0 13524 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1667941163
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1667941163
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1667941163
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1667941163
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1667941163
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1667941163
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1667941163
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1667941163
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1667941163
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1667941163
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1667941163
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1667941163
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1667941163
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1667941163
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1667941163
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1667941163
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1667941163
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1667941163
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1667941163
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1667941163
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1667941163
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1667941163
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1667941163
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1667941163
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1667941163
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1667941163
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1667941163
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 1667941163
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_401
timestamp 1667941163
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1667941163
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1667941163
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_421
timestamp 1667941163
transform 1 0 39836 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_435
timestamp 1667941163
transform 1 0 41124 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_447
timestamp 1667941163
transform 1 0 42228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_459
timestamp 1667941163
transform 1 0 43332 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_471
timestamp 1667941163
transform 1 0 44436 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1667941163
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1667941163
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_489
timestamp 1667941163
transform 1 0 46092 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_514
timestamp 1667941163
transform 1 0 48392 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_3
timestamp 1667941163
transform 1 0 1380 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_79_32
timestamp 1667941163
transform 1 0 4048 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_79_50
timestamp 1667941163
transform 1 0 5704 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_79_57
timestamp 1667941163
transform 1 0 6348 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_62
timestamp 1667941163
transform 1 0 6808 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1667941163
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1667941163
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_93
timestamp 1667941163
transform 1 0 9660 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_101
timestamp 1667941163
transform 1 0 10396 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1667941163
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1667941163
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1667941163
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1667941163
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_137
timestamp 1667941163
transform 1 0 13708 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_79_146
timestamp 1667941163
transform 1 0 14536 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_152
timestamp 1667941163
transform 1 0 15088 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_156
timestamp 1667941163
transform 1 0 15456 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1667941163
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1667941163
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1667941163
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1667941163
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1667941163
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1667941163
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1667941163
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1667941163
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_249
timestamp 1667941163
transform 1 0 24012 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_260
timestamp 1667941163
transform 1 0 25024 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_267
timestamp 1667941163
transform 1 0 25668 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1667941163
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1667941163
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1667941163
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_305
timestamp 1667941163
transform 1 0 29164 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_314
timestamp 1667941163
transform 1 0 29992 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_326
timestamp 1667941163
transform 1 0 31096 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_334
timestamp 1667941163
transform 1 0 31832 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1667941163
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1667941163
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1667941163
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_376
timestamp 1667941163
transform 1 0 35696 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1667941163
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1667941163
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1667941163
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1667941163
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_417
timestamp 1667941163
transform 1 0 39468 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_421
timestamp 1667941163
transform 1 0 39836 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_425
timestamp 1667941163
transform 1 0 40204 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_440
timestamp 1667941163
transform 1 0 41584 0 -1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1667941163
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1667941163
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_473
timestamp 1667941163
transform 1 0 44620 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_481
timestamp 1667941163
transform 1 0 45356 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_487
timestamp 1667941163
transform 1 0 45908 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_494
timestamp 1667941163
transform 1 0 46552 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_79_501
timestamp 1667941163
transform 1 0 47196 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_505
timestamp 1667941163
transform 1 0 47564 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_79_510
timestamp 1667941163
transform 1 0 48024 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_80_3
timestamp 1667941163
transform 1 0 1380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_26
timestamp 1667941163
transform 1 0 3496 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_29
timestamp 1667941163
transform 1 0 3772 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_40
timestamp 1667941163
transform 1 0 4784 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_44
timestamp 1667941163
transform 1 0 5152 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_66
timestamp 1667941163
transform 1 0 7176 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_73
timestamp 1667941163
transform 1 0 7820 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_81
timestamp 1667941163
transform 1 0 8556 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1667941163
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1667941163
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1667941163
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_121
timestamp 1667941163
transform 1 0 12236 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_126
timestamp 1667941163
transform 1 0 12696 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_134
timestamp 1667941163
transform 1 0 13432 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_138
timestamp 1667941163
transform 1 0 13800 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_80_141
timestamp 1667941163
transform 1 0 14076 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_147
timestamp 1667941163
transform 1 0 14628 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_172
timestamp 1667941163
transform 1 0 16928 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_184
timestamp 1667941163
transform 1 0 18032 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1667941163
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1667941163
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1667941163
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_233
timestamp 1667941163
transform 1 0 22540 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_237
timestamp 1667941163
transform 1 0 22908 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_245
timestamp 1667941163
transform 1 0 23644 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_250
timestamp 1667941163
transform 1 0 24104 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_80_253
timestamp 1667941163
transform 1 0 24380 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_277
timestamp 1667941163
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_289
timestamp 1667941163
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_301
timestamp 1667941163
transform 1 0 28796 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_306
timestamp 1667941163
transform 1 0 29256 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_309
timestamp 1667941163
transform 1 0 29532 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_332
timestamp 1667941163
transform 1 0 31648 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_344
timestamp 1667941163
transform 1 0 32752 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_350
timestamp 1667941163
transform 1 0 33304 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_362
timestamp 1667941163
transform 1 0 34408 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_365
timestamp 1667941163
transform 1 0 34684 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_80_394
timestamp 1667941163
transform 1 0 37352 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_402
timestamp 1667941163
transform 1 0 38088 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_408
timestamp 1667941163
transform 1 0 38640 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_421
timestamp 1667941163
transform 1 0 39836 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_444
timestamp 1667941163
transform 1 0 41952 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_456
timestamp 1667941163
transform 1 0 43056 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_468
timestamp 1667941163
transform 1 0 44160 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_477
timestamp 1667941163
transform 1 0 44988 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_482
timestamp 1667941163
transform 1 0 45448 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_489
timestamp 1667941163
transform 1 0 46092 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_514
timestamp 1667941163
transform 1 0 48392 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_3
timestamp 1667941163
transform 1 0 1380 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_7
timestamp 1667941163
transform 1 0 1748 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_29
timestamp 1667941163
transform 1 0 3772 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_54
timestamp 1667941163
transform 1 0 6072 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_57
timestamp 1667941163
transform 1 0 6348 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_62
timestamp 1667941163
transform 1 0 6808 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_69
timestamp 1667941163
transform 1 0 7452 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_76
timestamp 1667941163
transform 1 0 8096 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_88
timestamp 1667941163
transform 1 0 9200 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_100
timestamp 1667941163
transform 1 0 10304 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_113
timestamp 1667941163
transform 1 0 11500 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_117
timestamp 1667941163
transform 1 0 11868 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_139
timestamp 1667941163
transform 1 0 13892 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_164
timestamp 1667941163
transform 1 0 16192 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_169
timestamp 1667941163
transform 1 0 16652 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_174
timestamp 1667941163
transform 1 0 17112 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_186
timestamp 1667941163
transform 1 0 18216 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_198
timestamp 1667941163
transform 1 0 19320 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_210
timestamp 1667941163
transform 1 0 20424 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_222
timestamp 1667941163
transform 1 0 21528 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_81_225
timestamp 1667941163
transform 1 0 21804 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_231
timestamp 1667941163
transform 1 0 22356 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_253
timestamp 1667941163
transform 1 0 24380 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_278
timestamp 1667941163
transform 1 0 26680 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1667941163
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_293
timestamp 1667941163
transform 1 0 28060 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_299
timestamp 1667941163
transform 1 0 28612 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_324
timestamp 1667941163
transform 1 0 30912 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_337
timestamp 1667941163
transform 1 0 32108 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_81_366
timestamp 1667941163
transform 1 0 34776 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_81_377
timestamp 1667941163
transform 1 0 35788 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_381
timestamp 1667941163
transform 1 0 36156 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1667941163
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1667941163
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_393
timestamp 1667941163
transform 1 0 37260 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_416
timestamp 1667941163
transform 1 0 39376 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1667941163
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1667941163
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_449
timestamp 1667941163
transform 1 0 42412 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_472
timestamp 1667941163
transform 1 0 44528 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_480
timestamp 1667941163
transform 1 0 45264 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_502
timestamp 1667941163
transform 1 0 47288 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_505
timestamp 1667941163
transform 1 0 47564 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_81_510
timestamp 1667941163
transform 1 0 48024 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_82_3
timestamp 1667941163
transform 1 0 1380 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_9
timestamp 1667941163
transform 1 0 1932 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_19
timestamp 1667941163
transform 1 0 2852 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_26
timestamp 1667941163
transform 1 0 3496 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_29
timestamp 1667941163
transform 1 0 3772 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_43
timestamp 1667941163
transform 1 0 5060 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_50
timestamp 1667941163
transform 1 0 5704 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_82_57
timestamp 1667941163
transform 1 0 6348 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_62
timestamp 1667941163
transform 1 0 6808 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_69
timestamp 1667941163
transform 1 0 7452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_81
timestamp 1667941163
transform 1 0 8556 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_82_85
timestamp 1667941163
transform 1 0 8924 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1667941163
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_109
timestamp 1667941163
transform 1 0 11132 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_113
timestamp 1667941163
transform 1 0 11500 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_121
timestamp 1667941163
transform 1 0 12236 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_127
timestamp 1667941163
transform 1 0 12788 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_138
timestamp 1667941163
transform 1 0 13800 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_141
timestamp 1667941163
transform 1 0 14076 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_164
timestamp 1667941163
transform 1 0 16192 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_169
timestamp 1667941163
transform 1 0 16652 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_177
timestamp 1667941163
transform 1 0 17388 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_182
timestamp 1667941163
transform 1 0 17848 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_194
timestamp 1667941163
transform 1 0 18952 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_197
timestamp 1667941163
transform 1 0 19228 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_203
timestamp 1667941163
transform 1 0 19780 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_215
timestamp 1667941163
transform 1 0 20884 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_223
timestamp 1667941163
transform 1 0 21620 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_225
timestamp 1667941163
transform 1 0 21804 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_233
timestamp 1667941163
transform 1 0 22540 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_238
timestamp 1667941163
transform 1 0 23000 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_250
timestamp 1667941163
transform 1 0 24104 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_253
timestamp 1667941163
transform 1 0 24380 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_261
timestamp 1667941163
transform 1 0 25116 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_268
timestamp 1667941163
transform 1 0 25760 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_281
timestamp 1667941163
transform 1 0 26956 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_293
timestamp 1667941163
transform 1 0 28060 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_305
timestamp 1667941163
transform 1 0 29164 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_82_309
timestamp 1667941163
transform 1 0 29532 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_315
timestamp 1667941163
transform 1 0 30084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_327
timestamp 1667941163
transform 1 0 31188 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_335
timestamp 1667941163
transform 1 0 31924 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_337
timestamp 1667941163
transform 1 0 32108 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_343
timestamp 1667941163
transform 1 0 32660 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_350
timestamp 1667941163
transform 1 0 33304 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_362
timestamp 1667941163
transform 1 0 34408 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1667941163
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1667941163
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_389
timestamp 1667941163
transform 1 0 36892 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_393
timestamp 1667941163
transform 1 0 37260 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_408
timestamp 1667941163
transform 1 0 38640 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_421
timestamp 1667941163
transform 1 0 39836 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_426
timestamp 1667941163
transform 1 0 40296 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_434
timestamp 1667941163
transform 1 0 41032 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_439
timestamp 1667941163
transform 1 0 41492 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_447
timestamp 1667941163
transform 1 0 42228 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_449
timestamp 1667941163
transform 1 0 42412 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_455
timestamp 1667941163
transform 1 0 42964 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_467
timestamp 1667941163
transform 1 0 44068 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1667941163
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_477
timestamp 1667941163
transform 1 0 44988 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_502
timestamp 1667941163
transform 1 0 47288 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_82_505
timestamp 1667941163
transform 1 0 47564 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_82_514
timestamp 1667941163
transform 1 0 48392 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1667941163
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1667941163
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1667941163
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1667941163
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1667941163
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1667941163
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1667941163
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1667941163
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1667941163
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1667941163
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1667941163
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1667941163
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1667941163
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1667941163
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1667941163
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1667941163
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1667941163
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1667941163
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1667941163
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1667941163
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1667941163
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1667941163
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1667941163
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1667941163
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1667941163
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1667941163
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1667941163
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1667941163
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1667941163
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1667941163
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1667941163
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1667941163
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1667941163
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1667941163
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1667941163
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1667941163
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1667941163
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1667941163
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1667941163
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1667941163
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1667941163
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1667941163
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1667941163
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1667941163
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1667941163
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1667941163
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1667941163
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1667941163
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1667941163
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1667941163
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1667941163
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1667941163
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1667941163
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1667941163
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1667941163
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1667941163
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1667941163
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1667941163
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1667941163
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1667941163
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1667941163
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1667941163
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1667941163
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1667941163
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1667941163
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1667941163
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1667941163
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1667941163
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1667941163
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1667941163
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1667941163
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1667941163
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1667941163
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1667941163
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1667941163
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1667941163
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1667941163
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1667941163
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1667941163
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1667941163
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1667941163
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1667941163
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1667941163
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1667941163
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1667941163
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1667941163
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1667941163
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1667941163
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1667941163
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1667941163
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1667941163
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1667941163
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1667941163
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1667941163
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1667941163
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1667941163
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1667941163
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1667941163
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1667941163
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1667941163
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1667941163
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1667941163
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1667941163
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1667941163
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1667941163
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1667941163
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1667941163
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1667941163
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1667941163
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1667941163
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1667941163
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1667941163
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1667941163
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1667941163
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1667941163
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1667941163
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1667941163
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1667941163
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1667941163
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1667941163
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1667941163
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1667941163
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1667941163
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1667941163
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1667941163
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1667941163
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1667941163
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1667941163
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1667941163
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1667941163
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1667941163
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1667941163
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1667941163
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1667941163
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1667941163
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1667941163
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1667941163
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1667941163
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1667941163
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1667941163
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1667941163
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1667941163
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1667941163
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1667941163
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1667941163
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1667941163
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1667941163
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1667941163
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1667941163
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1667941163
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1667941163
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1667941163
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1667941163
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1667941163
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1667941163
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1667941163
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1667941163
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1667941163
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1667941163
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1667941163
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1667941163
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1667941163
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1667941163
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1667941163
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1667941163
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1667941163
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1667941163
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1667941163
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1667941163
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1667941163
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1667941163
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1667941163
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1667941163
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1667941163
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1667941163
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1667941163
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1667941163
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1667941163
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1667941163
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1667941163
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1667941163
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1667941163
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1667941163
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1667941163
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1667941163
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1667941163
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1667941163
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1667941163
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1667941163
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1667941163
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1667941163
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1667941163
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1667941163
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1667941163
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1667941163
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1667941163
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1667941163
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1667941163
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1667941163
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1667941163
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1667941163
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1667941163
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1667941163
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1667941163
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1667941163
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1667941163
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1667941163
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1667941163
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1667941163
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1667941163
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1667941163
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1667941163
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1667941163
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1667941163
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1667941163
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1667941163
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1667941163
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1667941163
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1667941163
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1667941163
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1667941163
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1667941163
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1667941163
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1667941163
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1667941163
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1667941163
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1667941163
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1667941163
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1667941163
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1667941163
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1667941163
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1667941163
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1667941163
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1667941163
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1667941163
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1667941163
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1667941163
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1667941163
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1667941163
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1667941163
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1667941163
transform 1 0 42320 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1667941163
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1667941163
transform 1 0 47472 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_6  _0951_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2024 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  _0952_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  _0953_
timestamp 1667941163
transform 1 0 5428 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0954_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2760 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0955_
timestamp 1667941163
transform 1 0 47748 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0956_
timestamp 1667941163
transform 1 0 2116 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0957_
timestamp 1667941163
transform 1 0 2760 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0958_
timestamp 1667941163
transform 1 0 39928 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0959_
timestamp 1667941163
transform 1 0 47012 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0960_
timestamp 1667941163
transform 1 0 2208 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0961_
timestamp 1667941163
transform 1 0 47748 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0962_
timestamp 1667941163
transform 1 0 45816 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0963_
timestamp 1667941163
transform 1 0 47748 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0964_
timestamp 1667941163
transform 1 0 40020 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0965_
timestamp 1667941163
transform 1 0 10396 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0966_
timestamp 1667941163
transform 1 0 39928 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0967_
timestamp 1667941163
transform 1 0 10396 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0968_
timestamp 1667941163
transform 1 0 32476 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0969_
timestamp 1667941163
transform 1 0 40756 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0970_
timestamp 1667941163
transform 1 0 28244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1667941163
transform 1 0 36248 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0972_
timestamp 1667941163
transform 1 0 10212 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1667941163
transform 1 0 38364 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0974_
timestamp 1667941163
transform 1 0 16100 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0975_
timestamp 1667941163
transform 1 0 3496 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0976_
timestamp 1667941163
transform 1 0 47748 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0977_
timestamp 1667941163
transform 1 0 2760 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0978_
timestamp 1667941163
transform 1 0 2760 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0979_
timestamp 1667941163
transform 1 0 6532 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0980_
timestamp 1667941163
transform 1 0 47748 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0981_
timestamp 1667941163
transform 1 0 47748 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0982_
timestamp 1667941163
transform 1 0 47748 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0983_
timestamp 1667941163
transform 1 0 15180 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0984_
timestamp 1667941163
transform 1 0 47748 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp 1667941163
transform 1 0 39008 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _0986_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3956 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _0987_
timestamp 1667941163
transform 1 0 41308 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0988_
timestamp 1667941163
transform 1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0989_
timestamp 1667941163
transform 1 0 43792 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0990_
timestamp 1667941163
transform 1 0 2484 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1667941163
transform 1 0 47748 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0992_
timestamp 1667941163
transform 1 0 12420 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0993_
timestamp 1667941163
transform 1 0 1932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0994_
timestamp 1667941163
transform 1 0 10488 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0995_
timestamp 1667941163
transform 1 0 2484 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0996_
timestamp 1667941163
transform 1 0 47748 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0997_
timestamp 1667941163
transform 1 0 6164 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0998_
timestamp 1667941163
transform 1 0 47012 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0999_
timestamp 1667941163
transform 1 0 47012 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1000_
timestamp 1667941163
transform 1 0 2760 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1001_
timestamp 1667941163
transform 1 0 13524 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1002_
timestamp 1667941163
transform 1 0 46368 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1003_
timestamp 1667941163
transform 1 0 12972 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1004_
timestamp 1667941163
transform 1 0 35420 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1005_
timestamp 1667941163
transform 1 0 14352 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1006_
timestamp 1667941163
transform 1 0 47012 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1007_
timestamp 1667941163
transform 1 0 7544 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1008_
timestamp 1667941163
transform 1 0 4600 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1009_
timestamp 1667941163
transform 1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1010_
timestamp 1667941163
transform 1 0 24748 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1011_
timestamp 1667941163
transform 1 0 25392 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1012_
timestamp 1667941163
transform 1 0 48116 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1013_
timestamp 1667941163
transform 1 0 47748 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1014_
timestamp 1667941163
transform 1 0 28980 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1015_
timestamp 1667941163
transform 1 0 41584 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1016_
timestamp 1667941163
transform 1 0 47748 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1017_
timestamp 1667941163
transform 1 0 6532 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1018_
timestamp 1667941163
transform 1 0 41400 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1019_
timestamp 1667941163
transform 1 0 3956 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1020_
timestamp 1667941163
transform 1 0 2208 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1021_
timestamp 1667941163
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1022_
timestamp 1667941163
transform 1 0 8280 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1023_
timestamp 1667941163
transform 1 0 10488 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1024_
timestamp 1667941163
transform 1 0 2208 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1025_
timestamp 1667941163
transform 1 0 2208 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1026_
timestamp 1667941163
transform 1 0 19320 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1027_
timestamp 1667941163
transform 1 0 2208 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1028_
timestamp 1667941163
transform 1 0 2208 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1667941163
transform 1 0 2208 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1030_
timestamp 1667941163
transform 1 0 4416 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1031_
timestamp 1667941163
transform 1 0 45172 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1032_
timestamp 1667941163
transform 1 0 3220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1033_
timestamp 1667941163
transform 1 0 46736 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1034_
timestamp 1667941163
transform 1 0 9568 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1035_
timestamp 1667941163
transform 1 0 46276 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1036_
timestamp 1667941163
transform 1 0 46000 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1037_
timestamp 1667941163
transform 1 0 46736 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1038_
timestamp 1667941163
transform 1 0 22080 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1039_
timestamp 1667941163
transform 1 0 17296 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1040_
timestamp 1667941163
transform 1 0 4968 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1041_
timestamp 1667941163
transform 1 0 2392 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1042_
timestamp 1667941163
transform 1 0 20332 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1043_
timestamp 1667941163
transform 1 0 3956 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1044_
timestamp 1667941163
transform 1 0 47012 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1045_
timestamp 1667941163
transform 1 0 47748 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1046_
timestamp 1667941163
transform 1 0 5428 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1047_
timestamp 1667941163
transform 1 0 47012 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1048_
timestamp 1667941163
transform 1 0 3956 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1049_
timestamp 1667941163
transform 1 0 47748 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1050_
timestamp 1667941163
transform 1 0 29716 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1051_
timestamp 1667941163
transform 1 0 12972 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1052_
timestamp 1667941163
transform 1 0 3956 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1053_
timestamp 1667941163
transform 1 0 47012 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1054_
timestamp 1667941163
transform 1 0 2300 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1055_
timestamp 1667941163
transform 1 0 47012 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1056_
timestamp 1667941163
transform 1 0 7176 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1057_
timestamp 1667941163
transform 1 0 47472 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1058_
timestamp 1667941163
transform 1 0 44712 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1059_
timestamp 1667941163
transform 1 0 2300 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1060_
timestamp 1667941163
transform 1 0 47748 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1061_
timestamp 1667941163
transform 1 0 22632 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1062_
timestamp 1667941163
transform 1 0 33028 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1063_
timestamp 1667941163
transform 1 0 6624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1064_
timestamp 1667941163
transform 1 0 45816 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1065_
timestamp 1667941163
transform 1 0 4692 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1066_
timestamp 1667941163
transform 1 0 46920 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1067_
timestamp 1667941163
transform 1 0 4784 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1068_
timestamp 1667941163
transform 1 0 18400 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1069_
timestamp 1667941163
transform 1 0 25300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1070_
timestamp 1667941163
transform 1 0 47748 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1071_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 12420 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1072_
timestamp 1667941163
transform 1 0 12972 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1073_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 13248 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1074_
timestamp 1667941163
transform 1 0 14720 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1075_
timestamp 1667941163
transform 1 0 13708 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1076_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11776 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1077_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14904 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1078_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 15180 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1079_
timestamp 1667941163
transform 1 0 15548 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1080_
timestamp 1667941163
transform 1 0 12420 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1081_
timestamp 1667941163
transform 1 0 12788 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1082_
timestamp 1667941163
transform 1 0 12328 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1083_
timestamp 1667941163
transform 1 0 13892 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1084_
timestamp 1667941163
transform 1 0 14260 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1085_
timestamp 1667941163
transform 1 0 15272 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1086_
timestamp 1667941163
transform 1 0 15824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1087_
timestamp 1667941163
transform 1 0 15548 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1088_
timestamp 1667941163
transform 1 0 14996 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1089_
timestamp 1667941163
transform 1 0 14536 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1090_
timestamp 1667941163
transform 1 0 13524 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1091_
timestamp 1667941163
transform 1 0 14352 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1092_
timestamp 1667941163
transform 1 0 12880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1093_
timestamp 1667941163
transform 1 0 12696 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1094_
timestamp 1667941163
transform 1 0 12052 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1095_
timestamp 1667941163
transform 1 0 12236 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1096_
timestamp 1667941163
transform 1 0 11684 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1097_
timestamp 1667941163
transform 1 0 8740 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1098_
timestamp 1667941163
transform 1 0 9844 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1099_
timestamp 1667941163
transform 1 0 9384 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1100_
timestamp 1667941163
transform 1 0 9752 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1101_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 40204 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1102_
timestamp 1667941163
transform 1 0 40572 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _1103_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 25668 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1104_
timestamp 1667941163
transform 1 0 39376 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1105_
timestamp 1667941163
transform 1 0 39284 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1106_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 25668 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1107_
timestamp 1667941163
transform 1 0 26036 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _1108_
timestamp 1667941163
transform 1 0 40296 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1109_
timestamp 1667941163
transform 1 0 38456 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1110_
timestamp 1667941163
transform 1 0 38456 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _1111_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 40296 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1112_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 39744 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1113_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 39284 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1114_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 40020 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1115_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 39560 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1116_
timestamp 1667941163
transform 1 0 40020 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1117_
timestamp 1667941163
transform 1 0 25852 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1118_
timestamp 1667941163
transform 1 0 26036 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1119_
timestamp 1667941163
transform 1 0 39100 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1120_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 38916 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1121_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 36708 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1122_
timestamp 1667941163
transform 1 0 36340 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1123_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 36248 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1124_
timestamp 1667941163
transform 1 0 36432 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1125_
timestamp 1667941163
transform 1 0 37076 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1126_
timestamp 1667941163
transform 1 0 39284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1127_
timestamp 1667941163
transform 1 0 37904 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1128_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 36156 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1129_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 35788 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1130_
timestamp 1667941163
transform 1 0 35052 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1131_
timestamp 1667941163
transform 1 0 35880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1132_
timestamp 1667941163
transform 1 0 35696 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1133_
timestamp 1667941163
transform 1 0 35788 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1134_
timestamp 1667941163
transform 1 0 34868 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1135_
timestamp 1667941163
transform 1 0 34684 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1136_
timestamp 1667941163
transform 1 0 33488 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1137_
timestamp 1667941163
transform 1 0 33396 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1138_
timestamp 1667941163
transform 1 0 31556 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1139_
timestamp 1667941163
transform 1 0 32292 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1140_
timestamp 1667941163
transform 1 0 32660 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1141_
timestamp 1667941163
transform 1 0 34868 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1142_
timestamp 1667941163
transform 1 0 35972 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a311oi_4  _1143_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 35328 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2_1  _1144_
timestamp 1667941163
transform 1 0 33672 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1145_
timestamp 1667941163
transform 1 0 33672 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1146_
timestamp 1667941163
transform 1 0 32752 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1147_
timestamp 1667941163
transform 1 0 30820 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1148_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 33764 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1149_
timestamp 1667941163
transform 1 0 37444 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1150_
timestamp 1667941163
transform 1 0 36432 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1151_
timestamp 1667941163
transform 1 0 34868 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1152_
timestamp 1667941163
transform 1 0 34868 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1153_
timestamp 1667941163
transform 1 0 32476 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1154_
timestamp 1667941163
transform 1 0 35144 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1155_
timestamp 1667941163
transform 1 0 35696 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1156_
timestamp 1667941163
transform 1 0 36340 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1157_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 36432 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1158_
timestamp 1667941163
transform 1 0 36708 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _1159_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37444 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1160_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 36616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1161_
timestamp 1667941163
transform 1 0 42596 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1162_
timestamp 1667941163
transform 1 0 34868 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1163_
timestamp 1667941163
transform 1 0 35696 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1164_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 35328 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1165_
timestamp 1667941163
transform 1 0 34040 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1166_
timestamp 1667941163
transform 1 0 34684 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1167_
timestamp 1667941163
transform 1 0 35512 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1168_
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1169_
timestamp 1667941163
transform 1 0 34868 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1170_
timestamp 1667941163
transform 1 0 34592 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_1  _1171_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 33672 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1172_
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1173_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 33672 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1174_
timestamp 1667941163
transform 1 0 35420 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1175_
timestamp 1667941163
transform 1 0 33856 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1176_
timestamp 1667941163
transform 1 0 33764 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1177_
timestamp 1667941163
transform 1 0 28980 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1178_
timestamp 1667941163
transform 1 0 28152 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1179_
timestamp 1667941163
transform 1 0 29624 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1180_
timestamp 1667941163
transform 1 0 29348 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1181_
timestamp 1667941163
transform 1 0 28520 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1182_
timestamp 1667941163
transform 1 0 28244 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1183_
timestamp 1667941163
transform 1 0 28152 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1184_
timestamp 1667941163
transform 1 0 28060 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1185_
timestamp 1667941163
transform 1 0 27140 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1186_
timestamp 1667941163
transform 1 0 26404 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1187_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 28244 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1188_
timestamp 1667941163
transform 1 0 28796 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1189_
timestamp 1667941163
transform 1 0 27784 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1190_
timestamp 1667941163
transform 1 0 26036 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1191_
timestamp 1667941163
transform 1 0 26312 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1192_
timestamp 1667941163
transform 1 0 27140 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1193_
timestamp 1667941163
transform 1 0 26864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1194_
timestamp 1667941163
transform 1 0 27324 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1195_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 27508 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1196_
timestamp 1667941163
transform 1 0 27508 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1197_
timestamp 1667941163
transform 1 0 28520 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1198_
timestamp 1667941163
transform 1 0 28520 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1199_
timestamp 1667941163
transform 1 0 24380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1200_
timestamp 1667941163
transform 1 0 25392 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1201_
timestamp 1667941163
transform 1 0 26220 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1202_
timestamp 1667941163
transform 1 0 26864 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1203_
timestamp 1667941163
transform 1 0 25668 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1204_
timestamp 1667941163
transform 1 0 24564 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1205_
timestamp 1667941163
transform 1 0 24840 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1206_
timestamp 1667941163
transform 1 0 23460 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1207_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 27784 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1208_
timestamp 1667941163
transform 1 0 28520 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1209_
timestamp 1667941163
transform 1 0 32752 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1210_
timestamp 1667941163
transform 1 0 25024 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1211_
timestamp 1667941163
transform 1 0 27232 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1212_
timestamp 1667941163
transform 1 0 27508 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1213_
timestamp 1667941163
transform 1 0 28152 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1214_
timestamp 1667941163
transform 1 0 28980 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1215_
timestamp 1667941163
transform 1 0 29716 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1216_
timestamp 1667941163
transform 1 0 29532 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1217_
timestamp 1667941163
transform 1 0 28612 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1218_
timestamp 1667941163
transform 1 0 27140 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1219_
timestamp 1667941163
transform 1 0 28888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1220_
timestamp 1667941163
transform 1 0 27968 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1221_
timestamp 1667941163
transform 1 0 27876 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1222_
timestamp 1667941163
transform 1 0 29532 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1223_
timestamp 1667941163
transform 1 0 28520 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1224_
timestamp 1667941163
transform 1 0 26128 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1225_
timestamp 1667941163
transform 1 0 27140 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1226_
timestamp 1667941163
transform 1 0 40664 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1227_
timestamp 1667941163
transform 1 0 28796 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1228_
timestamp 1667941163
transform 1 0 31372 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1229_
timestamp 1667941163
transform 1 0 30728 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1230_
timestamp 1667941163
transform 1 0 31924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1231_
timestamp 1667941163
transform 1 0 30728 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1232_
timestamp 1667941163
transform 1 0 31372 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1233_
timestamp 1667941163
transform 1 0 31464 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1234_
timestamp 1667941163
transform 1 0 32292 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1235_
timestamp 1667941163
transform 1 0 33120 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1236_
timestamp 1667941163
transform 1 0 33764 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1237_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 33764 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1238_
timestamp 1667941163
transform 1 0 31464 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1239_
timestamp 1667941163
transform 1 0 32752 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1240_
timestamp 1667941163
transform 1 0 33764 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1241_
timestamp 1667941163
transform 1 0 33304 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1242_
timestamp 1667941163
transform 1 0 33764 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1243_
timestamp 1667941163
transform 1 0 21252 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1244_
timestamp 1667941163
transform 1 0 23828 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1245_
timestamp 1667941163
transform 1 0 24564 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1246_
timestamp 1667941163
transform 1 0 23460 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1247_
timestamp 1667941163
transform 1 0 20884 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1248_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 20332 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1249_
timestamp 1667941163
transform 1 0 13524 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1250_
timestamp 1667941163
transform 1 0 16836 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1251_
timestamp 1667941163
transform 1 0 14260 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1252_
timestamp 1667941163
transform 1 0 15088 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1253_
timestamp 1667941163
transform 1 0 21344 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1254_
timestamp 1667941163
transform 1 0 18492 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1255_
timestamp 1667941163
transform 1 0 28336 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1256_
timestamp 1667941163
transform 1 0 29716 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1257_
timestamp 1667941163
transform 1 0 28612 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1258_
timestamp 1667941163
transform 1 0 32292 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1259_
timestamp 1667941163
transform 1 0 31188 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1260_
timestamp 1667941163
transform 1 0 32016 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1261_
timestamp 1667941163
transform 1 0 32568 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1262_
timestamp 1667941163
transform 1 0 27876 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1263_
timestamp 1667941163
transform 1 0 13524 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1264_
timestamp 1667941163
transform 1 0 14628 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1265_
timestamp 1667941163
transform 1 0 16836 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1266_
timestamp 1667941163
transform 1 0 19412 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1267_
timestamp 1667941163
transform 1 0 14536 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1268_
timestamp 1667941163
transform 1 0 14536 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1269_
timestamp 1667941163
transform 1 0 15364 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _1270_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16928 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1271_
timestamp 1667941163
transform 1 0 13432 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1272_
timestamp 1667941163
transform 1 0 17388 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1273_
timestamp 1667941163
transform 1 0 14812 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1274_
timestamp 1667941163
transform 1 0 13432 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1275_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 15272 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1276_
timestamp 1667941163
transform 1 0 17204 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1277_
timestamp 1667941163
transform 1 0 15916 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1278_
timestamp 1667941163
transform 1 0 15364 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1279_
timestamp 1667941163
transform 1 0 16836 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1280_
timestamp 1667941163
transform 1 0 16284 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1281_
timestamp 1667941163
transform 1 0 15180 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1282_
timestamp 1667941163
transform 1 0 15456 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1283_
timestamp 1667941163
transform 1 0 22172 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1284_
timestamp 1667941163
transform 1 0 23276 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1285_
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1286_
timestamp 1667941163
transform 1 0 22080 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1287_
timestamp 1667941163
transform 1 0 27508 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1288_
timestamp 1667941163
transform 1 0 28060 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1289_
timestamp 1667941163
transform 1 0 26220 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1290_
timestamp 1667941163
transform 1 0 25852 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1291_
timestamp 1667941163
transform 1 0 26864 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1292_
timestamp 1667941163
transform 1 0 26036 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1293_
timestamp 1667941163
transform 1 0 22540 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1294_
timestamp 1667941163
transform 1 0 23368 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1295_
timestamp 1667941163
transform 1 0 23184 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1296_
timestamp 1667941163
transform 1 0 24564 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1297_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 23460 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1298_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 25300 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_4  _1299_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24104 0 -1 39168
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_4  _1300_
timestamp 1667941163
transform 1 0 30820 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1301_
timestamp 1667941163
transform 1 0 33580 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1302_
timestamp 1667941163
transform 1 0 33580 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1303_
timestamp 1667941163
transform 1 0 35512 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1304_
timestamp 1667941163
transform 1 0 33028 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1305_
timestamp 1667941163
transform 1 0 25668 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1306_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 26404 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1307_
timestamp 1667941163
transform 1 0 17848 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1308_
timestamp 1667941163
transform 1 0 18676 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1309_
timestamp 1667941163
transform 1 0 19872 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1310_
timestamp 1667941163
transform 1 0 24564 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1311_
timestamp 1667941163
transform 1 0 33672 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1312_
timestamp 1667941163
transform 1 0 19136 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _1313_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 33856 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1314_
timestamp 1667941163
transform 1 0 33488 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1315_
timestamp 1667941163
transform 1 0 34868 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1316_
timestamp 1667941163
transform 1 0 34500 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1317_
timestamp 1667941163
transform 1 0 34408 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1318_
timestamp 1667941163
transform 1 0 32936 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1319_
timestamp 1667941163
transform 1 0 28152 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1320_
timestamp 1667941163
transform 1 0 33764 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1321_
timestamp 1667941163
transform 1 0 30452 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1322_
timestamp 1667941163
transform 1 0 30912 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1323_
timestamp 1667941163
transform 1 0 31096 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1324_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 31924 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _1325_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 32292 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1326_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 30176 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1327_
timestamp 1667941163
transform 1 0 30820 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1328_
timestamp 1667941163
transform 1 0 28796 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1329_
timestamp 1667941163
transform 1 0 29716 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1330_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 20240 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1331_
timestamp 1667941163
transform 1 0 29808 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1332_
timestamp 1667941163
transform 1 0 29716 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1333_
timestamp 1667941163
transform 1 0 30820 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1334_
timestamp 1667941163
transform 1 0 29808 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1335_
timestamp 1667941163
transform 1 0 30360 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1336_
timestamp 1667941163
transform 1 0 33028 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _1337_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 32292 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _1338_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 30728 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1339_
timestamp 1667941163
transform 1 0 30912 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1340_
timestamp 1667941163
transform 1 0 30452 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1341_
timestamp 1667941163
transform 1 0 31372 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1342_
timestamp 1667941163
transform 1 0 29716 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1343_
timestamp 1667941163
transform 1 0 33028 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1344_
timestamp 1667941163
transform 1 0 30452 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1345_
timestamp 1667941163
transform 1 0 33856 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1346_
timestamp 1667941163
transform 1 0 34868 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1347_
timestamp 1667941163
transform 1 0 32016 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1348_
timestamp 1667941163
transform 1 0 34040 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1349_
timestamp 1667941163
transform 1 0 33396 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1350_
timestamp 1667941163
transform 1 0 32844 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1351_
timestamp 1667941163
transform 1 0 33672 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1352_
timestamp 1667941163
transform 1 0 32476 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _1353_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 33212 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1354_
timestamp 1667941163
transform 1 0 33856 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1355_
timestamp 1667941163
transform 1 0 32292 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1356_
timestamp 1667941163
transform 1 0 33856 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1357_
timestamp 1667941163
transform 1 0 32476 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1358_
timestamp 1667941163
transform 1 0 33304 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1359_
timestamp 1667941163
transform 1 0 32752 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1360_
timestamp 1667941163
transform 1 0 29348 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1361_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 32292 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1362_
timestamp 1667941163
transform 1 0 32200 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _1363_
timestamp 1667941163
transform 1 0 32292 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__a31oi_1  _1364_
timestamp 1667941163
transform 1 0 32292 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1365_
timestamp 1667941163
transform 1 0 27600 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1366_
timestamp 1667941163
transform 1 0 25484 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1367_
timestamp 1667941163
transform 1 0 26496 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1368_
timestamp 1667941163
transform 1 0 26680 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1369_
timestamp 1667941163
transform 1 0 27140 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1370_
timestamp 1667941163
transform 1 0 26036 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1371_
timestamp 1667941163
transform 1 0 27140 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1372_
timestamp 1667941163
transform 1 0 27048 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1373_
timestamp 1667941163
transform 1 0 25116 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1374_
timestamp 1667941163
transform 1 0 25484 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1375_
timestamp 1667941163
transform 1 0 27140 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1376_
timestamp 1667941163
transform 1 0 26588 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _1377_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 25392 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1378_
timestamp 1667941163
transform 1 0 22356 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1379_
timestamp 1667941163
transform 1 0 22540 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1380_
timestamp 1667941163
transform 1 0 23552 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1381_
timestamp 1667941163
transform 1 0 23184 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1382_
timestamp 1667941163
transform 1 0 24104 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1383_
timestamp 1667941163
transform 1 0 22448 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1384_
timestamp 1667941163
transform 1 0 22264 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _1385_
timestamp 1667941163
transform 1 0 24196 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1386_
timestamp 1667941163
transform 1 0 23276 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1387_
timestamp 1667941163
transform 1 0 22632 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1388_
timestamp 1667941163
transform 1 0 24564 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1389_
timestamp 1667941163
transform 1 0 21804 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_4  _1390_
timestamp 1667941163
transform 1 0 22540 0 1 41344
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_4  _1391_
timestamp 1667941163
transform 1 0 24196 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _1392_
timestamp 1667941163
transform 1 0 16836 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1393_
timestamp 1667941163
transform 1 0 16836 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1394_
timestamp 1667941163
transform 1 0 15916 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1395_
timestamp 1667941163
transform 1 0 15916 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1396_
timestamp 1667941163
transform 1 0 17296 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1397_
timestamp 1667941163
transform 1 0 15548 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1398_
timestamp 1667941163
transform 1 0 14720 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1399_
timestamp 1667941163
transform 1 0 17020 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1400_
timestamp 1667941163
transform 1 0 19412 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1401_
timestamp 1667941163
transform 1 0 20516 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1402_
timestamp 1667941163
transform 1 0 19412 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1403_
timestamp 1667941163
transform 1 0 16928 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1404_
timestamp 1667941163
transform 1 0 16836 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1405_
timestamp 1667941163
transform 1 0 19412 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1406_
timestamp 1667941163
transform 1 0 19228 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1407_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19412 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1408_
timestamp 1667941163
transform 1 0 31188 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1409_
timestamp 1667941163
transform 1 0 31280 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1410_
timestamp 1667941163
transform 1 0 29900 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1411_
timestamp 1667941163
transform 1 0 30544 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1412_
timestamp 1667941163
transform 1 0 31832 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1413_
timestamp 1667941163
transform 1 0 31648 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1414_
timestamp 1667941163
transform 1 0 31096 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1415_
timestamp 1667941163
transform 1 0 28796 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _1416_
timestamp 1667941163
transform 1 0 25852 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1417_
timestamp 1667941163
transform 1 0 28796 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1418_
timestamp 1667941163
transform 1 0 27600 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1419_
timestamp 1667941163
transform 1 0 27508 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1420_
timestamp 1667941163
transform 1 0 19872 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1421_
timestamp 1667941163
transform 1 0 19412 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _1422_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 18768 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1423_
timestamp 1667941163
transform 1 0 20148 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1424_
timestamp 1667941163
transform 1 0 17664 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1425_
timestamp 1667941163
transform 1 0 16100 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1426_
timestamp 1667941163
transform 1 0 15548 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1427_
timestamp 1667941163
transform 1 0 13248 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1428_
timestamp 1667941163
transform 1 0 12696 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1429_
timestamp 1667941163
transform 1 0 15640 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1430_
timestamp 1667941163
transform 1 0 15364 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1431_
timestamp 1667941163
transform 1 0 14812 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1432_
timestamp 1667941163
transform 1 0 13432 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1433_
timestamp 1667941163
transform 1 0 12788 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1434_
timestamp 1667941163
transform 1 0 16560 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1435_
timestamp 1667941163
transform 1 0 18032 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1436_
timestamp 1667941163
transform 1 0 16836 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1437_
timestamp 1667941163
transform 1 0 16192 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1438_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17020 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1439_
timestamp 1667941163
transform 1 0 18216 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  _1440_
timestamp 1667941163
transform 1 0 13432 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1441_
timestamp 1667941163
transform 1 0 14168 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1442_
timestamp 1667941163
transform 1 0 14536 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1443_
timestamp 1667941163
transform 1 0 15180 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1444_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14352 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1445_
timestamp 1667941163
transform 1 0 12972 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1446_
timestamp 1667941163
transform 1 0 12512 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1447_
timestamp 1667941163
transform 1 0 15732 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1448_
timestamp 1667941163
transform 1 0 18676 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1449_
timestamp 1667941163
transform 1 0 17664 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1450_
timestamp 1667941163
transform 1 0 17664 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1451_
timestamp 1667941163
transform 1 0 18584 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1452_
timestamp 1667941163
transform 1 0 16008 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1453_
timestamp 1667941163
transform 1 0 16928 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1454_
timestamp 1667941163
transform 1 0 15272 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1455_
timestamp 1667941163
transform 1 0 15364 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1456_
timestamp 1667941163
transform 1 0 13800 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1457_
timestamp 1667941163
transform 1 0 12420 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1458_
timestamp 1667941163
transform 1 0 17572 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1459_
timestamp 1667941163
transform 1 0 22908 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1460_
timestamp 1667941163
transform 1 0 21988 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1461_
timestamp 1667941163
transform 1 0 22724 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1462_
timestamp 1667941163
transform 1 0 23184 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1463_
timestamp 1667941163
transform 1 0 20976 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1464_
timestamp 1667941163
transform 1 0 22080 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1465_
timestamp 1667941163
transform 1 0 22172 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1466_
timestamp 1667941163
transform 1 0 22080 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1467_
timestamp 1667941163
transform 1 0 20424 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1468_
timestamp 1667941163
transform 1 0 19964 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1469_
timestamp 1667941163
transform 1 0 23000 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1470_
timestamp 1667941163
transform 1 0 22264 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _1471_
timestamp 1667941163
transform 1 0 21344 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1472_
timestamp 1667941163
transform 1 0 21804 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1473_
timestamp 1667941163
transform 1 0 22632 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1474_
timestamp 1667941163
transform 1 0 22632 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1475_
timestamp 1667941163
transform 1 0 22356 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1476_
timestamp 1667941163
transform 1 0 22724 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1477_
timestamp 1667941163
transform 1 0 22172 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1478_
timestamp 1667941163
transform 1 0 23460 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1479_
timestamp 1667941163
transform 1 0 24840 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1480_
timestamp 1667941163
transform 1 0 24564 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1481_
timestamp 1667941163
transform 1 0 25024 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1482_
timestamp 1667941163
transform 1 0 25208 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1483_
timestamp 1667941163
transform 1 0 24656 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1484_
timestamp 1667941163
transform 1 0 24380 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1485_
timestamp 1667941163
transform 1 0 26404 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1486_
timestamp 1667941163
transform 1 0 25944 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1487_
timestamp 1667941163
transform 1 0 25668 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1488_
timestamp 1667941163
transform 1 0 26680 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1489_
timestamp 1667941163
transform 1 0 25852 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1490_
timestamp 1667941163
transform 1 0 27048 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _1491_
timestamp 1667941163
transform 1 0 23920 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1492_
timestamp 1667941163
transform 1 0 23092 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1493_
timestamp 1667941163
transform 1 0 23368 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1494_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24564 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1495_
timestamp 1667941163
transform 1 0 23368 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _1496_
timestamp 1667941163
transform 1 0 23184 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1497_
timestamp 1667941163
transform 1 0 31004 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1498_
timestamp 1667941163
transform 1 0 27416 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1499_
timestamp 1667941163
transform 1 0 33396 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1500_
timestamp 1667941163
transform 1 0 32568 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1501_
timestamp 1667941163
transform 1 0 33672 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1502_
timestamp 1667941163
transform 1 0 32752 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1503_
timestamp 1667941163
transform 1 0 33672 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1504_
timestamp 1667941163
transform 1 0 33580 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1505_
timestamp 1667941163
transform 1 0 32292 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1506_
timestamp 1667941163
transform 1 0 31280 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1507_
timestamp 1667941163
transform 1 0 25484 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1508_
timestamp 1667941163
transform 1 0 22448 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1509_
timestamp 1667941163
transform 1 0 29716 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1510_
timestamp 1667941163
transform 1 0 29348 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1511_
timestamp 1667941163
transform 1 0 31004 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1512_
timestamp 1667941163
transform 1 0 30820 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1513_
timestamp 1667941163
transform 1 0 30820 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1514_
timestamp 1667941163
transform 1 0 30084 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1515_
timestamp 1667941163
transform 1 0 30820 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1516_
timestamp 1667941163
transform 1 0 30452 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1517_
timestamp 1667941163
transform 1 0 27508 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1518_
timestamp 1667941163
transform 1 0 27140 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1519_
timestamp 1667941163
transform 1 0 22264 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1520_
timestamp 1667941163
transform 1 0 22172 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1521_
timestamp 1667941163
transform 1 0 27600 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1522_
timestamp 1667941163
transform 1 0 27140 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1523_
timestamp 1667941163
transform 1 0 21988 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1524_
timestamp 1667941163
transform 1 0 21988 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1525_
timestamp 1667941163
transform 1 0 21988 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1526_
timestamp 1667941163
transform 1 0 22632 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1527_
timestamp 1667941163
transform 1 0 21988 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1528_
timestamp 1667941163
transform 1 0 20976 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1529_
timestamp 1667941163
transform 1 0 32292 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1530_
timestamp 1667941163
transform 1 0 30360 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1531_
timestamp 1667941163
transform 1 0 29716 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1532_
timestamp 1667941163
transform 1 0 32200 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1533_
timestamp 1667941163
transform 1 0 32476 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1534_
timestamp 1667941163
transform 1 0 9108 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1535_
timestamp 1667941163
transform 1 0 6532 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1536_
timestamp 1667941163
transform 1 0 7452 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1537_
timestamp 1667941163
transform 1 0 7268 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1538_
timestamp 1667941163
transform 1 0 8188 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1539_
timestamp 1667941163
transform 1 0 9476 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1540_
timestamp 1667941163
transform 1 0 8556 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1541_
timestamp 1667941163
transform 1 0 8188 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1542_
timestamp 1667941163
transform 1 0 5520 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1543_
timestamp 1667941163
transform 1 0 5980 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1544_
timestamp 1667941163
transform 1 0 5060 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1545_
timestamp 1667941163
transform 1 0 4876 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1546_
timestamp 1667941163
transform 1 0 5152 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1547_
timestamp 1667941163
transform 1 0 4968 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1548_
timestamp 1667941163
transform 1 0 4508 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1549_
timestamp 1667941163
transform 1 0 6348 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1550_
timestamp 1667941163
transform 1 0 5428 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1551_
timestamp 1667941163
transform 1 0 6532 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1552_
timestamp 1667941163
transform 1 0 6808 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1553_
timestamp 1667941163
transform 1 0 7728 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1554_
timestamp 1667941163
transform 1 0 8096 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1555_
timestamp 1667941163
transform 1 0 7360 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1556_
timestamp 1667941163
transform 1 0 32384 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1557_
timestamp 1667941163
transform 1 0 29624 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1558_
timestamp 1667941163
transform 1 0 30452 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1559_
timestamp 1667941163
transform 1 0 29716 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1560_
timestamp 1667941163
transform 1 0 32660 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1561_
timestamp 1667941163
transform 1 0 36524 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1562_
timestamp 1667941163
transform 1 0 37812 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1563_
timestamp 1667941163
transform 1 0 36984 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1564_
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1565_
timestamp 1667941163
transform 1 0 37444 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1566_
timestamp 1667941163
transform 1 0 36156 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1567_
timestamp 1667941163
transform 1 0 36984 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1568_
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1569_
timestamp 1667941163
transform 1 0 36064 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1570_
timestamp 1667941163
transform 1 0 35144 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1571_
timestamp 1667941163
transform 1 0 35328 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1572_
timestamp 1667941163
transform 1 0 39192 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1573_
timestamp 1667941163
transform 1 0 39100 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1574_
timestamp 1667941163
transform 1 0 39284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1575_
timestamp 1667941163
transform 1 0 38732 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1576_
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1577_
timestamp 1667941163
transform 1 0 36432 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1578_
timestamp 1667941163
transform 1 0 37444 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _1579_
timestamp 1667941163
transform 1 0 36616 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1580_
timestamp 1667941163
transform 1 0 37720 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1581_
timestamp 1667941163
transform 1 0 37996 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1582_
timestamp 1667941163
transform 1 0 41308 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1583_
timestamp 1667941163
transform 1 0 42044 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1584_
timestamp 1667941163
transform 1 0 41032 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1585_
timestamp 1667941163
transform 1 0 40112 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1586_
timestamp 1667941163
transform 1 0 40204 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o41a_1  _1587_
timestamp 1667941163
transform 1 0 38640 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a2111oi_4  _1588_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37536 0 1 10880
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _1589_
timestamp 1667941163
transform 1 0 43516 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1590_
timestamp 1667941163
transform 1 0 44252 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1591_
timestamp 1667941163
transform 1 0 44160 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1592_
timestamp 1667941163
transform 1 0 42780 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1593_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 42872 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1594_
timestamp 1667941163
transform 1 0 44896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1595_
timestamp 1667941163
transform 1 0 45172 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1596_
timestamp 1667941163
transform 1 0 43240 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1597_
timestamp 1667941163
transform 1 0 44252 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1598_
timestamp 1667941163
transform 1 0 44160 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1599_
timestamp 1667941163
transform 1 0 43056 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1600_
timestamp 1667941163
transform 1 0 43332 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1601_
timestamp 1667941163
transform 1 0 44068 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1602_
timestamp 1667941163
transform 1 0 45172 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1603_
timestamp 1667941163
transform 1 0 44896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1604_
timestamp 1667941163
transform 1 0 44252 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1605_
timestamp 1667941163
transform 1 0 43608 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1606_
timestamp 1667941163
transform 1 0 44344 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1607_
timestamp 1667941163
transform 1 0 45172 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1608_
timestamp 1667941163
transform 1 0 43516 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1609_
timestamp 1667941163
transform 1 0 44344 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1610_
timestamp 1667941163
transform 1 0 43884 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1611_
timestamp 1667941163
transform 1 0 43240 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _1612_
timestamp 1667941163
transform 1 0 44436 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1613_
timestamp 1667941163
transform 1 0 43700 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1614_
timestamp 1667941163
transform 1 0 43056 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1615_
timestamp 1667941163
transform 1 0 42688 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1616_
timestamp 1667941163
transform 1 0 40940 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1617_
timestamp 1667941163
transform 1 0 42228 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1618_
timestamp 1667941163
transform 1 0 40756 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _1619_
timestamp 1667941163
transform 1 0 41492 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1620_
timestamp 1667941163
transform 1 0 41216 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1621_
timestamp 1667941163
transform 1 0 40020 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1622_
timestamp 1667941163
transform 1 0 41124 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1623_
timestamp 1667941163
transform 1 0 42596 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1624_
timestamp 1667941163
transform 1 0 41584 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1625_
timestamp 1667941163
transform 1 0 41400 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1626_
timestamp 1667941163
transform 1 0 40112 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1627_
timestamp 1667941163
transform 1 0 39284 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _1628_
timestamp 1667941163
transform 1 0 42596 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1629_
timestamp 1667941163
transform 1 0 41492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1630_
timestamp 1667941163
transform 1 0 41400 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1631_
timestamp 1667941163
transform 1 0 40848 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1632_
timestamp 1667941163
transform 1 0 43976 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1633_
timestamp 1667941163
transform 1 0 42780 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1634_
timestamp 1667941163
transform 1 0 43424 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1635_
timestamp 1667941163
transform 1 0 43424 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_1  _1636_
timestamp 1667941163
transform 1 0 42412 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1637_
timestamp 1667941163
transform 1 0 42780 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1638_
timestamp 1667941163
transform 1 0 42872 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1639_
timestamp 1667941163
transform 1 0 43700 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1640_
timestamp 1667941163
transform 1 0 43240 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1641_
timestamp 1667941163
transform 1 0 43608 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1642_
timestamp 1667941163
transform 1 0 45172 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1643_
timestamp 1667941163
transform 1 0 44160 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1644_
timestamp 1667941163
transform 1 0 44252 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _1645_
timestamp 1667941163
transform 1 0 43976 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1646_
timestamp 1667941163
transform 1 0 44068 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1647_
timestamp 1667941163
transform 1 0 41860 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _1648_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 43148 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1649_
timestamp 1667941163
transform 1 0 42596 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1650_
timestamp 1667941163
transform 1 0 22540 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1651_
timestamp 1667941163
transform 1 0 22080 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1652_
timestamp 1667941163
transform 1 0 20148 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1653_
timestamp 1667941163
transform 1 0 19780 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1654_
timestamp 1667941163
transform 1 0 21252 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1655_
timestamp 1667941163
transform 1 0 18032 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1656_
timestamp 1667941163
transform 1 0 21160 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1657_
timestamp 1667941163
transform 1 0 20240 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1658_
timestamp 1667941163
transform 1 0 22356 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1659_
timestamp 1667941163
transform 1 0 20240 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1660_
timestamp 1667941163
transform 1 0 19688 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1661_
timestamp 1667941163
transform 1 0 19780 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1662_
timestamp 1667941163
transform 1 0 17756 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1663_
timestamp 1667941163
transform 1 0 16836 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1664_
timestamp 1667941163
transform 1 0 17756 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1665_
timestamp 1667941163
transform 1 0 18032 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1666_
timestamp 1667941163
transform 1 0 17020 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1667_
timestamp 1667941163
transform 1 0 16928 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1668_
timestamp 1667941163
transform -1 0 18308 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1669_
timestamp 1667941163
transform 1 0 18676 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1670_
timestamp 1667941163
transform 1 0 18216 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1671_
timestamp 1667941163
transform 1 0 19412 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1672_
timestamp 1667941163
transform 1 0 18492 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1673_
timestamp 1667941163
transform 1 0 19136 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1674_
timestamp 1667941163
transform 1 0 17020 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1675_
timestamp 1667941163
transform 1 0 16836 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1676_
timestamp 1667941163
transform 1 0 16100 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1677_
timestamp 1667941163
transform 1 0 17112 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1678_
timestamp 1667941163
transform 1 0 18308 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1679_
timestamp 1667941163
transform 1 0 16836 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1680_
timestamp 1667941163
transform 1 0 18676 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1681_
timestamp 1667941163
transform 1 0 18308 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1682_
timestamp 1667941163
transform 1 0 19412 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1683_
timestamp 1667941163
transform 1 0 24472 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1684_
timestamp 1667941163
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_2  _1685_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 23092 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1686_
timestamp 1667941163
transform 1 0 24564 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1687_
timestamp 1667941163
transform 1 0 25760 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1688_
timestamp 1667941163
transform 1 0 25576 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1689_
timestamp 1667941163
transform 1 0 24564 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1690_
timestamp 1667941163
transform 1 0 24564 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1691_
timestamp 1667941163
transform 1 0 24380 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1692_
timestamp 1667941163
transform 1 0 25208 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1693_
timestamp 1667941163
transform 1 0 24288 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1694_
timestamp 1667941163
transform 1 0 23460 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1695_
timestamp 1667941163
transform 1 0 23092 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1696_
timestamp 1667941163
transform 1 0 26956 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1697_
timestamp 1667941163
transform 1 0 37904 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1698_
timestamp 1667941163
transform 1 0 39008 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1699_
timestamp 1667941163
transform 1 0 37444 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1700_
timestamp 1667941163
transform 1 0 38548 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1701_
timestamp 1667941163
transform 1 0 38088 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1702_
timestamp 1667941163
transform 1 0 37996 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1703_
timestamp 1667941163
transform 1 0 31096 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1704_
timestamp 1667941163
transform 1 0 31280 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1705_
timestamp 1667941163
transform 1 0 29808 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1706_
timestamp 1667941163
transform 1 0 29900 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1707_
timestamp 1667941163
transform 1 0 37628 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1708_
timestamp 1667941163
transform 1 0 37720 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1709_
timestamp 1667941163
transform 1 0 38456 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1710_
timestamp 1667941163
transform 1 0 38640 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1711_
timestamp 1667941163
transform 1 0 30820 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1712_
timestamp 1667941163
transform 1 0 32292 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1713_
timestamp 1667941163
transform 1 0 30084 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1714_
timestamp 1667941163
transform 1 0 26588 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1715_
timestamp 1667941163
transform 1 0 27140 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1716_
timestamp 1667941163
transform 1 0 22724 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1717_
timestamp 1667941163
transform 1 0 24564 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1718_
timestamp 1667941163
transform 1 0 24748 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1719_
timestamp 1667941163
transform 1 0 24656 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1720_
timestamp 1667941163
transform 1 0 23184 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1721_
timestamp 1667941163
transform 1 0 23184 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1722_
timestamp 1667941163
transform 1 0 22264 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1723_
timestamp 1667941163
transform 1 0 22448 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1724_
timestamp 1667941163
transform 1 0 22540 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1725_
timestamp 1667941163
transform 1 0 22356 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1726_
timestamp 1667941163
transform 1 0 24288 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1727_
timestamp 1667941163
transform 1 0 24564 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1728_
timestamp 1667941163
transform 1 0 25024 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1729_
timestamp 1667941163
transform 1 0 25392 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1730_
timestamp 1667941163
transform 1 0 37168 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1731_
timestamp 1667941163
transform 1 0 23092 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1732_
timestamp 1667941163
transform 1 0 23276 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1733_
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _1734_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24656 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1735_
timestamp 1667941163
transform 1 0 26220 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1736_
timestamp 1667941163
transform 1 0 30360 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1737_
timestamp 1667941163
transform 1 0 30176 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1738_
timestamp 1667941163
transform 1 0 30636 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1739_
timestamp 1667941163
transform 1 0 30636 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1740_
timestamp 1667941163
transform 1 0 25484 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1741_
timestamp 1667941163
transform 1 0 27140 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1742_
timestamp 1667941163
transform 1 0 27140 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1743_
timestamp 1667941163
transform 1 0 18216 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1744_
timestamp 1667941163
transform 1 0 18032 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1745_
timestamp 1667941163
transform 1 0 12328 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1746_
timestamp 1667941163
transform 1 0 11960 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1747_
timestamp 1667941163
transform 1 0 14720 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1748_
timestamp 1667941163
transform 1 0 14260 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1749_
timestamp 1667941163
transform 1 0 18400 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1750_
timestamp 1667941163
transform 1 0 17848 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1751_
timestamp 1667941163
transform 1 0 12512 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1752_
timestamp 1667941163
transform 1 0 12328 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1753_
timestamp 1667941163
transform 1 0 15456 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1754_
timestamp 1667941163
transform 1 0 16652 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1755_
timestamp 1667941163
transform 1 0 12420 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1756_
timestamp 1667941163
transform 1 0 12144 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1757_
timestamp 1667941163
transform 1 0 25852 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1758_
timestamp 1667941163
transform 1 0 26128 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1759_
timestamp 1667941163
transform 1 0 20516 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1760_
timestamp 1667941163
transform 1 0 20332 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1761_
timestamp 1667941163
transform 1 0 20424 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1762_
timestamp 1667941163
transform 1 0 19964 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1763_
timestamp 1667941163
transform 1 0 27692 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1764_
timestamp 1667941163
transform 1 0 21068 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1765_
timestamp 1667941163
transform 1 0 20148 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1766_
timestamp 1667941163
transform 1 0 26772 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1767_
timestamp 1667941163
transform 1 0 27140 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1768_
timestamp 1667941163
transform 1 0 26956 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1769_
timestamp 1667941163
transform 1 0 26956 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1770_
timestamp 1667941163
transform 1 0 28244 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1771_
timestamp 1667941163
transform 1 0 24288 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1772_
timestamp 1667941163
transform 1 0 24656 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1773_
timestamp 1667941163
transform 1 0 24564 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1774_
timestamp 1667941163
transform 1 0 28520 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1775_
timestamp 1667941163
transform 1 0 28980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1776_
timestamp 1667941163
transform 1 0 28520 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1777_
timestamp 1667941163
transform 1 0 28428 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1778_
timestamp 1667941163
transform 1 0 28520 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1779_
timestamp 1667941163
transform 1 0 28704 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1780_
timestamp 1667941163
transform 1 0 17756 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1781_
timestamp 1667941163
transform 1 0 17480 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1782_
timestamp 1667941163
transform 1 0 15456 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1783_
timestamp 1667941163
transform 1 0 15180 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1784_
timestamp 1667941163
transform 1 0 14352 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1785_
timestamp 1667941163
transform 1 0 13892 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1786_
timestamp 1667941163
transform 1 0 21528 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1787_
timestamp 1667941163
transform 1 0 21160 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1788_
timestamp 1667941163
transform 1 0 21988 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1789_
timestamp 1667941163
transform 1 0 15640 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1790_
timestamp 1667941163
transform 1 0 14352 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1791_
timestamp 1667941163
transform 1 0 19412 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1792_
timestamp 1667941163
transform 1 0 18400 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1793_
timestamp 1667941163
transform 1 0 16376 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1794_
timestamp 1667941163
transform 1 0 16836 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1795_
timestamp 1667941163
transform 1 0 24380 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1796_
timestamp 1667941163
transform 1 0 24380 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1797_
timestamp 1667941163
transform 1 0 22448 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1798_
timestamp 1667941163
transform 1 0 22264 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1799_
timestamp 1667941163
transform 1 0 21620 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1800_
timestamp 1667941163
transform 1 0 20976 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1801_
timestamp 1667941163
transform 1 0 22448 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1802_
timestamp 1667941163
transform 1 0 22080 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1803_
timestamp 1667941163
transform 1 0 24656 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1804_
timestamp 1667941163
transform 1 0 23552 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1805_
timestamp 1667941163
transform 1 0 24840 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1806_
timestamp 1667941163
transform 1 0 23920 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1807_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 40020 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1808_
timestamp 1667941163
transform 1 0 40020 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1809_
timestamp 1667941163
transform 1 0 36156 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1810_
timestamp 1667941163
transform 1 0 33212 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1811_
timestamp 1667941163
transform 1 0 30544 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1812_
timestamp 1667941163
transform 1 0 35880 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1813_
timestamp 1667941163
transform 1 0 37444 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1814_
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1815_
timestamp 1667941163
transform 1 0 28980 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1816_
timestamp 1667941163
transform 1 0 25208 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1817_
timestamp 1667941163
transform 1 0 28704 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1818_
timestamp 1667941163
transform 1 0 23000 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1819_
timestamp 1667941163
transform 1 0 26496 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1820_
timestamp 1667941163
transform 1 0 26128 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1821_
timestamp 1667941163
transform 1 0 31004 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1822_
timestamp 1667941163
transform 1 0 33856 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1823_
timestamp 1667941163
transform 1 0 34960 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1824_
timestamp 1667941163
transform 1 0 35052 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1825_
timestamp 1667941163
transform 1 0 29256 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1826_
timestamp 1667941163
transform 1 0 27784 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1827_
timestamp 1667941163
transform 1 0 28980 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1828_
timestamp 1667941163
transform 1 0 35052 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1829_
timestamp 1667941163
transform 1 0 34868 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1830_
timestamp 1667941163
transform 1 0 30912 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1831_
timestamp 1667941163
transform 1 0 27140 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1832_
timestamp 1667941163
transform 1 0 25208 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1833_
timestamp 1667941163
transform 1 0 20608 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1834_
timestamp 1667941163
transform 1 0 20792 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1835_
timestamp 1667941163
transform 1 0 15456 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1836_
timestamp 1667941163
transform 1 0 14076 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1837_
timestamp 1667941163
transform 1 0 18768 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1838_
timestamp 1667941163
transform 1 0 18400 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1839_
timestamp 1667941163
transform 1 0 30268 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1840_
timestamp 1667941163
transform 1 0 32292 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1841_
timestamp 1667941163
transform 1 0 27324 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1842_
timestamp 1667941163
transform 1 0 18308 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1843_
timestamp 1667941163
transform 1 0 12328 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1844_
timestamp 1667941163
transform 1 0 12328 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1845_
timestamp 1667941163
transform 1 0 17480 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1846_
timestamp 1667941163
transform 1 0 12052 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1847_
timestamp 1667941163
transform 1 0 19412 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1848_
timestamp 1667941163
transform 1 0 11960 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1849_
timestamp 1667941163
transform 1 0 24288 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1850_
timestamp 1667941163
transform 1 0 19412 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1851_
timestamp 1667941163
transform 1 0 21988 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1852_
timestamp 1667941163
transform 1 0 20792 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1853_
timestamp 1667941163
transform 1 0 24564 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1854_
timestamp 1667941163
transform 1 0 27140 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1855_
timestamp 1667941163
transform 1 0 32292 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1856_
timestamp 1667941163
transform 1 0 33672 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1857_
timestamp 1667941163
transform 1 0 33764 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1858_
timestamp 1667941163
transform 1 0 31096 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1859_
timestamp 1667941163
transform 1 0 29164 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1860_
timestamp 1667941163
transform 1 0 30636 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1861_
timestamp 1667941163
transform 1 0 30360 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1862_
timestamp 1667941163
transform 1 0 30268 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1863_
timestamp 1667941163
transform 1 0 27048 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1864_
timestamp 1667941163
transform 1 0 21804 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1865_
timestamp 1667941163
transform 1 0 27140 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1866_
timestamp 1667941163
transform 1 0 20792 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1867_
timestamp 1667941163
transform 1 0 20700 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1868_
timestamp 1667941163
transform 1 0 20792 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1869_
timestamp 1667941163
transform 1 0 29716 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1870_
timestamp 1667941163
transform 1 0 32292 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1871_
timestamp 1667941163
transform 1 0 15272 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1872_
timestamp 1667941163
transform 1 0 11868 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1873_
timestamp 1667941163
transform 1 0 12236 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1874_
timestamp 1667941163
transform 1 0 14168 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1875_
timestamp 1667941163
transform 1 0 14904 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1876_
timestamp 1667941163
transform 1 0 14260 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1877_
timestamp 1667941163
transform 1 0 13800 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1878_
timestamp 1667941163
transform 1 0 12052 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1879_
timestamp 1667941163
transform 1 0 11500 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1880_
timestamp 1667941163
transform 1 0 11684 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1881_
timestamp 1667941163
transform 1 0 6900 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1882_
timestamp 1667941163
transform 1 0 9108 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1883_
timestamp 1667941163
transform 1 0 7176 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1884_
timestamp 1667941163
transform 1 0 4324 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1885_
timestamp 1667941163
transform 1 0 4324 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1886_
timestamp 1667941163
transform 1 0 4324 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1887_
timestamp 1667941163
transform 1 0 4324 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1888_
timestamp 1667941163
transform 1 0 5244 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1889_
timestamp 1667941163
transform 1 0 7084 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1890_
timestamp 1667941163
transform 1 0 8004 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1891_
timestamp 1667941163
transform 1 0 37444 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1892_
timestamp 1667941163
transform 1 0 34868 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1893_
timestamp 1667941163
transform 1 0 37444 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1894_
timestamp 1667941163
transform 1 0 40204 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1895_
timestamp 1667941163
transform 1 0 45172 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1896_
timestamp 1667941163
transform 1 0 42688 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1897_
timestamp 1667941163
transform 1 0 45632 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1898_
timestamp 1667941163
transform 1 0 42596 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1899_
timestamp 1667941163
transform 1 0 39376 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1900_
timestamp 1667941163
transform 1 0 39744 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1901_
timestamp 1667941163
transform 1 0 40388 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1902_
timestamp 1667941163
transform 1 0 43516 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1903_
timestamp 1667941163
transform 1 0 43700 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1904_
timestamp 1667941163
transform 1 0 44344 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1905_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 44804 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1906_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 41860 0 1 19584
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1907_
timestamp 1667941163
transform 1 0 19412 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1908_
timestamp 1667941163
transform 1 0 20056 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1909_
timestamp 1667941163
transform 1 0 19320 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1910_
timestamp 1667941163
transform 1 0 17388 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1911_
timestamp 1667941163
transform 1 0 16008 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1912_
timestamp 1667941163
transform 1 0 16928 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1913_
timestamp 1667941163
transform 1 0 18492 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1914_
timestamp 1667941163
transform 1 0 16008 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1915_
timestamp 1667941163
transform 1 0 16376 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1916_
timestamp 1667941163
transform 1 0 18400 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1917_
timestamp 1667941163
transform 1 0 25116 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1918_
timestamp 1667941163
transform 1 0 23828 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1919_
timestamp 1667941163
transform 1 0 39284 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1920_
timestamp 1667941163
transform 1 0 38088 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1921_
timestamp 1667941163
transform 1 0 37628 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1922_
timestamp 1667941163
transform 1 0 31188 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1923_
timestamp 1667941163
transform 1 0 29440 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1924_
timestamp 1667941163
transform 1 0 37444 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1925_
timestamp 1667941163
transform 1 0 38088 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1926_
timestamp 1667941163
transform 1 0 32108 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1927_
timestamp 1667941163
transform 1 0 27140 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1928_
timestamp 1667941163
transform 1 0 23368 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1929_
timestamp 1667941163
transform 1 0 24288 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1930_
timestamp 1667941163
transform 1 0 22632 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1931_
timestamp 1667941163
transform 1 0 21896 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1932_
timestamp 1667941163
transform 1 0 21804 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1933_
timestamp 1667941163
transform 1 0 23920 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1934_
timestamp 1667941163
transform 1 0 24656 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1935_
timestamp 1667941163
transform 1 0 37444 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1936_
timestamp 1667941163
transform 1 0 29900 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1937_
timestamp 1667941163
transform 1 0 30728 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1938_
timestamp 1667941163
transform 1 0 27140 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1939_
timestamp 1667941163
transform 1 0 17480 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1940_
timestamp 1667941163
transform 1 0 11776 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1941_
timestamp 1667941163
transform 1 0 12880 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1942_
timestamp 1667941163
transform 1 0 16560 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1943_
timestamp 1667941163
transform 1 0 12052 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1944_
timestamp 1667941163
transform 1 0 14812 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1945_
timestamp 1667941163
transform 1 0 11960 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1946_
timestamp 1667941163
transform 1 0 25392 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1947_
timestamp 1667941163
transform 1 0 19688 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1948_
timestamp 1667941163
transform 1 0 19504 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1949_
timestamp 1667941163
transform 1 0 20056 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1950_
timestamp 1667941163
transform 1 0 27140 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1951_
timestamp 1667941163
transform 1 0 27140 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1952_
timestamp 1667941163
transform 1 0 28520 0 -1 36992
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1953_
timestamp 1667941163
transform 1 0 28336 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1954_
timestamp 1667941163
transform 1 0 28980 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1955_
timestamp 1667941163
transform 1 0 28980 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1956_
timestamp 1667941163
transform 1 0 17204 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1957_
timestamp 1667941163
transform 1 0 14812 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1958_
timestamp 1667941163
transform 1 0 14260 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1959_
timestamp 1667941163
transform 1 0 20608 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1960_
timestamp 1667941163
transform 1 0 13800 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1961_
timestamp 1667941163
transform 1 0 18124 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1962_
timestamp 1667941163
transform 1 0 15732 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1963_
timestamp 1667941163
transform 1 0 24564 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1964_
timestamp 1667941163
transform 1 0 21988 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1965_
timestamp 1667941163
transform 1 0 20516 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1966_
timestamp 1667941163
transform 1 0 21988 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1967_
timestamp 1667941163
transform 1 0 24564 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1968_
timestamp 1667941163
transform 1 0 24564 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _2066__29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 7268 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2066_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 7268 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2067_
timestamp 1667941163
transform 1 0 2024 0 -1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2067__30
timestamp 1667941163
transform 1 0 2852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2068__31
timestamp 1667941163
transform 1 0 20608 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2068_
timestamp 1667941163
transform 1 0 19688 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2069__32
timestamp 1667941163
transform 1 0 2116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2069_
timestamp 1667941163
transform 1 0 2024 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2070__33
timestamp 1667941163
transform 1 0 44436 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2070_
timestamp 1667941163
transform 1 0 44896 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2071_
timestamp 1667941163
transform 1 0 3772 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2071__34
timestamp 1667941163
transform 1 0 2576 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2072__35
timestamp 1667941163
transform 1 0 47748 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2072_
timestamp 1667941163
transform 1 0 46460 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2073_
timestamp 1667941163
transform 1 0 10212 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2074_
timestamp 1667941163
transform 1 0 46184 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2075_
timestamp 1667941163
transform 1 0 45908 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2076_
timestamp 1667941163
transform 1 0 46460 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2077_
timestamp 1667941163
transform 1 0 21988 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2078_
timestamp 1667941163
transform 1 0 17204 0 -1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2079_
timestamp 1667941163
transform 1 0 4876 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2080_
timestamp 1667941163
transform 1 0 20332 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2081_
timestamp 1667941163
transform 1 0 3772 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2082_
timestamp 1667941163
transform 1 0 45356 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2082__36
timestamp 1667941163
transform 1 0 47748 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2083__37
timestamp 1667941163
transform 1 0 47748 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2083_
timestamp 1667941163
transform 1 0 46460 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2084__38
timestamp 1667941163
transform 1 0 6532 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2084_
timestamp 1667941163
transform 1 0 5244 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2085__39
timestamp 1667941163
transform 1 0 47012 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2085_
timestamp 1667941163
transform 1 0 46460 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2086__40
timestamp 1667941163
transform 1 0 2852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2086_
timestamp 1667941163
transform 1 0 2668 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2087__41
timestamp 1667941163
transform 1 0 47012 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2087_
timestamp 1667941163
transform 1 0 46460 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2088__42
timestamp 1667941163
transform 1 0 29808 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2088_
timestamp 1667941163
transform 1 0 29716 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2089__43
timestamp 1667941163
transform 1 0 12328 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2089_
timestamp 1667941163
transform 1 0 12328 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2090__44
timestamp 1667941163
transform 1 0 47748 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2090_
timestamp 1667941163
transform 1 0 46460 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2091__45
timestamp 1667941163
transform 1 0 2944 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2091_
timestamp 1667941163
transform 1 0 1564 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2092_
timestamp 1667941163
transform 1 0 46460 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2092__46
timestamp 1667941163
transform 1 0 47012 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2093__47
timestamp 1667941163
transform 1 0 7820 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2093_
timestamp 1667941163
transform 1 0 1564 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2094__48
timestamp 1667941163
transform 1 0 44068 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2094_
timestamp 1667941163
transform 1 0 45172 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2095__49
timestamp 1667941163
transform 1 0 5336 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2095_
timestamp 1667941163
transform 1 0 5980 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2096__50
timestamp 1667941163
transform 1 0 47748 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2096_
timestamp 1667941163
transform 1 0 46460 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2097_
timestamp 1667941163
transform 1 0 45356 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2097__51
timestamp 1667941163
transform 1 0 45632 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2098_
timestamp 1667941163
transform 1 0 46460 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2098__52
timestamp 1667941163
transform 1 0 46276 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2099__53
timestamp 1667941163
transform 1 0 33028 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2099_
timestamp 1667941163
transform 1 0 32844 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2100_
timestamp 1667941163
transform 1 0 6624 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2100__54
timestamp 1667941163
transform 1 0 6624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2101_
timestamp 1667941163
transform 1 0 1564 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2101__55
timestamp 1667941163
transform 1 0 1656 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2102__56
timestamp 1667941163
transform 1 0 47012 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2102_
timestamp 1667941163
transform 1 0 46460 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2103__57
timestamp 1667941163
transform 1 0 22724 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2103_
timestamp 1667941163
transform 1 0 22448 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2104_
timestamp 1667941163
transform 1 0 45356 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2104__58
timestamp 1667941163
transform 1 0 45172 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2105__59
timestamp 1667941163
transform 1 0 4324 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2105_
timestamp 1667941163
transform 1 0 4140 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2106__60
timestamp 1667941163
transform 1 0 18400 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2106_
timestamp 1667941163
transform 1 0 17296 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2107_
timestamp 1667941163
transform 1 0 1564 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2107__61
timestamp 1667941163
transform 1 0 2116 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2108__62
timestamp 1667941163
transform 1 0 47012 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2108_
timestamp 1667941163
transform 1 0 46460 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2109__63
timestamp 1667941163
transform 1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2109_
timestamp 1667941163
transform 1 0 1840 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2110__64
timestamp 1667941163
transform 1 0 2116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2110_
timestamp 1667941163
transform 1 0 2024 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2111__65
timestamp 1667941163
transform 1 0 40020 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2111_
timestamp 1667941163
transform 1 0 39928 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2112__66
timestamp 1667941163
transform 1 0 47748 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2112_
timestamp 1667941163
transform 1 0 46460 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2113__67
timestamp 1667941163
transform 1 0 2024 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2113_
timestamp 1667941163
transform 1 0 2024 0 -1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2114__68
timestamp 1667941163
transform 1 0 47748 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2114_
timestamp 1667941163
transform 1 0 46460 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2115__69
timestamp 1667941163
transform 1 0 45816 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2115_
timestamp 1667941163
transform 1 0 45356 0 -1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2116_
timestamp 1667941163
transform 1 0 45908 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2116__70
timestamp 1667941163
transform 1 0 43792 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2117_
timestamp 1667941163
transform 1 0 10120 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2118__71
timestamp 1667941163
transform 1 0 40020 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2118_
timestamp 1667941163
transform 1 0 40020 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2119_
timestamp 1667941163
transform 1 0 10028 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2120__72
timestamp 1667941163
transform 1 0 31832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2120_
timestamp 1667941163
transform 1 0 32292 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2121__73
timestamp 1667941163
transform 1 0 41308 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2121_
timestamp 1667941163
transform 1 0 41308 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2122__74
timestamp 1667941163
transform 1 0 27232 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2122_
timestamp 1667941163
transform 1 0 27140 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2123_
timestamp 1667941163
transform 1 0 37444 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2123__75
timestamp 1667941163
transform 1 0 36248 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2124__76
timestamp 1667941163
transform 1 0 9568 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2124_
timestamp 1667941163
transform 1 0 9844 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2125__77
timestamp 1667941163
transform 1 0 38364 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2125_
timestamp 1667941163
transform 1 0 39744 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2126__78
timestamp 1667941163
transform 1 0 16836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2126_
timestamp 1667941163
transform 1 0 16744 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2127__79
timestamp 1667941163
transform 1 0 45816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2127_
timestamp 1667941163
transform 1 0 45356 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2128_
timestamp 1667941163
transform 1 0 1564 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2128__80
timestamp 1667941163
transform 1 0 2116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2129_
timestamp 1667941163
transform 1 0 1564 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2129__81
timestamp 1667941163
transform 1 0 2116 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2130__82
timestamp 1667941163
transform 1 0 7176 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2130_
timestamp 1667941163
transform 1 0 2116 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2131__83
timestamp 1667941163
transform 1 0 47748 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2131_
timestamp 1667941163
transform 1 0 46460 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2132__84
timestamp 1667941163
transform 1 0 47012 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2132_
timestamp 1667941163
transform 1 0 46460 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2133__85
timestamp 1667941163
transform 1 0 47472 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2133_
timestamp 1667941163
transform 1 0 46460 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2134__86
timestamp 1667941163
transform 1 0 16836 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2134_
timestamp 1667941163
transform 1 0 14996 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2135__87
timestamp 1667941163
transform 1 0 47748 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2135_
timestamp 1667941163
transform 1 0 46460 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2136__88
timestamp 1667941163
transform 1 0 26036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2136_
timestamp 1667941163
transform 1 0 25944 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2137__89
timestamp 1667941163
transform 1 0 39008 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2137_
timestamp 1667941163
transform 1 0 39008 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2138__90
timestamp 1667941163
transform 1 0 41216 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2138_
timestamp 1667941163
transform 1 0 42596 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2139__91
timestamp 1667941163
transform 1 0 25208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2139_
timestamp 1667941163
transform 1 0 24748 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2140__92
timestamp 1667941163
transform 1 0 45724 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2140_
timestamp 1667941163
transform 1 0 43056 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2141__93
timestamp 1667941163
transform 1 0 1840 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2141_
timestamp 1667941163
transform 1 0 2116 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2142__94
timestamp 1667941163
transform 1 0 47748 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2142_
timestamp 1667941163
transform 1 0 46460 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2143__95
timestamp 1667941163
transform 1 0 12512 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2143_
timestamp 1667941163
transform 1 0 11960 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2144__96
timestamp 1667941163
transform 1 0 3956 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2144_
timestamp 1667941163
transform 1 0 3956 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2145_
timestamp 1667941163
transform 1 0 10488 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2145__97
timestamp 1667941163
transform 1 0 10488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2146__98
timestamp 1667941163
transform 1 0 2116 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2146_
timestamp 1667941163
transform 1 0 1564 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2147__99
timestamp 1667941163
transform 1 0 47012 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2147_
timestamp 1667941163
transform 1 0 46460 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2148_
timestamp 1667941163
transform 1 0 46460 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2148__100
timestamp 1667941163
transform 1 0 47748 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2149__101
timestamp 1667941163
transform 1 0 47748 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2149_
timestamp 1667941163
transform 1 0 46460 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2150__102
timestamp 1667941163
transform 1 0 1564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2150_
timestamp 1667941163
transform 1 0 2208 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2151_
timestamp 1667941163
transform 1 0 14260 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2151__103
timestamp 1667941163
transform 1 0 13524 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2152__104
timestamp 1667941163
transform 1 0 44436 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2152_
timestamp 1667941163
transform 1 0 45356 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2153__105
timestamp 1667941163
transform 1 0 12972 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2153_
timestamp 1667941163
transform 1 0 12972 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2154__106
timestamp 1667941163
transform 1 0 35512 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2154_
timestamp 1667941163
transform 1 0 35420 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2155_
timestamp 1667941163
transform 1 0 14260 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2155__107
timestamp 1667941163
transform 1 0 14260 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2156__108
timestamp 1667941163
transform 1 0 47748 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2156_
timestamp 1667941163
transform 1 0 46460 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2157__109
timestamp 1667941163
transform 1 0 7176 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2157_
timestamp 1667941163
transform 1 0 1840 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2158__110
timestamp 1667941163
transform 1 0 4784 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2158_
timestamp 1667941163
transform 1 0 4140 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2159_
timestamp 1667941163
transform 1 0 24656 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2159__111
timestamp 1667941163
transform 1 0 23828 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2160__112
timestamp 1667941163
transform 1 0 25484 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2160_
timestamp 1667941163
transform 1 0 24748 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2161_
timestamp 1667941163
transform 1 0 45356 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2161__113
timestamp 1667941163
transform 1 0 47748 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2162__114
timestamp 1667941163
transform 1 0 47748 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2162_
timestamp 1667941163
transform 1 0 46460 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2163_
timestamp 1667941163
transform 1 0 28980 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2163__115
timestamp 1667941163
transform 1 0 28336 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2164__116
timestamp 1667941163
transform 1 0 43056 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2164_
timestamp 1667941163
transform 1 0 42596 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2165__117
timestamp 1667941163
transform 1 0 47748 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2165_
timestamp 1667941163
transform 1 0 46460 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2166__118
timestamp 1667941163
transform 1 0 3220 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2166_
timestamp 1667941163
transform 1 0 4140 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2167__119
timestamp 1667941163
transform 1 0 40756 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2167_
timestamp 1667941163
transform 1 0 40756 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2168_
timestamp 1667941163
transform 1 0 1564 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2168__120
timestamp 1667941163
transform 1 0 2024 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2169__121
timestamp 1667941163
transform 1 0 19964 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2169_
timestamp 1667941163
transform 1 0 19596 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2170__122
timestamp 1667941163
transform 1 0 10488 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2170_
timestamp 1667941163
transform 1 0 10488 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2171__123
timestamp 1667941163
transform 1 0 2024 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2171_
timestamp 1667941163
transform 1 0 2024 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2172__124
timestamp 1667941163
transform 1 0 2024 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2172_
timestamp 1667941163
transform 1 0 2024 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _2173__125
timestamp 1667941163
transform 1 0 2024 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2173_
timestamp 1667941163
transform 1 0 2024 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i
timestamp 1667941163
transform 1 0 29716 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17940 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_wb_clk_i
timestamp 1667941163
transform 1 0 17940 0 -1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_wb_clk_i
timestamp 1667941163
transform 1 0 21988 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_wb_clk_i
timestamp 1667941163
transform 1 0 23092 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_wb_clk_i
timestamp 1667941163
transform 1 0 19412 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_wb_clk_i
timestamp 1667941163
transform 1 0 19412 0 1 39168
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_wb_clk_i
timestamp 1667941163
transform 1 0 24564 0 -1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_wb_clk_i
timestamp 1667941163
transform 1 0 25668 0 1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_wb_clk_i
timestamp 1667941163
transform 1 0 32476 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_wb_clk_i
timestamp 1667941163
transform 1 0 32936 0 1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_wb_clk_i
timestamp 1667941163
transform 1 0 40112 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_wb_clk_i
timestamp 1667941163
transform 1 0 40020 0 1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_wb_clk_i
timestamp 1667941163
transform 1 0 33304 0 1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_wb_clk_i
timestamp 1667941163
transform 1 0 31924 0 1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_wb_clk_i
timestamp 1667941163
transform 1 0 36524 0 1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_wb_clk_i
timestamp 1667941163
transform 1 0 35880 0 -1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  fanout26
timestamp 1667941163
transform 1 0 7820 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14260 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout28
timestamp 1667941163
transform 1 0 20240 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1667941163
transform 1 0 1564 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 1667941163
transform 1 0 9108 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  input3
timestamp 1667941163
transform 1 0 47840 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1667941163
transform 1 0 32292 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input5
timestamp 1667941163
transform 1 0 24564 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input6
timestamp 1667941163
transform 1 0 43884 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input7
timestamp 1667941163
transform 1 0 17480 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input8
timestamp 1667941163
transform 1 0 20056 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1667941163
transform 1 0 1564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input10
timestamp 1667941163
transform 1 0 47840 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input11
timestamp 1667941163
transform 1 0 47840 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input12
timestamp 1667941163
transform 1 0 2484 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input13
timestamp 1667941163
transform 1 0 14260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input14
timestamp 1667941163
transform 1 0 1564 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1667941163
transform 1 0 48024 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1667941163
transform 1 0 1564 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1667941163
transform 1 0 1564 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input19
timestamp 1667941163
transform 1 0 11684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input20
timestamp 1667941163
transform 1 0 1564 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1667941163
transform 1 0 38732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1667941163
transform 1 0 1564 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input23
timestamp 1667941163
transform 1 0 42596 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1667941163
transform 1 0 48024 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1667941163
transform 1 0 19412 0 1 46784
box -38 -48 406 592
<< labels >>
flabel metal3 s 200 46188 800 46428 0 FreeSans 960 0 0 0 active
port 0 nsew signal input
flabel metal2 s 15446 200 15558 800 0 FreeSans 448 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 27682 49200 27794 49800 0 FreeSans 448 90 0 0 io_in[10]
port 2 nsew signal input
flabel metal2 s -10 49200 102 49800 0 FreeSans 448 90 0 0 io_in[11]
port 3 nsew signal input
flabel metal3 s 49200 42108 49800 42348 0 FreeSans 960 0 0 0 io_in[12]
port 4 nsew signal input
flabel metal2 s 23818 200 23930 800 0 FreeSans 448 90 0 0 io_in[13]
port 5 nsew signal input
flabel metal2 s 18666 49200 18778 49800 0 FreeSans 448 90 0 0 io_in[14]
port 6 nsew signal input
flabel metal3 s 49200 44148 49800 44388 0 FreeSans 960 0 0 0 io_in[15]
port 7 nsew signal input
flabel metal3 s 49200 4028 49800 4268 0 FreeSans 960 0 0 0 io_in[16]
port 8 nsew signal input
flabel metal2 s 10294 49200 10406 49800 0 FreeSans 448 90 0 0 io_in[17]
port 9 nsew signal input
flabel metal2 s 12226 49200 12338 49800 0 FreeSans 448 90 0 0 io_in[18]
port 10 nsew signal input
flabel metal2 s 43138 200 43250 800 0 FreeSans 448 90 0 0 io_in[19]
port 11 nsew signal input
flabel metal3 s 200 16268 800 16508 0 FreeSans 960 0 0 0 io_in[1]
port 12 nsew signal input
flabel metal3 s 200 29188 800 29428 0 FreeSans 960 0 0 0 io_in[20]
port 13 nsew signal input
flabel metal3 s 200 18988 800 19228 0 FreeSans 960 0 0 0 io_in[21]
port 14 nsew signal input
flabel metal3 s 49200 15588 49800 15828 0 FreeSans 960 0 0 0 io_in[22]
port 15 nsew signal input
flabel metal2 s 9006 49200 9118 49800 0 FreeSans 448 90 0 0 io_in[23]
port 16 nsew signal input
flabel metal2 s 6430 49200 6542 49800 0 FreeSans 448 90 0 0 io_in[24]
port 17 nsew signal input
flabel metal2 s 37342 200 37454 800 0 FreeSans 448 90 0 0 io_in[25]
port 18 nsew signal input
flabel metal2 s 36698 200 36810 800 0 FreeSans 448 90 0 0 io_in[26]
port 19 nsew signal input
flabel metal3 s 49200 10828 49800 11068 0 FreeSans 960 0 0 0 io_in[27]
port 20 nsew signal input
flabel metal2 s 32834 200 32946 800 0 FreeSans 448 90 0 0 io_in[28]
port 21 nsew signal input
flabel metal2 s 49578 49200 49690 49800 0 FreeSans 448 90 0 0 io_in[29]
port 22 nsew signal input
flabel metal2 s 16090 200 16202 800 0 FreeSans 448 90 0 0 io_in[2]
port 23 nsew signal input
flabel metal3 s 49200 19668 49800 19908 0 FreeSans 960 0 0 0 io_in[30]
port 24 nsew signal input
flabel metal3 s 200 44148 800 44388 0 FreeSans 960 0 0 0 io_in[31]
port 25 nsew signal input
flabel metal2 s 30902 200 31014 800 0 FreeSans 448 90 0 0 io_in[32]
port 26 nsew signal input
flabel metal3 s 200 25788 800 26028 0 FreeSans 960 0 0 0 io_in[33]
port 27 nsew signal input
flabel metal2 s 37986 49200 38098 49800 0 FreeSans 448 90 0 0 io_in[34]
port 28 nsew signal input
flabel metal2 s 43138 49200 43250 49800 0 FreeSans 448 90 0 0 io_in[35]
port 29 nsew signal input
flabel metal3 s 49200 31228 49800 31468 0 FreeSans 960 0 0 0 io_in[36]
port 30 nsew signal input
flabel metal2 s 44426 49200 44538 49800 0 FreeSans 448 90 0 0 io_in[37]
port 31 nsew signal input
flabel metal2 s 28970 49200 29082 49800 0 FreeSans 448 90 0 0 io_in[3]
port 32 nsew signal input
flabel metal3 s 49200 30548 49800 30788 0 FreeSans 960 0 0 0 io_in[4]
port 33 nsew signal input
flabel metal3 s 49200 48228 49800 48468 0 FreeSans 960 0 0 0 io_in[5]
port 34 nsew signal input
flabel metal3 s 200 30548 800 30788 0 FreeSans 960 0 0 0 io_in[6]
port 35 nsew signal input
flabel metal3 s 200 21028 800 21268 0 FreeSans 960 0 0 0 io_in[7]
port 36 nsew signal input
flabel metal3 s 49200 33268 49800 33508 0 FreeSans 960 0 0 0 io_in[8]
port 37 nsew signal input
flabel metal2 s 8362 49200 8474 49800 0 FreeSans 448 90 0 0 io_in[9]
port 38 nsew signal input
flabel metal2 s 26394 200 26506 800 0 FreeSans 448 90 0 0 io_oeb[0]
port 39 nsew signal bidirectional
flabel metal3 s 200 16948 800 17188 0 FreeSans 960 0 0 0 io_oeb[10]
port 40 nsew signal bidirectional
flabel metal3 s 49200 28508 49800 28748 0 FreeSans 960 0 0 0 io_oeb[11]
port 41 nsew signal bidirectional
flabel metal3 s 49200 14908 49800 15148 0 FreeSans 960 0 0 0 io_oeb[12]
port 42 nsew signal bidirectional
flabel metal3 s 49200 13548 49800 13788 0 FreeSans 960 0 0 0 io_oeb[13]
port 43 nsew signal bidirectional
flabel metal3 s 200 4708 800 4948 0 FreeSans 960 0 0 0 io_oeb[14]
port 44 nsew signal bidirectional
flabel metal2 s 14158 49200 14270 49800 0 FreeSans 448 90 0 0 io_oeb[15]
port 45 nsew signal bidirectional
flabel metal3 s 49200 1988 49800 2228 0 FreeSans 960 0 0 0 io_oeb[16]
port 46 nsew signal bidirectional
flabel metal2 s 13514 200 13626 800 0 FreeSans 448 90 0 0 io_oeb[17]
port 47 nsew signal bidirectional
flabel metal2 s 36054 49200 36166 49800 0 FreeSans 448 90 0 0 io_oeb[18]
port 48 nsew signal bidirectional
flabel metal2 s 14802 49200 14914 49800 0 FreeSans 448 90 0 0 io_oeb[19]
port 49 nsew signal bidirectional
flabel metal2 s 39274 200 39386 800 0 FreeSans 448 90 0 0 io_oeb[1]
port 50 nsew signal bidirectional
flabel metal3 s 49200 21708 49800 21948 0 FreeSans 960 0 0 0 io_oeb[20]
port 51 nsew signal bidirectional
flabel metal2 s 1922 49200 2034 49800 0 FreeSans 448 90 0 0 io_oeb[21]
port 52 nsew signal bidirectional
flabel metal2 s 5142 200 5254 800 0 FreeSans 448 90 0 0 io_oeb[22]
port 53 nsew signal bidirectional
flabel metal2 s 25106 49200 25218 49800 0 FreeSans 448 90 0 0 io_oeb[23]
port 54 nsew signal bidirectional
flabel metal2 s 25750 49200 25862 49800 0 FreeSans 448 90 0 0 io_oeb[24]
port 55 nsew signal bidirectional
flabel metal2 s 47646 200 47758 800 0 FreeSans 448 90 0 0 io_oeb[25]
port 56 nsew signal bidirectional
flabel metal3 s 49200 39388 49800 39628 0 FreeSans 960 0 0 0 io_oeb[26]
port 57 nsew signal bidirectional
flabel metal2 s 29614 49200 29726 49800 0 FreeSans 448 90 0 0 io_oeb[27]
port 58 nsew signal bidirectional
flabel metal2 s 41850 200 41962 800 0 FreeSans 448 90 0 0 io_oeb[28]
port 59 nsew signal bidirectional
flabel metal3 s 49200 32588 49800 32828 0 FreeSans 960 0 0 0 io_oeb[29]
port 60 nsew signal bidirectional
flabel metal2 s 41850 49200 41962 49800 0 FreeSans 448 90 0 0 io_oeb[2]
port 61 nsew signal bidirectional
flabel metal2 s 2566 49200 2678 49800 0 FreeSans 448 90 0 0 io_oeb[30]
port 62 nsew signal bidirectional
flabel metal2 s 41206 200 41318 800 0 FreeSans 448 90 0 0 io_oeb[31]
port 63 nsew signal bidirectional
flabel metal3 s 200 25108 800 25348 0 FreeSans 960 0 0 0 io_oeb[32]
port 64 nsew signal bidirectional
flabel metal2 s 48934 200 49046 800 0 FreeSans 448 90 0 0 io_oeb[33]
port 65 nsew signal bidirectional
flabel metal2 s 10938 49200 11050 49800 0 FreeSans 448 90 0 0 io_oeb[34]
port 66 nsew signal bidirectional
flabel metal3 s 200 21708 800 21948 0 FreeSans 960 0 0 0 io_oeb[35]
port 67 nsew signal bidirectional
flabel metal3 s 200 11508 800 11748 0 FreeSans 960 0 0 0 io_oeb[36]
port 68 nsew signal bidirectional
flabel metal3 s 200 18308 800 18548 0 FreeSans 960 0 0 0 io_oeb[37]
port 69 nsew signal bidirectional
flabel metal2 s 25750 200 25862 800 0 FreeSans 448 90 0 0 io_oeb[3]
port 70 nsew signal bidirectional
flabel metal3 s 49200 -52 49800 188 0 FreeSans 960 0 0 0 io_oeb[4]
port 71 nsew signal bidirectional
flabel metal3 s 200 32588 800 32828 0 FreeSans 960 0 0 0 io_oeb[5]
port 72 nsew signal bidirectional
flabel metal3 s 49200 17628 49800 17868 0 FreeSans 960 0 0 0 io_oeb[6]
port 73 nsew signal bidirectional
flabel metal2 s 12870 49200 12982 49800 0 FreeSans 448 90 0 0 io_oeb[7]
port 74 nsew signal bidirectional
flabel metal2 s 4498 200 4610 800 0 FreeSans 448 90 0 0 io_oeb[8]
port 75 nsew signal bidirectional
flabel metal2 s 10938 200 11050 800 0 FreeSans 448 90 0 0 io_oeb[9]
port 76 nsew signal bidirectional
flabel metal3 s 49200 46868 49800 47108 0 FreeSans 960 0 0 0 io_out[0]
port 77 nsew signal bidirectional
flabel metal3 s 49200 27828 49800 28068 0 FreeSans 960 0 0 0 io_out[10]
port 78 nsew signal bidirectional
flabel metal3 s 200 2668 800 2908 0 FreeSans 960 0 0 0 io_out[11]
port 79 nsew signal bidirectional
flabel metal3 s 200 7428 800 7668 0 FreeSans 960 0 0 0 io_out[12]
port 80 nsew signal bidirectional
flabel metal2 s 40562 200 40674 800 0 FreeSans 448 90 0 0 io_out[13]
port 81 nsew signal bidirectional
flabel metal3 s 49200 40068 49800 40308 0 FreeSans 960 0 0 0 io_out[14]
port 82 nsew signal bidirectional
flabel metal3 s 200 41428 800 41668 0 FreeSans 960 0 0 0 io_out[15]
port 83 nsew signal bidirectional
flabel metal3 s 49200 26468 49800 26708 0 FreeSans 960 0 0 0 io_out[16]
port 84 nsew signal bidirectional
flabel metal2 s 46358 49200 46470 49800 0 FreeSans 448 90 0 0 io_out[17]
port 85 nsew signal bidirectional
flabel metal2 s 47002 200 47114 800 0 FreeSans 448 90 0 0 io_out[18]
port 86 nsew signal bidirectional
flabel metal3 s 200 23748 800 23988 0 FreeSans 960 0 0 0 io_out[19]
port 87 nsew signal bidirectional
flabel metal2 s 33478 49200 33590 49800 0 FreeSans 448 90 0 0 io_out[1]
port 88 nsew signal bidirectional
flabel metal2 s 40562 49200 40674 49800 0 FreeSans 448 90 0 0 io_out[20]
port 89 nsew signal bidirectional
flabel metal3 s 200 40748 800 40988 0 FreeSans 960 0 0 0 io_out[21]
port 90 nsew signal bidirectional
flabel metal2 s 32190 200 32302 800 0 FreeSans 448 90 0 0 io_out[22]
port 91 nsew signal bidirectional
flabel metal3 s 49200 22388 49800 22628 0 FreeSans 960 0 0 0 io_out[23]
port 92 nsew signal bidirectional
flabel metal2 s 27682 200 27794 800 0 FreeSans 448 90 0 0 io_out[24]
port 93 nsew signal bidirectional
flabel metal2 s 36698 49200 36810 49800 0 FreeSans 448 90 0 0 io_out[25]
port 94 nsew signal bidirectional
flabel metal3 s 200 5388 800 5628 0 FreeSans 960 0 0 0 io_out[26]
port 95 nsew signal bidirectional
flabel metal2 s 38630 49200 38742 49800 0 FreeSans 448 90 0 0 io_out[27]
port 96 nsew signal bidirectional
flabel metal2 s 17378 200 17490 800 0 FreeSans 448 90 0 0 io_out[28]
port 97 nsew signal bidirectional
flabel metal3 s 49200 1308 49800 1548 0 FreeSans 960 0 0 0 io_out[29]
port 98 nsew signal bidirectional
flabel metal2 s 7074 200 7186 800 0 FreeSans 448 90 0 0 io_out[2]
port 99 nsew signal bidirectional
flabel metal3 s 200 6748 800 6988 0 FreeSans 960 0 0 0 io_out[30]
port 100 nsew signal bidirectional
flabel metal3 s 200 14228 800 14468 0 FreeSans 960 0 0 0 io_out[31]
port 101 nsew signal bidirectional
flabel metal3 s 200 47548 800 47788 0 FreeSans 960 0 0 0 io_out[32]
port 102 nsew signal bidirectional
flabel metal3 s 49200 6748 49800 6988 0 FreeSans 960 0 0 0 io_out[33]
port 103 nsew signal bidirectional
flabel metal3 s 49200 41428 49800 41668 0 FreeSans 960 0 0 0 io_out[34]
port 104 nsew signal bidirectional
flabel metal3 s 49200 38028 49800 38268 0 FreeSans 960 0 0 0 io_out[35]
port 105 nsew signal bidirectional
flabel metal2 s 15446 49200 15558 49800 0 FreeSans 448 90 0 0 io_out[36]
port 106 nsew signal bidirectional
flabel metal3 s 49200 44828 49800 45068 0 FreeSans 960 0 0 0 io_out[37]
port 107 nsew signal bidirectional
flabel metal3 s 200 43468 800 43708 0 FreeSans 960 0 0 0 io_out[3]
port 108 nsew signal bidirectional
flabel metal3 s 49200 29188 49800 29428 0 FreeSans 960 0 0 0 io_out[4]
port 109 nsew signal bidirectional
flabel metal2 s 23174 49200 23286 49800 0 FreeSans 448 90 0 0 io_out[5]
port 110 nsew signal bidirectional
flabel metal2 s 48290 49200 48402 49800 0 FreeSans 448 90 0 0 io_out[6]
port 111 nsew signal bidirectional
flabel metal3 s 200 20348 800 20588 0 FreeSans 960 0 0 0 io_out[7]
port 112 nsew signal bidirectional
flabel metal2 s 19310 200 19422 800 0 FreeSans 448 90 0 0 io_out[8]
port 113 nsew signal bidirectional
flabel metal3 s 200 14908 800 15148 0 FreeSans 960 0 0 0 io_out[9]
port 114 nsew signal bidirectional
flabel metal3 s 49200 8108 49800 8348 0 FreeSans 960 0 0 0 la1_data_in[0]
port 115 nsew signal input
flabel metal2 s 21886 200 21998 800 0 FreeSans 448 90 0 0 la1_data_in[10]
port 116 nsew signal input
flabel metal3 s 49200 6068 49800 6308 0 FreeSans 960 0 0 0 la1_data_in[11]
port 117 nsew signal input
flabel metal3 s 200 37348 800 37588 0 FreeSans 960 0 0 0 la1_data_in[12]
port 118 nsew signal input
flabel metal2 s 34122 200 34234 800 0 FreeSans 448 90 0 0 la1_data_in[13]
port 119 nsew signal input
flabel metal3 s 200 13548 800 13788 0 FreeSans 960 0 0 0 la1_data_in[14]
port 120 nsew signal input
flabel metal2 s 16734 49200 16846 49800 0 FreeSans 448 90 0 0 la1_data_in[15]
port 121 nsew signal input
flabel metal2 s 31546 49200 31658 49800 0 FreeSans 448 90 0 0 la1_data_in[16]
port 122 nsew signal input
flabel metal2 s 23818 49200 23930 49800 0 FreeSans 448 90 0 0 la1_data_in[17]
port 123 nsew signal input
flabel metal2 s 43782 200 43894 800 0 FreeSans 448 90 0 0 la1_data_in[18]
port 124 nsew signal input
flabel metal2 s 17378 49200 17490 49800 0 FreeSans 448 90 0 0 la1_data_in[19]
port 125 nsew signal input
flabel metal2 s 19954 200 20066 800 0 FreeSans 448 90 0 0 la1_data_in[1]
port 126 nsew signal input
flabel metal3 s 200 36668 800 36908 0 FreeSans 960 0 0 0 la1_data_in[20]
port 127 nsew signal input
flabel metal2 s 48934 49200 49046 49800 0 FreeSans 448 90 0 0 la1_data_in[21]
port 128 nsew signal input
flabel metal3 s 49200 8788 49800 9028 0 FreeSans 960 0 0 0 la1_data_in[22]
port 129 nsew signal input
flabel metal3 s 200 628 800 868 0 FreeSans 960 0 0 0 la1_data_in[23]
port 130 nsew signal input
flabel metal2 s 14158 200 14270 800 0 FreeSans 448 90 0 0 la1_data_in[24]
port 131 nsew signal input
flabel metal3 s 200 38708 800 38948 0 FreeSans 960 0 0 0 la1_data_in[25]
port 132 nsew signal input
flabel metal3 s 49200 3348 49800 3588 0 FreeSans 960 0 0 0 la1_data_in[26]
port 133 nsew signal input
flabel metal2 s 28970 200 29082 800 0 FreeSans 448 90 0 0 la1_data_in[27]
port 134 nsew signal input
flabel metal3 s 200 33948 800 34188 0 FreeSans 960 0 0 0 la1_data_in[28]
port 135 nsew signal input
flabel metal2 s 1278 49200 1390 49800 0 FreeSans 448 90 0 0 la1_data_in[29]
port 136 nsew signal input
flabel metal2 s 11582 200 11694 800 0 FreeSans 448 90 0 0 la1_data_in[2]
port 137 nsew signal input
flabel metal2 s 1278 200 1390 800 0 FreeSans 448 90 0 0 la1_data_in[30]
port 138 nsew signal input
flabel metal2 s 38630 200 38742 800 0 FreeSans 448 90 0 0 la1_data_in[31]
port 139 nsew signal input
flabel metal3 s 200 31908 800 32148 0 FreeSans 960 0 0 0 la1_data_in[3]
port 140 nsew signal input
flabel metal2 s 42494 49200 42606 49800 0 FreeSans 448 90 0 0 la1_data_in[4]
port 141 nsew signal input
flabel metal3 s 49200 24428 49800 24668 0 FreeSans 960 0 0 0 la1_data_in[5]
port 142 nsew signal input
flabel metal2 s 19310 49200 19422 49800 0 FreeSans 448 90 0 0 la1_data_in[6]
port 143 nsew signal input
flabel metal3 s 200 23068 800 23308 0 FreeSans 960 0 0 0 la1_data_in[7]
port 144 nsew signal input
flabel metal2 s 20598 49200 20710 49800 0 FreeSans 448 90 0 0 la1_data_in[8]
port 145 nsew signal input
flabel metal3 s 200 34628 800 34868 0 FreeSans 960 0 0 0 la1_data_in[9]
port 146 nsew signal input
flabel metal2 s 7718 200 7830 800 0 FreeSans 448 90 0 0 la1_data_out[0]
port 147 nsew signal bidirectional
flabel metal3 s 49200 12188 49800 12428 0 FreeSans 960 0 0 0 la1_data_out[10]
port 148 nsew signal bidirectional
flabel metal2 s 22530 200 22642 800 0 FreeSans 448 90 0 0 la1_data_out[11]
port 149 nsew signal bidirectional
flabel metal3 s 49200 46188 49800 46428 0 FreeSans 960 0 0 0 la1_data_out[12]
port 150 nsew signal bidirectional
flabel metal2 s 4498 49200 4610 49800 0 FreeSans 448 90 0 0 la1_data_out[13]
port 151 nsew signal bidirectional
flabel metal2 s 27038 49200 27150 49800 0 FreeSans 448 90 0 0 la1_data_out[14]
port 152 nsew signal bidirectional
flabel metal3 s 200 1308 800 1548 0 FreeSans 960 0 0 0 la1_data_out[15]
port 153 nsew signal bidirectional
flabel metal3 s 49200 16948 49800 17188 0 FreeSans 960 0 0 0 la1_data_out[16]
port 154 nsew signal bidirectional
flabel metal3 s 49200 35988 49800 36228 0 FreeSans 960 0 0 0 la1_data_out[17]
port 155 nsew signal bidirectional
flabel metal2 s 5786 49200 5898 49800 0 FreeSans 448 90 0 0 la1_data_out[18]
port 156 nsew signal bidirectional
flabel metal3 s 49200 25788 49800 26028 0 FreeSans 960 0 0 0 la1_data_out[19]
port 157 nsew signal bidirectional
flabel metal3 s 200 45508 800 45748 0 FreeSans 960 0 0 0 la1_data_out[1]
port 158 nsew signal bidirectional
flabel metal3 s 200 10148 800 10388 0 FreeSans 960 0 0 0 la1_data_out[20]
port 159 nsew signal bidirectional
flabel metal3 s 49200 42788 49800 43028 0 FreeSans 960 0 0 0 la1_data_out[21]
port 160 nsew signal bidirectional
flabel metal2 s 30258 49200 30370 49800 0 FreeSans 448 90 0 0 la1_data_out[22]
port 161 nsew signal bidirectional
flabel metal2 s 12870 200 12982 800 0 FreeSans 448 90 0 0 la1_data_out[23]
port 162 nsew signal bidirectional
flabel metal3 s 49200 18988 49800 19228 0 FreeSans 960 0 0 0 la1_data_out[24]
port 163 nsew signal bidirectional
flabel metal3 s 200 3348 800 3588 0 FreeSans 960 0 0 0 la1_data_out[25]
port 164 nsew signal bidirectional
flabel metal3 s 49200 5388 49800 5628 0 FreeSans 960 0 0 0 la1_data_out[26]
port 165 nsew signal bidirectional
flabel metal3 s 200 48228 800 48468 0 FreeSans 960 0 0 0 la1_data_out[27]
port 166 nsew signal bidirectional
flabel metal2 s 45070 200 45182 800 0 FreeSans 448 90 0 0 la1_data_out[28]
port 167 nsew signal bidirectional
flabel metal2 s 6430 200 6542 800 0 FreeSans 448 90 0 0 la1_data_out[29]
port 168 nsew signal bidirectional
flabel metal2 s 20598 200 20710 800 0 FreeSans 448 90 0 0 la1_data_out[2]
port 169 nsew signal bidirectional
flabel metal3 s 49200 12868 49800 13108 0 FreeSans 960 0 0 0 la1_data_out[30]
port 170 nsew signal bidirectional
flabel metal3 s 49200 48908 49800 49148 0 FreeSans 960 0 0 0 la1_data_out[31]
port 171 nsew signal bidirectional
flabel metal3 s 200 9468 800 9708 0 FreeSans 960 0 0 0 la1_data_out[3]
port 172 nsew signal bidirectional
flabel metal2 s 45714 200 45826 800 0 FreeSans 448 90 0 0 la1_data_out[4]
port 173 nsew signal bidirectional
flabel metal2 s 3210 200 3322 800 0 FreeSans 448 90 0 0 la1_data_out[5]
port 174 nsew signal bidirectional
flabel metal3 s 49200 20348 49800 20588 0 FreeSans 960 0 0 0 la1_data_out[6]
port 175 nsew signal bidirectional
flabel metal2 s 634 200 746 800 0 FreeSans 448 90 0 0 la1_data_out[7]
port 176 nsew signal bidirectional
flabel metal3 s 49200 37348 49800 37588 0 FreeSans 960 0 0 0 la1_data_out[8]
port 177 nsew signal bidirectional
flabel metal2 s 47002 49200 47114 49800 0 FreeSans 448 90 0 0 la1_data_out[9]
port 178 nsew signal bidirectional
flabel metal2 s 49578 200 49690 800 0 FreeSans 448 90 0 0 la1_oenb[0]
port 179 nsew signal input
flabel metal2 s 45070 49200 45182 49800 0 FreeSans 448 90 0 0 la1_oenb[10]
port 180 nsew signal input
flabel metal3 s 200 27828 800 28068 0 FreeSans 960 0 0 0 la1_oenb[11]
port 181 nsew signal input
flabel metal3 s 200 29868 800 30108 0 FreeSans 960 0 0 0 la1_oenb[12]
port 182 nsew signal input
flabel metal2 s 30258 200 30370 800 0 FreeSans 448 90 0 0 la1_oenb[13]
port 183 nsew signal input
flabel metal2 s -10 200 102 800 0 FreeSans 448 90 0 0 la1_oenb[14]
port 184 nsew signal input
flabel metal2 s 35410 200 35522 800 0 FreeSans 448 90 0 0 la1_oenb[15]
port 185 nsew signal input
flabel metal3 s 200 35988 800 36228 0 FreeSans 960 0 0 0 la1_oenb[16]
port 186 nsew signal input
flabel metal2 s 3854 49200 3966 49800 0 FreeSans 448 90 0 0 la1_oenb[17]
port 187 nsew signal input
flabel metal2 s 21886 49200 21998 49800 0 FreeSans 448 90 0 0 la1_oenb[18]
port 188 nsew signal input
flabel metal3 s 200 27148 800 27388 0 FreeSans 960 0 0 0 la1_oenb[19]
port 189 nsew signal input
flabel metal2 s 9006 200 9118 800 0 FreeSans 448 90 0 0 la1_oenb[1]
port 190 nsew signal input
flabel metal2 s 2566 200 2678 800 0 FreeSans 448 90 0 0 la1_oenb[20]
port 191 nsew signal input
flabel metal2 s 32190 49200 32302 49800 0 FreeSans 448 90 0 0 la1_oenb[21]
port 192 nsew signal input
flabel metal2 s 21242 49200 21354 49800 0 FreeSans 448 90 0 0 la1_oenb[22]
port 193 nsew signal input
flabel metal2 s 24462 200 24574 800 0 FreeSans 448 90 0 0 la1_oenb[23]
port 194 nsew signal input
flabel metal2 s 39918 49200 40030 49800 0 FreeSans 448 90 0 0 la1_oenb[24]
port 195 nsew signal input
flabel metal3 s 49200 10148 49800 10388 0 FreeSans 960 0 0 0 la1_oenb[25]
port 196 nsew signal input
flabel metal3 s 200 39388 800 39628 0 FreeSans 960 0 0 0 la1_oenb[26]
port 197 nsew signal input
flabel metal3 s 49200 35308 49800 35548 0 FreeSans 960 0 0 0 la1_oenb[27]
port 198 nsew signal input
flabel metal2 s 9650 200 9762 800 0 FreeSans 448 90 0 0 la1_oenb[28]
port 199 nsew signal input
flabel metal2 s 18022 200 18134 800 0 FreeSans 448 90 0 0 la1_oenb[29]
port 200 nsew signal input
flabel metal3 s 200 8108 800 8348 0 FreeSans 960 0 0 0 la1_oenb[2]
port 201 nsew signal input
flabel metal3 s 49200 34628 49800 34868 0 FreeSans 960 0 0 0 la1_oenb[30]
port 202 nsew signal input
flabel metal2 s 28326 200 28438 800 0 FreeSans 448 90 0 0 la1_oenb[31]
port 203 nsew signal input
flabel metal2 s 35410 49200 35522 49800 0 FreeSans 448 90 0 0 la1_oenb[3]
port 204 nsew signal input
flabel metal2 s 34122 49200 34234 49800 0 FreeSans 448 90 0 0 la1_oenb[4]
port 205 nsew signal input
flabel metal3 s 200 49588 800 49828 0 FreeSans 960 0 0 0 la1_oenb[5]
port 206 nsew signal input
flabel metal2 s 7718 49200 7830 49800 0 FreeSans 448 90 0 0 la1_oenb[6]
port 207 nsew signal input
flabel metal2 s 34766 200 34878 800 0 FreeSans 448 90 0 0 la1_oenb[7]
port 208 nsew signal input
flabel metal3 s 200 12188 800 12428 0 FreeSans 960 0 0 0 la1_oenb[8]
port 209 nsew signal input
flabel metal3 s 200 42788 800 43028 0 FreeSans 960 0 0 0 la1_oenb[9]
port 210 nsew signal input
flabel metal4 s 4208 2128 4528 47376 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 34928 2128 35248 47376 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 19568 2128 19888 47376 0 FreeSans 1920 90 0 0 vssd1
port 212 nsew ground bidirectional
flabel metal3 s 49200 23748 49800 23988 0 FreeSans 960 0 0 0 wb_clk_i
port 213 nsew signal input
rlabel metal1 24978 47328 24978 47328 0 vccd1
rlabel metal1 24978 46784 24978 46784 0 vssd1
rlabel metal2 15226 20434 15226 20434 0 _0000_
rlabel metal2 12466 21046 12466 21046 0 _0001_
rlabel metal2 12558 22406 12558 22406 0 _0002_
rlabel metal2 14306 22406 14306 22406 0 _0003_
rlabel metal1 15359 18734 15359 18734 0 _0004_
rlabel metal1 14807 17238 14807 17238 0 _0005_
rlabel via1 14117 15062 14117 15062 0 _0006_
rlabel metal2 12926 15878 12926 15878 0 _0007_
rlabel metal2 12098 17442 12098 17442 0 _0008_
rlabel metal1 11776 18938 11776 18938 0 _0009_
rlabel metal1 39820 24106 39820 24106 0 _0010_
rlabel via1 40337 20910 40337 20910 0 _0011_
rlabel metal1 36519 21930 36519 21930 0 _0012_
rlabel via1 33529 26962 33529 26962 0 _0013_
rlabel metal2 31602 21794 31602 21794 0 _0014_
rlabel metal1 35972 19482 35972 19482 0 _0015_
rlabel metal2 36846 16966 36846 16966 0 _0016_
rlabel metal1 35047 15062 35047 15062 0 _0017_
rlabel metal1 29118 21114 29118 21114 0 _0018_
rlabel metal2 26818 19142 26818 19142 0 _0019_
rlabel metal1 29118 14586 29118 14586 0 _0020_
rlabel metal2 23506 17000 23506 17000 0 _0021_
rlabel metal1 27876 11730 27876 11730 0 _0022_
rlabel metal1 27181 10030 27181 10030 0 _0023_
rlabel metal2 32338 11288 32338 11288 0 _0024_
rlabel via1 34173 12818 34173 12818 0 _0025_
rlabel metal1 34576 41174 34576 41174 0 _0026_
rlabel metal2 34454 42466 34454 42466 0 _0027_
rlabel metal1 30217 42262 30217 42262 0 _0028_
rlabel metal1 28929 42602 28929 42602 0 _0029_
rlabel metal2 29762 38726 29762 38726 0 _0030_
rlabel metal1 35420 38522 35420 38522 0 _0031_
rlabel metal1 34944 37162 34944 37162 0 _0032_
rlabel metal1 32011 36074 32011 36074 0 _0033_
rlabel metal2 27738 40256 27738 40256 0 _0034_
rlabel metal1 25801 42602 25801 42602 0 _0035_
rlabel metal1 21707 40426 21707 40426 0 _0036_
rlabel metal1 21891 42602 21891 42602 0 _0037_
rlabel metal1 15865 41514 15865 41514 0 _0038_
rlabel metal1 14577 41174 14577 41174 0 _0039_
rlabel metal2 19458 41990 19458 41990 0 _0040_
rlabel metal1 19085 40018 19085 40018 0 _0041_
rlabel via1 30585 34646 30585 34646 0 _0042_
rlabel metal1 32512 32402 32512 32402 0 _0043_
rlabel metal1 27600 28730 27600 28730 0 _0044_
rlabel metal1 18993 36822 18993 36822 0 _0045_
rlabel via1 12645 37230 12645 37230 0 _0046_
rlabel metal2 12834 35938 12834 35938 0 _0047_
rlabel metal1 18860 28186 18860 28186 0 _0048_
rlabel metal2 12558 27234 12558 27234 0 _0049_
rlabel metal1 19320 30090 19320 30090 0 _0050_
rlabel metal2 12466 31518 12466 31518 0 _0051_
rlabel metal1 24508 29138 24508 29138 0 _0052_
rlabel metal2 20010 27846 20010 27846 0 _0053_
rlabel metal2 22126 34918 22126 34918 0 _0054_
rlabel metal1 22678 37706 22678 37706 0 _0055_
rlabel metal2 24426 34850 24426 34850 0 _0056_
rlabel metal1 27549 37910 27549 37910 0 _0057_
rlabel metal2 32614 23970 32614 23970 0 _0058_
rlabel via1 33989 21590 33989 21590 0 _0059_
rlabel metal1 33764 22746 33764 22746 0 _0060_
rlabel metal1 31372 24922 31372 24922 0 _0061_
rlabel via1 29481 22610 29481 22610 0 _0062_
rlabel via1 30953 19822 30953 19822 0 _0063_
rlabel metal1 30390 18326 30390 18326 0 _0064_
rlabel metal1 30544 15674 30544 15674 0 _0065_
rlabel metal1 27268 24174 27268 24174 0 _0066_
rlabel metal1 22167 18666 22167 18666 0 _0067_
rlabel metal1 27360 13906 27360 13906 0 _0068_
rlabel metal1 21569 16558 21569 16558 0 _0069_
rlabel metal1 21845 12206 21845 12206 0 _0070_
rlabel viali 21109 13294 21109 13294 0 _0071_
rlabel via1 30033 13974 30033 13974 0 _0072_
rlabel via1 32609 13974 32609 13974 0 _0073_
rlabel metal2 7314 29410 7314 29410 0 _0074_
rlabel metal2 9522 30498 9522 30498 0 _0075_
rlabel metal1 7861 30702 7861 30702 0 _0076_
rlabel metal2 6026 31110 6026 31110 0 _0077_
rlabel metal1 4779 29614 4779 29614 0 _0078_
rlabel metal1 4825 28118 4825 28118 0 _0079_
rlabel metal1 5515 27030 5515 27030 0 _0080_
rlabel metal1 6067 26350 6067 26350 0 _0081_
rlabel metal2 7774 26146 7774 26146 0 _0082_
rlabel metal1 7850 27030 7850 27030 0 _0083_
rlabel metal2 37582 13702 37582 13702 0 _0084_
rlabel metal1 35553 10030 35553 10030 0 _0085_
rlabel metal1 37899 9554 37899 9554 0 _0086_
rlabel metal1 40296 9486 40296 9486 0 _0087_
rlabel metal2 45770 13702 45770 13702 0 _0088_
rlabel metal2 43102 15266 43102 15266 0 _0089_
rlabel metal1 45846 10710 45846 10710 0 _0090_
rlabel metal1 43097 9622 43097 9622 0 _0091_
rlabel metal1 40112 12954 40112 12954 0 _0092_
rlabel metal2 39330 15878 39330 15878 0 _0093_
rlabel metal1 40802 17850 40802 17850 0 _0094_
rlabel metal1 43562 16762 43562 16762 0 _0095_
rlabel metal1 43920 22610 43920 22610 0 _0096_
rlabel metal2 45218 21726 45218 21726 0 _0097_
rlabel metal1 44880 18326 44880 18326 0 _0098_
rlabel metal1 42412 18938 42412 18938 0 _0099_
rlabel metal1 20511 23018 20511 23018 0 _0100_
rlabel metal2 22402 21692 22402 21692 0 _0101_
rlabel metal1 19534 20502 19534 20502 0 _0102_
rlabel metal2 17802 21794 17802 21794 0 _0103_
rlabel metal1 16647 23018 16647 23018 0 _0104_
rlabel metal1 17751 18666 17751 18666 0 _0105_
rlabel metal1 18993 15062 18993 15062 0 _0106_
rlabel metal1 16222 14314 16222 14314 0 _0107_
rlabel metal1 16785 16490 16785 16490 0 _0108_
rlabel metal1 19085 17238 19085 17238 0 _0109_
rlabel metal2 25714 24310 25714 24310 0 _0110_
rlabel metal1 24375 21590 24375 21590 0 _0111_
rlabel metal1 39314 25942 39314 25942 0 _0112_
rlabel metal2 38594 27234 38594 27234 0 _0113_
rlabel metal2 38042 25058 38042 25058 0 _0114_
rlabel metal2 31326 26690 31326 26690 0 _0115_
rlabel metal1 29849 24854 29849 24854 0 _0116_
rlabel metal2 37766 20230 37766 20230 0 _0117_
rlabel metal1 38543 17646 38543 17646 0 _0118_
rlabel metal1 32384 16218 32384 16218 0 _0119_
rlabel metal1 27232 20570 27232 20570 0 _0120_
rlabel metal1 24145 18326 24145 18326 0 _0121_
rlabel via1 24605 13906 24605 13906 0 _0122_
rlabel metal2 23230 14994 23230 14994 0 _0123_
rlabel metal2 22494 10914 22494 10914 0 _0124_
rlabel metal2 22402 9826 22402 9826 0 _0125_
rlabel metal2 24610 10438 24610 10438 0 _0126_
rlabel metal1 25203 11050 25203 11050 0 _0127_
rlabel metal1 37566 15062 37566 15062 0 _0128_
rlabel metal2 30222 30838 30222 30838 0 _0129_
rlabel metal1 30856 28526 30856 28526 0 _0130_
rlabel metal1 27232 26010 27232 26010 0 _0131_
rlabel metal1 17935 32878 17935 32878 0 _0132_
rlabel metal1 12052 33626 12052 33626 0 _0133_
rlabel metal2 14306 33286 14306 33286 0 _0134_
rlabel metal2 17894 26146 17894 26146 0 _0135_
rlabel metal2 12374 25058 12374 25058 0 _0136_
rlabel metal1 15911 25194 15911 25194 0 _0137_
rlabel via1 12277 30226 12277 30226 0 _0138_
rlabel metal2 26174 29410 26174 29410 0 _0139_
rlabel metal1 20189 26350 20189 26350 0 _0140_
rlabel metal1 19913 33558 19913 33558 0 _0141_
rlabel metal2 20194 37094 20194 37094 0 _0142_
rlabel metal1 27360 32402 27360 32402 0 _0143_
rlabel metal1 27216 34646 27216 34646 0 _0144_
rlabel metal1 28474 36346 28474 36346 0 _0145_
rlabel metal2 29026 35190 29026 35190 0 _0146_
rlabel metal1 29200 32402 29200 32402 0 _0147_
rlabel metal1 29010 27030 29010 27030 0 _0148_
rlabel metal2 17526 38454 17526 38454 0 _0149_
rlabel metal1 15364 37978 15364 37978 0 _0150_
rlabel metal2 13938 39202 13938 39202 0 _0151_
rlabel metal1 21477 24174 21477 24174 0 _0152_
rlabel metal2 14398 24582 14398 24582 0 _0153_
rlabel via1 18441 24854 18441 24854 0 _0154_
rlabel metal2 16882 33762 16882 33762 0 _0155_
rlabel via1 24881 27370 24881 27370 0 _0156_
rlabel via1 22305 26282 22305 26282 0 _0157_
rlabel metal2 21022 31586 21022 31586 0 _0158_
rlabel metal1 22208 32402 22208 32402 0 _0159_
rlabel metal1 24554 31790 24554 31790 0 _0160_
rlabel metal2 23966 32674 23966 32674 0 _0161_
rlabel metal1 23598 19856 23598 19856 0 _0162_
rlabel metal1 23598 20434 23598 20434 0 _0163_
rlabel metal1 24242 19754 24242 19754 0 _0164_
rlabel metal1 21252 13838 21252 13838 0 _0165_
rlabel metal2 23598 18938 23598 18938 0 _0166_
rlabel metal1 32706 13260 32706 13260 0 _0167_
rlabel metal1 34132 21998 34132 21998 0 _0168_
rlabel metal1 18630 17646 18630 17646 0 _0169_
rlabel metal2 32798 24140 32798 24140 0 _0170_
rlabel metal1 32982 22032 32982 22032 0 _0171_
rlabel metal1 33764 22610 33764 22610 0 _0172_
rlabel metal1 31924 24786 31924 24786 0 _0173_
rlabel metal1 21528 32878 21528 32878 0 _0174_
rlabel metal1 22264 12818 22264 12818 0 _0175_
rlabel metal1 29670 23290 29670 23290 0 _0176_
rlabel metal2 31050 19958 31050 19958 0 _0177_
rlabel metal1 30636 17850 30636 17850 0 _0178_
rlabel metal2 30682 15674 30682 15674 0 _0179_
rlabel metal2 27554 24310 27554 24310 0 _0180_
rlabel metal1 22356 18394 22356 18394 0 _0181_
rlabel metal2 27646 13872 27646 13872 0 _0182_
rlabel metal2 22218 16694 22218 16694 0 _0183_
rlabel metal2 22862 13124 22862 13124 0 _0184_
rlabel metal1 21620 13906 21620 13906 0 _0185_
rlabel metal1 37858 20876 37858 20876 0 _0186_
rlabel metal2 30406 13872 30406 13872 0 _0187_
rlabel metal1 32476 13498 32476 13498 0 _0188_
rlabel metal1 7774 29104 7774 29104 0 _0189_
rlabel metal1 5014 27438 5014 27438 0 _0190_
rlabel metal2 7498 29614 7498 29614 0 _0191_
rlabel metal2 8694 29750 8694 29750 0 _0192_
rlabel metal1 8740 30362 8740 30362 0 _0193_
rlabel metal1 6118 30362 6118 30362 0 _0194_
rlabel metal1 5106 30260 5106 30260 0 _0195_
rlabel metal1 5428 28526 5428 28526 0 _0196_
rlabel metal1 6578 27472 6578 27472 0 _0197_
rlabel metal1 6348 26962 6348 26962 0 _0198_
rlabel metal1 7636 25874 7636 25874 0 _0199_
rlabel metal2 7590 27132 7590 27132 0 _0200_
rlabel metal1 32844 10642 32844 10642 0 _0201_
rlabel metal1 30360 10778 30360 10778 0 _0202_
rlabel metal1 36662 11084 36662 11084 0 _0203_
rlabel metal1 29854 10234 29854 10234 0 _0204_
rlabel metal1 36754 11186 36754 11186 0 _0205_
rlabel metal1 36478 12274 36478 12274 0 _0206_
rlabel metal1 38548 14382 38548 14382 0 _0207_
rlabel metal1 37398 12410 37398 12410 0 _0208_
rlabel metal2 37490 12988 37490 12988 0 _0209_
rlabel metal1 36524 12750 36524 12750 0 _0210_
rlabel metal2 36754 12988 36754 12988 0 _0211_
rlabel metal1 35650 11118 35650 11118 0 _0212_
rlabel metal2 35466 11628 35466 11628 0 _0213_
rlabel metal2 35558 10846 35558 10846 0 _0214_
rlabel metal2 39514 9350 39514 9350 0 _0215_
rlabel metal1 39376 9554 39376 9554 0 _0216_
rlabel metal2 38502 10268 38502 10268 0 _0217_
rlabel metal2 38962 14960 38962 14960 0 _0218_
rlabel metal1 38364 10778 38364 10778 0 _0219_
rlabel metal1 37766 11730 37766 11730 0 _0220_
rlabel metal1 38226 10676 38226 10676 0 _0221_
rlabel metal1 38318 10064 38318 10064 0 _0222_
rlabel metal2 38226 10268 38226 10268 0 _0223_
rlabel metal1 41998 9486 41998 9486 0 _0224_
rlabel metal2 40342 10914 40342 10914 0 _0225_
rlabel metal1 40848 9622 40848 9622 0 _0226_
rlabel metal2 40434 9996 40434 9996 0 _0227_
rlabel metal2 38686 10880 38686 10880 0 _0228_
rlabel metal2 41354 11662 41354 11662 0 _0229_
rlabel metal1 44390 13260 44390 13260 0 _0230_
rlabel metal1 44298 14450 44298 14450 0 _0231_
rlabel metal2 43194 12988 43194 12988 0 _0232_
rlabel metal1 44068 12750 44068 12750 0 _0233_
rlabel metal1 44942 12852 44942 12852 0 _0234_
rlabel metal2 45034 13090 45034 13090 0 _0235_
rlabel metal1 44252 12818 44252 12818 0 _0236_
rlabel metal1 44528 14586 44528 14586 0 _0237_
rlabel metal1 43286 14926 43286 14926 0 _0238_
rlabel metal1 43516 13702 43516 13702 0 _0239_
rlabel metal1 44620 12614 44620 12614 0 _0240_
rlabel metal1 45632 10234 45632 10234 0 _0241_
rlabel metal1 44712 9894 44712 9894 0 _0242_
rlabel metal1 44528 11730 44528 11730 0 _0243_
rlabel metal2 44206 11084 44206 11084 0 _0244_
rlabel metal1 45172 11118 45172 11118 0 _0245_
rlabel metal1 44252 10030 44252 10030 0 _0246_
rlabel metal1 43470 10132 43470 10132 0 _0247_
rlabel metal2 43562 10234 43562 10234 0 _0248_
rlabel metal2 45034 10744 45034 10744 0 _0249_
rlabel metal1 41446 12240 41446 12240 0 _0250_
rlabel metal2 43102 11526 43102 11526 0 _0251_
rlabel metal2 41170 12036 41170 12036 0 _0252_
rlabel metal1 41446 13872 41446 13872 0 _0253_
rlabel metal1 41676 13294 41676 13294 0 _0254_
rlabel metal1 41860 15470 41860 15470 0 _0255_
rlabel metal2 40342 13022 40342 13022 0 _0256_
rlabel metal2 40250 13362 40250 13362 0 _0257_
rlabel metal2 41630 15113 41630 15113 0 _0258_
rlabel metal1 42320 15946 42320 15946 0 _0259_
rlabel metal1 40342 14824 40342 14824 0 _0260_
rlabel metal2 41446 15232 41446 15232 0 _0261_
rlabel metal2 40526 15130 40526 15130 0 _0262_
rlabel metal2 43286 17306 43286 17306 0 _0263_
rlabel metal2 41630 17340 41630 17340 0 _0264_
rlabel metal2 41078 17476 41078 17476 0 _0265_
rlabel metal1 43194 17714 43194 17714 0 _0266_
rlabel metal1 43240 16558 43240 16558 0 _0267_
rlabel metal1 42972 20774 42972 20774 0 _0268_
rlabel metal1 43516 22134 43516 22134 0 _0269_
rlabel metal1 42964 21658 42964 21658 0 _0270_
rlabel metal1 43470 22406 43470 22406 0 _0271_
rlabel metal1 43838 21114 43838 21114 0 _0272_
rlabel metal1 43654 21896 43654 21896 0 _0273_
rlabel metal1 44160 19822 44160 19822 0 _0274_
rlabel metal2 44298 18938 44298 18938 0 _0275_
rlabel metal1 44114 18768 44114 18768 0 _0276_
rlabel metal2 42826 19040 42826 19040 0 _0277_
rlabel metal2 43102 18938 43102 18938 0 _0278_
rlabel metal1 22586 22678 22586 22678 0 _0279_
rlabel metal1 19320 18190 19320 18190 0 _0280_
rlabel metal2 20194 23256 20194 23256 0 _0281_
rlabel metal2 21482 23290 21482 23290 0 _0282_
rlabel metal1 20010 19414 20010 19414 0 _0283_
rlabel metal1 20930 22134 20930 22134 0 _0284_
rlabel metal1 20746 22032 20746 22032 0 _0285_
rlabel metal2 20102 19448 20102 19448 0 _0286_
rlabel metal1 20102 19482 20102 19482 0 _0287_
rlabel metal1 17526 22474 17526 22474 0 _0288_
rlabel metal1 18032 21522 18032 21522 0 _0289_
rlabel metal2 18078 23426 18078 23426 0 _0290_
rlabel metal2 17526 24004 17526 24004 0 _0291_
rlabel metal1 18722 19448 18722 19448 0 _0292_
rlabel metal2 19090 19958 19090 19958 0 _0293_
rlabel metal1 18538 15368 18538 15368 0 _0294_
rlabel metal2 18906 15878 18906 15878 0 _0295_
rlabel metal2 17158 15096 17158 15096 0 _0296_
rlabel metal1 16951 15130 16951 15130 0 _0297_
rlabel metal1 17756 16150 17756 16150 0 _0298_
rlabel metal1 17710 17170 17710 17170 0 _0299_
rlabel metal2 18722 17918 18722 17918 0 _0300_
rlabel metal1 19642 17680 19642 17680 0 _0301_
rlabel metal1 24656 20910 24656 20910 0 _0302_
rlabel metal1 25346 24174 25346 24174 0 _0303_
rlabel metal1 24886 26996 24886 26996 0 _0304_
rlabel metal2 16882 32606 16882 32606 0 _0305_
rlabel metal2 25622 24004 25622 24004 0 _0306_
rlabel metal1 24840 21114 24840 21114 0 _0307_
rlabel metal1 25070 20502 25070 20502 0 _0308_
rlabel metal1 24656 19346 24656 19346 0 _0309_
rlabel metal2 32706 18054 32706 18054 0 _0310_
rlabel metal1 23414 21522 23414 21522 0 _0311_
rlabel metal1 23690 14960 23690 14960 0 _0312_
rlabel metal2 38962 16864 38962 16864 0 _0313_
rlabel metal1 39238 26384 39238 26384 0 _0314_
rlabel metal1 38778 26928 38778 26928 0 _0315_
rlabel metal2 38226 25228 38226 25228 0 _0316_
rlabel metal2 31510 26316 31510 26316 0 _0317_
rlabel metal1 29992 24378 29992 24378 0 _0318_
rlabel metal2 37950 20298 37950 20298 0 _0319_
rlabel metal2 38502 18564 38502 18564 0 _0320_
rlabel metal2 32522 16524 32522 16524 0 _0321_
rlabel metal1 26818 22032 26818 22032 0 _0322_
rlabel metal2 27370 21148 27370 21148 0 _0323_
rlabel metal2 24794 19074 24794 19074 0 _0324_
rlabel metal1 24840 13498 24840 13498 0 _0325_
rlabel metal2 23414 14586 23414 14586 0 _0326_
rlabel metal2 22678 11084 22678 11084 0 _0327_
rlabel metal2 22586 10812 22586 10812 0 _0328_
rlabel metal2 24794 10778 24794 10778 0 _0329_
rlabel metal2 25622 11900 25622 11900 0 _0330_
rlabel metal2 23690 24786 23690 24786 0 _0331_
rlabel metal1 20608 34034 20608 34034 0 _0332_
rlabel metal1 18400 33286 18400 33286 0 _0333_
rlabel metal1 20930 32912 20930 32912 0 _0334_
rlabel metal1 18676 32402 18676 32402 0 _0335_
rlabel metal2 30406 30396 30406 30396 0 _0336_
rlabel metal1 30774 28186 30774 28186 0 _0337_
rlabel metal1 18492 32402 18492 32402 0 _0338_
rlabel metal2 27370 26044 27370 26044 0 _0339_
rlabel metal2 18262 33014 18262 33014 0 _0340_
rlabel metal1 12282 33082 12282 33082 0 _0341_
rlabel metal2 14490 33082 14490 33082 0 _0342_
rlabel metal2 18078 26180 18078 26180 0 _0343_
rlabel metal2 12558 25228 12558 25228 0 _0344_
rlabel metal2 16882 25466 16882 25466 0 _0345_
rlabel metal2 12466 30260 12466 30260 0 _0346_
rlabel metal2 26358 29580 26358 29580 0 _0347_
rlabel metal2 20562 26486 20562 26486 0 _0348_
rlabel metal1 20332 33082 20332 33082 0 _0349_
rlabel metal2 21298 36890 21298 36890 0 _0350_
rlabel metal2 20378 36618 20378 36618 0 _0351_
rlabel metal1 27094 31314 27094 31314 0 _0352_
rlabel metal1 27094 34170 27094 34170 0 _0353_
rlabel metal2 24702 23834 24702 23834 0 _0354_
rlabel metal1 24150 31994 24150 31994 0 _0355_
rlabel metal2 15594 38284 15594 38284 0 _0356_
rlabel metal2 29210 34748 29210 34748 0 _0357_
rlabel metal2 28566 32436 28566 32436 0 _0358_
rlabel metal2 28566 26962 28566 26962 0 _0359_
rlabel metal2 17710 38012 17710 38012 0 _0360_
rlabel metal2 15410 38012 15410 38012 0 _0361_
rlabel metal1 14260 38522 14260 38522 0 _0362_
rlabel metal1 21528 24922 21528 24922 0 _0363_
rlabel metal1 22218 24718 22218 24718 0 _0364_
rlabel metal1 14582 24208 14582 24208 0 _0365_
rlabel metal1 18630 25228 18630 25228 0 _0366_
rlabel metal1 16744 33082 16744 33082 0 _0367_
rlabel metal1 24518 27098 24518 27098 0 _0368_
rlabel metal2 22494 26486 22494 26486 0 _0369_
rlabel metal1 21436 32742 21436 32742 0 _0370_
rlabel metal2 22310 31484 22310 31484 0 _0371_
rlabel metal1 24242 31450 24242 31450 0 _0372_
rlabel metal1 24518 32402 24518 32402 0 _0373_
rlabel metal2 4922 44608 4922 44608 0 _0374_
rlabel metal1 6118 4114 6118 4114 0 _0375_
rlabel metal2 6302 4216 6302 4216 0 _0376_
rlabel metal2 16146 4590 16146 4590 0 _0377_
rlabel metal1 3542 43214 3542 43214 0 _0378_
rlabel metal2 1978 3332 1978 3332 0 _0379_
rlabel metal2 6578 3808 6578 3808 0 _0380_
rlabel metal1 4784 3570 4784 3570 0 _0381_
rlabel metal1 2300 17646 2300 17646 0 _0382_
rlabel metal1 5106 3672 5106 3672 0 _0383_
rlabel metal1 3542 44778 3542 44778 0 _0384_
rlabel metal1 2530 5678 2530 5678 0 _0385_
rlabel metal1 13478 18870 13478 18870 0 _0386_
rlabel metal1 14260 22134 14260 22134 0 _0387_
rlabel metal1 13984 17102 13984 17102 0 _0388_
rlabel metal1 14030 19244 14030 19244 0 _0389_
rlabel metal1 14720 19142 14720 19142 0 _0390_
rlabel metal1 13938 21454 13938 21454 0 _0391_
rlabel metal2 15410 20026 15410 20026 0 _0392_
rlabel metal1 13248 20434 13248 20434 0 _0393_
rlabel metal2 12834 21556 12834 21556 0 _0394_
rlabel metal2 13938 21828 13938 21828 0 _0395_
rlabel metal1 16008 19822 16008 19822 0 _0396_
rlabel metal2 15226 17850 15226 17850 0 _0397_
rlabel metal1 14168 15470 14168 15470 0 _0398_
rlabel metal2 13110 15674 13110 15674 0 _0399_
rlabel metal2 12742 16966 12742 16966 0 _0400_
rlabel metal2 12282 18564 12282 18564 0 _0401_
rlabel metal1 9476 27914 9476 27914 0 _0402_
rlabel metal1 10396 20366 10396 20366 0 _0403_
rlabel metal1 40526 23290 40526 23290 0 _0404_
rlabel metal1 40526 23834 40526 23834 0 _0405_
rlabel metal1 40066 19822 40066 19822 0 _0406_
rlabel metal2 39422 24004 39422 24004 0 _0407_
rlabel metal2 26174 21386 26174 21386 0 _0408_
rlabel metal1 40710 20434 40710 20434 0 _0409_
rlabel metal1 40986 12716 40986 12716 0 _0410_
rlabel metal1 39974 22678 39974 22678 0 _0411_
rlabel metal2 39330 22406 39330 22406 0 _0412_
rlabel metal1 40250 22406 40250 22406 0 _0413_
rlabel metal2 40986 21726 40986 21726 0 _0414_
rlabel via1 40258 21930 40258 21930 0 _0415_
rlabel metal1 39563 21522 39563 21522 0 _0416_
rlabel metal1 40572 20026 40572 20026 0 _0417_
rlabel metal2 26174 16966 26174 16966 0 _0418_
rlabel metal1 35098 22066 35098 22066 0 _0419_
rlabel metal1 39468 22202 39468 22202 0 _0420_
rlabel metal1 37306 22984 37306 22984 0 _0421_
rlabel metal2 36386 24378 36386 24378 0 _0422_
rlabel metal2 36018 25534 36018 25534 0 _0423_
rlabel metal2 36478 23358 36478 23358 0 _0424_
rlabel metal2 36570 23290 36570 23290 0 _0425_
rlabel metal1 37076 23086 37076 23086 0 _0426_
rlabel metal1 37720 16558 37720 16558 0 _0427_
rlabel metal1 35466 19346 35466 19346 0 _0428_
rlabel metal2 35834 22780 35834 22780 0 _0429_
rlabel via1 36210 25942 36210 25942 0 _0430_
rlabel metal1 35880 27098 35880 27098 0 _0431_
rlabel metal1 35466 26350 35466 26350 0 _0432_
rlabel metal1 35788 24786 35788 24786 0 _0433_
rlabel metal1 35328 26010 35328 26010 0 _0434_
rlabel metal1 34362 26010 34362 26010 0 _0435_
rlabel metal1 33580 26010 33580 26010 0 _0436_
rlabel metal1 33442 19822 33442 19822 0 _0437_
rlabel metal2 32706 21658 32706 21658 0 _0438_
rlabel metal1 33350 20842 33350 20842 0 _0439_
rlabel metal2 36478 26350 36478 26350 0 _0440_
rlabel metal2 36938 25466 36938 25466 0 _0441_
rlabel metal1 33948 20910 33948 20910 0 _0442_
rlabel metal1 33488 20570 33488 20570 0 _0443_
rlabel metal1 33672 21114 33672 21114 0 _0444_
rlabel metal1 30866 21454 30866 21454 0 _0445_
rlabel metal1 35098 19788 35098 19788 0 _0446_
rlabel metal2 36662 18768 36662 18768 0 _0447_
rlabel metal1 35098 18768 35098 18768 0 _0448_
rlabel metal1 35328 19890 35328 19890 0 _0449_
rlabel metal2 35374 19516 35374 19516 0 _0450_
rlabel metal1 35190 19380 35190 19380 0 _0451_
rlabel metal1 35650 17748 35650 17748 0 _0452_
rlabel metal1 35098 17646 35098 17646 0 _0453_
rlabel metal2 36662 17306 36662 17306 0 _0454_
rlabel metal2 36754 17136 36754 17136 0 _0455_
rlabel metal1 37122 16626 37122 16626 0 _0456_
rlabel via1 40723 9554 40723 9554 0 _0457_
rlabel metal1 35420 16762 35420 16762 0 _0458_
rlabel metal1 34776 16558 34776 16558 0 _0459_
rlabel metal1 35157 16218 35157 16218 0 _0460_
rlabel metal1 34868 16082 34868 16082 0 _0461_
rlabel metal1 35374 15878 35374 15878 0 _0462_
rlabel metal1 35098 15504 35098 15504 0 _0463_
rlabel metal1 34086 15470 34086 15470 0 _0464_
rlabel metal2 33718 17884 33718 17884 0 _0465_
rlabel metal2 33166 18496 33166 18496 0 _0466_
rlabel metal2 33902 19482 33902 19482 0 _0467_
rlabel metal2 33994 18326 33994 18326 0 _0468_
rlabel metal1 33902 17272 33902 17272 0 _0469_
rlabel viali 34025 18292 34025 18292 0 _0470_
rlabel metal2 34178 18530 34178 18530 0 _0471_
rlabel metal1 29532 20570 29532 20570 0 _0472_
rlabel metal1 29670 20400 29670 20400 0 _0473_
rlabel metal2 29394 19788 29394 19788 0 _0474_
rlabel metal2 29486 19584 29486 19584 0 _0475_
rlabel metal1 28842 19482 28842 19482 0 _0476_
rlabel metal1 28244 20026 28244 20026 0 _0477_
rlabel metal2 28290 18564 28290 18564 0 _0478_
rlabel via1 27554 18938 27554 18938 0 _0479_
rlabel metal1 27830 18700 27830 18700 0 _0480_
rlabel metal1 28888 18938 28888 18938 0 _0481_
rlabel metal2 28106 18564 28106 18564 0 _0482_
rlabel metal1 26082 18802 26082 18802 0 _0483_
rlabel metal1 26910 14586 26910 14586 0 _0484_
rlabel metal1 27830 16014 27830 16014 0 _0485_
rlabel metal1 27738 15436 27738 15436 0 _0486_
rlabel metal1 28014 18224 28014 18224 0 _0487_
rlabel metal2 27278 17306 27278 17306 0 _0488_
rlabel metal1 28336 15470 28336 15470 0 _0489_
rlabel metal2 28566 14858 28566 14858 0 _0490_
rlabel metal2 26450 15674 26450 15674 0 _0491_
rlabel metal1 26266 15504 26266 15504 0 _0492_
rlabel metal2 26266 15878 26266 15878 0 _0493_
rlabel metal2 25990 16320 25990 16320 0 _0494_
rlabel metal1 26312 16218 26312 16218 0 _0495_
rlabel metal1 24610 16456 24610 16456 0 _0496_
rlabel metal1 24288 16558 24288 16558 0 _0497_
rlabel metal2 28198 17340 28198 17340 0 _0498_
rlabel metal1 30498 18224 30498 18224 0 _0499_
rlabel metal2 31924 14212 31924 14212 0 _0500_
rlabel metal1 27278 16116 27278 16116 0 _0501_
rlabel via1 29946 11730 29946 11730 0 _0502_
rlabel metal1 29210 11152 29210 11152 0 _0503_
rlabel metal1 28796 11118 28796 11118 0 _0504_
rlabel metal2 29762 11424 29762 11424 0 _0505_
rlabel metal2 29026 11526 29026 11526 0 _0506_
rlabel metal1 29348 11730 29348 11730 0 _0507_
rlabel via2 27186 11747 27186 11747 0 _0508_
rlabel metal1 28888 9554 28888 9554 0 _0509_
rlabel metal1 29946 10064 29946 10064 0 _0510_
rlabel metal1 29578 9588 29578 9588 0 _0511_
rlabel metal1 29946 9690 29946 9690 0 _0512_
rlabel metal1 28980 9350 28980 9350 0 _0513_
rlabel metal1 26864 10642 26864 10642 0 _0514_
rlabel metal1 36938 13294 36938 13294 0 _0515_
rlabel metal1 31786 9996 31786 9996 0 _0516_
rlabel metal2 32154 9690 32154 9690 0 _0517_
rlabel metal1 33258 10574 33258 10574 0 _0518_
rlabel metal2 32062 9248 32062 9248 0 _0519_
rlabel metal2 32614 10880 32614 10880 0 _0520_
rlabel metal1 31832 9418 31832 9418 0 _0521_
rlabel metal1 32430 11730 32430 11730 0 _0522_
rlabel metal1 33120 10642 33120 10642 0 _0523_
rlabel metal2 34086 10574 34086 10574 0 _0524_
rlabel metal1 32982 9962 32982 9962 0 _0525_
rlabel metal1 32292 10098 32292 10098 0 _0526_
rlabel metal1 33580 10234 33580 10234 0 _0527_
rlabel metal2 33994 12002 33994 12002 0 _0528_
rlabel metal1 33580 13158 33580 13158 0 _0529_
rlabel metal2 20746 29546 20746 29546 0 _0530_
rlabel metal1 21804 29614 21804 29614 0 _0531_
rlabel metal1 23506 28560 23506 28560 0 _0532_
rlabel metal2 20654 30022 20654 30022 0 _0533_
rlabel metal2 21298 28288 21298 28288 0 _0534_
rlabel metal1 18400 29750 18400 29750 0 _0535_
rlabel metal1 14628 30566 14628 30566 0 _0536_
rlabel metal1 16928 30770 16928 30770 0 _0537_
rlabel metal1 15318 30736 15318 30736 0 _0538_
rlabel metal2 21666 29852 21666 29852 0 _0539_
rlabel metal1 22494 34544 22494 34544 0 _0540_
rlabel metal1 18124 34918 18124 34918 0 _0541_
rlabel metal2 28106 29478 28106 29478 0 _0542_
rlabel metal2 30130 30226 30130 30226 0 _0543_
rlabel metal1 28934 30226 28934 30226 0 _0544_
rlabel metal2 32154 32300 32154 32300 0 _0545_
rlabel metal1 32476 31994 32476 31994 0 _0546_
rlabel metal1 32522 30906 32522 30906 0 _0547_
rlabel metal1 31556 31926 31556 31926 0 _0548_
rlabel metal1 19780 35122 19780 35122 0 _0549_
rlabel metal1 16376 35734 16376 35734 0 _0550_
rlabel metal1 15594 35666 15594 35666 0 _0551_
rlabel metal2 16974 36006 16974 36006 0 _0552_
rlabel metal2 17710 35428 17710 35428 0 _0553_
rlabel metal2 15042 34442 15042 34442 0 _0554_
rlabel metal1 15410 34544 15410 34544 0 _0555_
rlabel metal1 16422 35054 16422 35054 0 _0556_
rlabel metal1 16836 34918 16836 34918 0 _0557_
rlabel metal2 13570 27676 13570 27676 0 _0558_
rlabel metal1 17940 27302 17940 27302 0 _0559_
rlabel metal1 15318 33830 15318 33830 0 _0560_
rlabel metal2 14214 26724 14214 26724 0 _0561_
rlabel metal1 16146 29138 16146 29138 0 _0562_
rlabel metal1 17112 27098 17112 27098 0 _0563_
rlabel metal1 15870 27098 15870 27098 0 _0564_
rlabel metal1 15686 29138 15686 29138 0 _0565_
rlabel metal1 16744 31858 16744 31858 0 _0566_
rlabel metal1 16928 30838 16928 30838 0 _0567_
rlabel metal2 15778 29920 15778 29920 0 _0568_
rlabel metal1 17526 29682 17526 29682 0 _0569_
rlabel metal1 22586 36006 22586 36006 0 _0570_
rlabel metal1 22586 34000 22586 34000 0 _0571_
rlabel metal1 22356 34578 22356 34578 0 _0572_
rlabel metal2 22310 34884 22310 34884 0 _0573_
rlabel metal1 27278 37842 27278 37842 0 _0574_
rlabel metal1 26312 37842 26312 37842 0 _0575_
rlabel metal1 25898 37298 25898 37298 0 _0576_
rlabel metal1 26588 35802 26588 35802 0 _0577_
rlabel metal1 25162 36142 25162 36142 0 _0578_
rlabel metal1 25300 38726 25300 38726 0 _0579_
rlabel metal1 23322 38862 23322 38862 0 _0580_
rlabel metal1 23598 37774 23598 37774 0 _0581_
rlabel via1 22870 38182 22870 38182 0 _0582_
rlabel metal2 25070 38726 25070 38726 0 _0583_
rlabel metal1 24242 38182 24242 38182 0 _0584_
rlabel metal2 25346 38454 25346 38454 0 _0585_
rlabel metal1 32522 39916 32522 39916 0 _0586_
rlabel metal1 32384 38930 32384 38930 0 _0587_
rlabel metal1 34730 41650 34730 41650 0 _0588_
rlabel metal1 34270 42262 34270 42262 0 _0589_
rlabel metal1 33994 40630 33994 40630 0 _0590_
rlabel metal1 33764 41038 33764 41038 0 _0591_
rlabel metal1 26266 26010 26266 26010 0 _0592_
rlabel metal1 18906 37162 18906 37162 0 _0593_
rlabel metal1 21528 34986 21528 34986 0 _0594_
rlabel metal2 20010 37842 20010 37842 0 _0595_
rlabel metal1 19688 38182 19688 38182 0 _0596_
rlabel metal2 33166 36176 33166 36176 0 _0597_
rlabel metal2 33902 40902 33902 40902 0 _0598_
rlabel metal1 34454 40970 34454 40970 0 _0599_
rlabel metal1 34454 43214 34454 43214 0 _0600_
rlabel metal1 35420 41718 35420 41718 0 _0601_
rlabel metal2 34638 42636 34638 42636 0 _0602_
rlabel metal2 32338 42228 32338 42228 0 _0603_
rlabel metal1 34316 38386 34316 38386 0 _0604_
rlabel metal1 32430 42636 32430 42636 0 _0605_
rlabel metal1 30912 43622 30912 43622 0 _0606_
rlabel metal2 31326 42636 31326 42636 0 _0607_
rlabel metal2 31970 42976 31970 42976 0 _0608_
rlabel metal2 30130 43520 30130 43520 0 _0609_
rlabel metal2 32798 42908 32798 42908 0 _0610_
rlabel metal2 33258 35802 33258 35802 0 _0611_
rlabel metal1 32890 42806 32890 42806 0 _0612_
rlabel metal1 29854 42738 29854 42738 0 _0613_
rlabel metal1 33580 38318 33580 38318 0 _0614_
rlabel metal2 30038 42874 30038 42874 0 _0615_
rlabel metal2 30590 38012 30590 38012 0 _0616_
rlabel metal1 30682 39440 30682 39440 0 _0617_
rlabel metal1 32154 39372 32154 39372 0 _0618_
rlabel metal2 32706 42432 32706 42432 0 _0619_
rlabel metal1 32660 40086 32660 40086 0 _0620_
rlabel metal2 30958 40800 30958 40800 0 _0621_
rlabel metal2 30498 40358 30498 40358 0 _0622_
rlabel metal1 30038 38216 30038 38216 0 _0623_
rlabel metal1 29946 38352 29946 38352 0 _0624_
rlabel metal1 32200 38522 32200 38522 0 _0625_
rlabel metal2 30498 39066 30498 39066 0 _0626_
rlabel metal1 34822 38318 34822 38318 0 _0627_
rlabel metal1 32660 37978 32660 37978 0 _0628_
rlabel metal1 33258 38284 33258 38284 0 _0629_
rlabel metal1 33764 36890 33764 36890 0 _0630_
rlabel metal1 33488 37230 33488 37230 0 _0631_
rlabel via1 33442 37910 33442 37910 0 _0632_
rlabel metal2 32982 37196 32982 37196 0 _0633_
rlabel metal2 33902 38012 33902 38012 0 _0634_
rlabel metal1 33396 35598 33396 35598 0 _0635_
rlabel metal1 32522 36754 32522 36754 0 _0636_
rlabel metal2 33074 36346 33074 36346 0 _0637_
rlabel metal1 32982 36074 32982 36074 0 _0638_
rlabel metal2 29486 40188 29486 40188 0 _0639_
rlabel metal2 32798 39508 32798 39508 0 _0640_
rlabel viali 32337 40040 32337 40040 0 _0641_
rlabel metal1 32522 39066 32522 39066 0 _0642_
rlabel metal2 27830 39780 27830 39780 0 _0643_
rlabel metal1 27186 39508 27186 39508 0 _0644_
rlabel metal2 26542 40018 26542 40018 0 _0645_
rlabel metal1 27048 40086 27048 40086 0 _0646_
rlabel metal1 26956 39610 26956 39610 0 _0647_
rlabel metal1 26128 42058 26128 42058 0 _0648_
rlabel metal1 27140 41242 27140 41242 0 _0649_
rlabel metal1 26450 43350 26450 43350 0 _0650_
rlabel metal1 25346 42330 25346 42330 0 _0651_
rlabel metal2 27186 41786 27186 41786 0 _0652_
rlabel metal2 24334 41276 24334 41276 0 _0653_
rlabel metal1 23690 41140 23690 41140 0 _0654_
rlabel metal1 23782 40528 23782 40528 0 _0655_
rlabel metal1 23644 40494 23644 40494 0 _0656_
rlabel metal1 24610 41106 24610 41106 0 _0657_
rlabel metal1 23368 41174 23368 41174 0 _0658_
rlabel metal1 22678 40562 22678 40562 0 _0659_
rlabel metal2 24242 41854 24242 41854 0 _0660_
rlabel metal1 22954 42568 22954 42568 0 _0661_
rlabel metal1 23092 42330 23092 42330 0 _0662_
rlabel metal1 23138 41616 23138 41616 0 _0663_
rlabel metal1 22770 41514 22770 41514 0 _0664_
rlabel metal2 17342 40834 17342 40834 0 _0665_
rlabel metal2 20562 39678 20562 39678 0 _0666_
rlabel metal2 16054 40902 16054 40902 0 _0667_
rlabel metal1 16514 41106 16514 41106 0 _0668_
rlabel metal2 16146 40698 16146 40698 0 _0669_
rlabel metal2 17710 41956 17710 41956 0 _0670_
rlabel metal2 14950 41786 14950 41786 0 _0671_
rlabel metal1 19826 41106 19826 41106 0 _0672_
rlabel metal1 19504 41650 19504 41650 0 _0673_
rlabel metal1 19520 40494 19520 40494 0 _0674_
rlabel metal1 17112 37434 17112 37434 0 _0675_
rlabel metal1 14030 36686 14030 36686 0 _0676_
rlabel metal1 19918 39066 19918 39066 0 _0677_
rlabel metal2 20102 40732 20102 40732 0 _0678_
rlabel metal1 31280 33082 31280 33082 0 _0679_
rlabel metal1 31188 34170 31188 34170 0 _0680_
rlabel metal1 30636 34170 30636 34170 0 _0681_
rlabel metal2 31878 32402 31878 32402 0 _0682_
rlabel metal1 31418 31994 31418 31994 0 _0683_
rlabel metal2 29302 29648 29302 29648 0 _0684_
rlabel metal1 16100 32334 16100 32334 0 _0685_
rlabel metal1 28474 29274 28474 29274 0 _0686_
rlabel metal2 27738 28730 27738 28730 0 _0687_
rlabel metal2 19550 35326 19550 35326 0 _0688_
rlabel metal2 19642 35462 19642 35462 0 _0689_
rlabel metal2 20010 36278 20010 36278 0 _0690_
rlabel metal1 16882 35598 16882 35598 0 _0691_
rlabel metal1 16330 36346 16330 36346 0 _0692_
rlabel metal1 14674 36890 14674 36890 0 _0693_
rlabel metal1 13110 36890 13110 36890 0 _0694_
rlabel metal2 15686 35292 15686 35292 0 _0695_
rlabel metal1 15594 35258 15594 35258 0 _0696_
rlabel metal1 14398 35802 14398 35802 0 _0697_
rlabel metal1 13248 35666 13248 35666 0 _0698_
rlabel metal1 18078 27472 18078 27472 0 _0699_
rlabel metal1 16514 28526 16514 28526 0 _0700_
rlabel metal1 17158 28050 17158 28050 0 _0701_
rlabel metal2 16238 28118 16238 28118 0 _0702_
rlabel metal1 18262 28118 18262 28118 0 _0703_
rlabel metal1 14076 26962 14076 26962 0 _0704_
rlabel metal2 14582 28356 14582 28356 0 _0705_
rlabel metal2 14582 27642 14582 27642 0 _0706_
rlabel metal1 14674 27404 14674 27404 0 _0707_
rlabel metal2 14398 27812 14398 27812 0 _0708_
rlabel metal2 12742 27404 12742 27404 0 _0709_
rlabel metal2 16974 29886 16974 29886 0 _0710_
rlabel metal1 18216 30838 18216 30838 0 _0711_
rlabel metal1 17940 30294 17940 30294 0 _0712_
rlabel metal2 18630 30396 18630 30396 0 _0713_
rlabel metal1 16560 30838 16560 30838 0 _0714_
rlabel metal1 16376 30906 16376 30906 0 _0715_
rlabel metal2 15870 31790 15870 31790 0 _0716_
rlabel metal1 14858 31450 14858 31450 0 _0717_
rlabel metal1 13248 31790 13248 31790 0 _0718_
rlabel metal2 22402 30736 22402 30736 0 _0719_
rlabel metal1 23046 29750 23046 29750 0 _0720_
rlabel metal2 22402 29580 22402 29580 0 _0721_
rlabel metal2 23230 29308 23230 29308 0 _0722_
rlabel metal1 22494 29036 22494 29036 0 _0723_
rlabel metal1 22264 28050 22264 28050 0 _0724_
rlabel metal2 22402 28492 22402 28492 0 _0725_
rlabel metal2 20930 28288 20930 28288 0 _0726_
rlabel metal2 20194 27914 20194 27914 0 _0727_
rlabel metal2 23414 34986 23414 34986 0 _0728_
rlabel metal2 22494 34442 22494 34442 0 _0729_
rlabel metal1 21758 33966 21758 33966 0 _0730_
rlabel metal1 22816 38454 22816 38454 0 _0731_
rlabel metal1 22540 38930 22540 38930 0 _0732_
rlabel metal1 22586 37910 22586 37910 0 _0733_
rlabel metal1 22816 33082 22816 33082 0 _0734_
rlabel metal1 24840 37230 24840 37230 0 _0735_
rlabel metal1 25576 37230 25576 37230 0 _0736_
rlabel metal1 25070 36210 25070 36210 0 _0737_
rlabel metal1 25576 34714 25576 34714 0 _0738_
rlabel metal1 25208 35802 25208 35802 0 _0739_
rlabel metal2 24610 35020 24610 35020 0 _0740_
rlabel metal1 26220 36822 26220 36822 0 _0741_
rlabel metal1 26499 36890 26499 36890 0 _0742_
rlabel metal1 26726 37128 26726 37128 0 _0743_
rlabel metal1 27186 37434 27186 37434 0 _0744_
rlabel metal2 25898 34527 25898 34527 0 _0745_
rlabel metal2 7498 3230 7498 3230 0 _0746_
rlabel metal2 2346 43520 2346 43520 0 _0747_
rlabel metal2 19918 3740 19918 3740 0 _0748_
rlabel metal2 2346 9316 2346 9316 0 _0749_
rlabel metal2 45126 3230 45126 3230 0 _0750_
rlabel metal1 3680 3706 3680 3706 0 _0751_
rlabel metal2 46690 20060 46690 20060 0 _0752_
rlabel metal1 10074 19754 10074 19754 0 _0753_
rlabel metal2 46414 22780 46414 22780 0 _0754_
rlabel metal2 46138 22882 46138 22882 0 _0755_
rlabel metal2 46690 17884 46690 17884 0 _0756_
rlabel metal2 22218 3876 22218 3876 0 _0757_
rlabel metal2 17434 43044 17434 43044 0 _0758_
rlabel metal2 5106 42466 5106 42466 0 _0759_
rlabel metal2 20562 43996 20562 43996 0 _0760_
rlabel metal2 4094 14756 4094 14756 0 _0761_
rlabel metal2 47150 16728 47150 16728 0 _0762_
rlabel metal1 47288 36074 47288 36074 0 _0763_
rlabel metal1 5520 46002 5520 46002 0 _0764_
rlabel metal2 47150 24990 47150 24990 0 _0765_
rlabel metal2 2898 10846 2898 10846 0 _0766_
rlabel metal1 47288 42602 47288 42602 0 _0767_
rlabel metal1 29900 45594 29900 45594 0 _0768_
rlabel metal2 12558 10846 12558 10846 0 _0769_
rlabel metal1 46920 18802 46920 18802 0 _0770_
rlabel metal2 1794 5100 1794 5100 0 _0771_
rlabel metal2 47610 5202 47610 5202 0 _0772_
rlabel metal1 1794 45832 1794 45832 0 _0773_
rlabel metal2 45402 4828 45402 4828 0 _0774_
rlabel metal1 5520 3434 5520 3434 0 _0775_
rlabel metal1 46920 12274 46920 12274 0 _0776_
rlabel metal1 45770 46138 45770 46138 0 _0777_
rlabel metal2 46690 46172 46690 46172 0 _0778_
rlabel metal2 33166 46308 33166 46308 0 _0779_
rlabel via1 6854 2363 6854 2363 0 _0780_
rlabel metal2 2438 43554 2438 43554 0 _0781_
rlabel metal1 47288 29682 47288 29682 0 _0782_
rlabel metal2 22770 46308 22770 46308 0 _0783_
rlabel metal1 46322 46478 46322 46478 0 _0784_
rlabel metal2 4922 20196 4922 20196 0 _0785_
rlabel metal2 18538 2788 18538 2788 0 _0786_
rlabel metal2 2898 15232 2898 15232 0 _0787_
rlabel metal1 47288 27370 47288 27370 0 _0788_
rlabel metal2 2070 3502 2070 3502 0 _0789_
rlabel metal2 2254 7582 2254 7582 0 _0790_
rlabel metal2 40158 3502 40158 3502 0 _0791_
rlabel metal2 47150 40222 47150 40222 0 _0792_
rlabel metal2 2346 40868 2346 40868 0 _0793_
rlabel metal1 47288 26282 47288 26282 0 _0794_
rlabel metal2 45954 40868 45954 40868 0 _0795_
rlabel metal2 46138 3740 46138 3740 0 _0796_
rlabel metal2 10534 22882 10534 22882 0 _0797_
rlabel metal1 40158 45594 40158 45594 0 _0798_
rlabel metal2 10258 21148 10258 21148 0 _0799_
rlabel metal2 32522 3230 32522 3230 0 _0800_
rlabel metal2 40894 21794 40894 21794 0 _0801_
rlabel metal2 27370 3230 27370 3230 0 _0802_
rlabel metal1 37030 45526 37030 45526 0 _0803_
rlabel metal2 10074 5100 10074 5100 0 _0804_
rlabel metal1 39238 46138 39238 46138 0 _0805_
rlabel metal1 16606 3434 16606 3434 0 _0806_
rlabel metal1 46736 5270 46736 5270 0 _0807_
rlabel metal1 2346 6426 2346 6426 0 _0808_
rlabel metal1 2346 14042 2346 14042 0 _0809_
rlabel metal1 4002 45526 4002 45526 0 _0810_
rlabel metal2 47886 6562 47886 6562 0 _0811_
rlabel metal1 47288 41650 47288 41650 0 _0812_
rlabel metal1 47288 37162 47288 37162 0 _0813_
rlabel metal1 15272 45594 15272 45594 0 _0814_
rlabel metal2 47886 44642 47886 44642 0 _0815_
rlabel metal1 25806 3434 25806 3434 0 _0816_
rlabel metal2 39238 5678 39238 5678 0 _0817_
rlabel metal1 42136 45526 42136 45526 0 _0818_
rlabel metal2 24978 3230 24978 3230 0 _0819_
rlabel metal2 43286 4318 43286 4318 0 _0820_
rlabel metal2 2346 32606 2346 32606 0 _0821_
rlabel metal1 46736 16490 46736 16490 0 _0822_
rlabel metal2 12558 46308 12558 46308 0 _0823_
rlabel via1 4186 2499 4186 2499 0 _0824_
rlabel metal2 10718 3740 10718 3740 0 _0825_
rlabel metal2 2622 16354 2622 16354 0 _0826_
rlabel metal1 47288 28458 47288 28458 0 _0827_
rlabel metal2 47150 15266 47150 15266 0 _0828_
rlabel metal1 46920 13362 46920 13362 0 _0829_
rlabel metal2 2898 4624 2898 4624 0 _0830_
rlabel metal1 13754 46138 13754 46138 0 _0831_
rlabel metal1 46046 2482 46046 2482 0 _0832_
rlabel metal2 13202 3230 13202 3230 0 _0833_
rlabel metal1 35604 45594 35604 45594 0 _0834_
rlabel metal2 14490 46308 14490 46308 0 _0835_
rlabel metal2 46690 21148 46690 21148 0 _0836_
rlabel metal2 2070 46308 2070 46308 0 _0837_
rlabel metal2 4370 3230 4370 3230 0 _0838_
rlabel metal2 24886 45730 24886 45730 0 _0839_
rlabel metal1 25254 45594 25254 45594 0 _0840_
rlabel metal1 46276 4046 46276 4046 0 _0841_
rlabel metal2 47886 39202 47886 39202 0 _0842_
rlabel metal1 29164 46138 29164 46138 0 _0843_
rlabel metal1 42320 2618 42320 2618 0 _0844_
rlabel metal2 47886 32674 47886 32674 0 _0845_
rlabel metal1 6302 45526 6302 45526 0 _0846_
rlabel metal2 41446 3740 41446 3740 0 _0847_
rlabel metal2 1794 25500 1794 25500 0 _0848_
rlabel metal1 19688 2618 19688 2618 0 _0849_
rlabel metal1 10672 44506 10672 44506 0 _0850_
rlabel metal2 2346 21284 2346 21284 0 _0851_
rlabel metal2 2346 11492 2346 11492 0 _0852_
rlabel metal1 2300 17850 2300 17850 0 _0853_
rlabel metal1 2346 42602 2346 42602 0 active
rlabel metal1 32476 14382 32476 14382 0 clknet_0_wb_clk_i
rlabel metal1 17802 21998 17802 21998 0 clknet_4_0_0_wb_clk_i
rlabel metal1 39422 13940 39422 13940 0 clknet_4_10_0_wb_clk_i
rlabel metal1 43746 22474 43746 22474 0 clknet_4_11_0_wb_clk_i
rlabel metal1 33718 21556 33718 21556 0 clknet_4_12_0_wb_clk_i
rlabel metal1 27186 21556 27186 21556 0 clknet_4_13_0_wb_clk_i
rlabel metal1 36754 21998 36754 21998 0 clknet_4_14_0_wb_clk_i
rlabel metal2 36662 32946 36662 32946 0 clknet_4_15_0_wb_clk_i
rlabel metal2 13846 25024 13846 25024 0 clknet_4_1_0_wb_clk_i
rlabel metal1 19642 16626 19642 16626 0 clknet_4_2_0_wb_clk_i
rlabel metal1 20102 21556 20102 21556 0 clknet_4_3_0_wb_clk_i
rlabel metal1 12098 36142 12098 36142 0 clknet_4_4_0_wb_clk_i
rlabel metal1 14214 39474 14214 39474 0 clknet_4_5_0_wb_clk_i
rlabel metal2 30314 35360 30314 35360 0 clknet_4_6_0_wb_clk_i
rlabel metal1 27140 34578 27140 34578 0 clknet_4_7_0_wb_clk_i
rlabel metal1 32798 12886 32798 12886 0 clknet_4_8_0_wb_clk_i
rlabel metal1 34362 14892 34362 14892 0 clknet_4_9_0_wb_clk_i
rlabel metal1 20102 40154 20102 40154 0 gps_channel0.ca_full_chip
rlabel metal1 9200 28050 9200 28050 0 gps_channel0.ca_gen.g1\[10\]
rlabel metal2 8326 29206 8326 29206 0 gps_channel0.ca_gen.g1\[1\]
rlabel metal1 9706 30022 9706 30022 0 gps_channel0.ca_gen.g1\[2\]
rlabel metal1 7682 30226 7682 30226 0 gps_channel0.ca_gen.g1\[3\]
rlabel metal2 5382 31008 5382 31008 0 gps_channel0.ca_gen.g1\[4\]
rlabel metal1 5474 28968 5474 28968 0 gps_channel0.ca_gen.g1\[5\]
rlabel metal1 4922 27642 4922 27642 0 gps_channel0.ca_gen.g1\[6\]
rlabel metal2 5750 27370 5750 27370 0 gps_channel0.ca_gen.g1\[7\]
rlabel metal2 6946 26078 6946 26078 0 gps_channel0.ca_gen.g1\[8\]
rlabel metal2 8418 27098 8418 27098 0 gps_channel0.ca_gen.g1\[9\]
rlabel metal1 12834 19482 12834 19482 0 gps_channel0.ca_gen.g2\[10\]
rlabel metal2 16054 21284 16054 21284 0 gps_channel0.ca_gen.g2\[1\]
rlabel metal2 13294 21862 13294 21862 0 gps_channel0.ca_gen.g2\[2\]
rlabel metal2 13202 21794 13202 21794 0 gps_channel0.ca_gen.g2\[3\]
rlabel metal1 15686 22066 15686 22066 0 gps_channel0.ca_gen.g2\[4\]
rlabel metal2 16054 18394 16054 18394 0 gps_channel0.ca_gen.g2\[5\]
rlabel metal1 14996 16966 14996 16966 0 gps_channel0.ca_gen.g2\[6\]
rlabel metal2 15226 15606 15226 15606 0 gps_channel0.ca_gen.g2\[7\]
rlabel metal2 13202 16898 13202 16898 0 gps_channel0.ca_gen.g2\[8\]
rlabel metal2 12742 18020 12742 18020 0 gps_channel0.ca_gen.g2\[9\]
rlabel metal1 19458 17306 19458 17306 0 gps_channel0.ca_gen.g2_init\[10\]
rlabel metal1 19228 20026 19228 20026 0 gps_channel0.ca_gen.g2_init\[1\]
rlabel metal1 20700 21658 20700 21658 0 gps_channel0.ca_gen.g2_init\[2\]
rlabel metal1 20562 20298 20562 20298 0 gps_channel0.ca_gen.g2_init\[3\]
rlabel metal2 18814 21658 18814 21658 0 gps_channel0.ca_gen.g2_init\[4\]
rlabel metal1 16514 21998 16514 21998 0 gps_channel0.ca_gen.g2_init\[5\]
rlabel metal1 18124 18598 18124 18598 0 gps_channel0.ca_gen.g2_init\[6\]
rlabel metal1 19136 15470 19136 15470 0 gps_channel0.ca_gen.g2_init\[7\]
rlabel metal1 17250 15470 17250 15470 0 gps_channel0.ca_gen.g2_init\[8\]
rlabel metal2 17526 16320 17526 16320 0 gps_channel0.ca_gen.g2_init\[9\]
rlabel metal2 31418 33932 31418 33932 0 gps_channel0.ca_nco.accumulator\[0\]
rlabel metal1 24656 29546 24656 29546 0 gps_channel0.ca_nco.accumulator\[10\]
rlabel metal2 20838 28288 20838 28288 0 gps_channel0.ca_nco.accumulator\[11\]
rlabel metal1 21390 34952 21390 34952 0 gps_channel0.ca_nco.accumulator\[12\]
rlabel metal2 22494 38012 22494 38012 0 gps_channel0.ca_nco.accumulator\[13\]
rlabel metal1 26128 35734 26128 35734 0 gps_channel0.ca_nco.accumulator\[14\]
rlabel metal1 28106 38284 28106 38284 0 gps_channel0.ca_nco.accumulator\[15\]
rlabel metal1 34546 40970 34546 40970 0 gps_channel0.ca_nco.accumulator\[16\]
rlabel metal1 33626 42806 33626 42806 0 gps_channel0.ca_nco.accumulator\[17\]
rlabel metal1 30728 43350 30728 43350 0 gps_channel0.ca_nco.accumulator\[18\]
rlabel metal1 30360 42738 30360 42738 0 gps_channel0.ca_nco.accumulator\[19\]
rlabel metal1 33212 32198 33212 32198 0 gps_channel0.ca_nco.accumulator\[1\]
rlabel metal1 34086 38386 34086 38386 0 gps_channel0.ca_nco.accumulator\[20\]
rlabel metal1 35190 38352 35190 38352 0 gps_channel0.ca_nco.accumulator\[21\]
rlabel metal1 32890 37128 32890 37128 0 gps_channel0.ca_nco.accumulator\[22\]
rlabel metal1 32522 36346 32522 36346 0 gps_channel0.ca_nco.accumulator\[23\]
rlabel metal1 26772 41174 26772 41174 0 gps_channel0.ca_nco.accumulator\[24\]
rlabel metal2 26174 41888 26174 41888 0 gps_channel0.ca_nco.accumulator\[25\]
rlabel metal1 21942 40698 21942 40698 0 gps_channel0.ca_nco.accumulator\[26\]
rlabel metal1 22218 42772 22218 42772 0 gps_channel0.ca_nco.accumulator\[27\]
rlabel metal1 17020 40426 17020 40426 0 gps_channel0.ca_nco.accumulator\[28\]
rlabel metal1 4922 42602 4922 42602 0 gps_channel0.ca_nco.accumulator\[29\]
rlabel metal1 28750 29512 28750 29512 0 gps_channel0.ca_nco.accumulator\[2\]
rlabel metal1 19688 41174 19688 41174 0 gps_channel0.ca_nco.accumulator\[30\]
rlabel metal1 18538 35020 18538 35020 0 gps_channel0.ca_nco.accumulator\[3\]
rlabel metal2 13662 36992 13662 36992 0 gps_channel0.ca_nco.accumulator\[4\]
rlabel metal2 13846 35904 13846 35904 0 gps_channel0.ca_nco.accumulator\[5\]
rlabel via1 18428 28050 18428 28050 0 gps_channel0.ca_nco.accumulator\[6\]
rlabel metal2 13478 26826 13478 26826 0 gps_channel0.ca_nco.accumulator\[7\]
rlabel via1 18796 30226 18796 30226 0 gps_channel0.ca_nco.accumulator\[8\]
rlabel metal2 13570 30906 13570 30906 0 gps_channel0.ca_nco.accumulator\[9\]
rlabel metal1 29992 35462 29992 35462 0 gps_channel0.ca_nco.phase_in\[0\]
rlabel metal1 25530 27302 25530 27302 0 gps_channel0.ca_nco.phase_in\[10\]
rlabel metal1 23046 26554 23046 26554 0 gps_channel0.ca_nco.phase_in\[11\]
rlabel metal2 22310 32980 22310 32980 0 gps_channel0.ca_nco.phase_in\[12\]
rlabel metal2 23414 32640 23414 32640 0 gps_channel0.ca_nco.phase_in\[13\]
rlabel metal2 25990 33252 25990 33252 0 gps_channel0.ca_nco.phase_in\[14\]
rlabel metal1 26174 33082 26174 33082 0 gps_channel0.ca_nco.phase_in\[15\]
rlabel metal2 30406 31994 30406 31994 0 gps_channel0.ca_nco.phase_in\[1\]
rlabel metal2 29210 27744 29210 27744 0 gps_channel0.ca_nco.phase_in\[2\]
rlabel metal2 18446 37536 18446 37536 0 gps_channel0.ca_nco.phase_in\[3\]
rlabel metal2 16146 37604 16146 37604 0 gps_channel0.ca_nco.phase_in\[4\]
rlabel metal1 15134 38318 15134 38318 0 gps_channel0.ca_nco.phase_in\[5\]
rlabel metal1 21482 25262 21482 25262 0 gps_channel0.ca_nco.phase_in\[6\]
rlabel metal1 15272 24650 15272 24650 0 gps_channel0.ca_nco.phase_in\[7\]
rlabel metal1 19458 24922 19458 24922 0 gps_channel0.ca_nco.phase_in\[8\]
rlabel metal1 17112 32878 17112 32878 0 gps_channel0.ca_nco.phase_in\[9\]
rlabel metal2 25898 26452 25898 26452 0 gps_channel0.ca_nco.phase_sync
rlabel metal1 31326 33422 31326 33422 0 gps_channel0.ca_nco.step\[0\]
rlabel metal1 24426 29614 24426 29614 0 gps_channel0.ca_nco.step\[10\]
rlabel metal1 21298 27438 21298 27438 0 gps_channel0.ca_nco.step\[11\]
rlabel metal2 20930 34544 20930 34544 0 gps_channel0.ca_nco.step\[12\]
rlabel metal2 21758 37434 21758 37434 0 gps_channel0.ca_nco.step\[13\]
rlabel metal2 27462 31994 27462 31994 0 gps_channel0.ca_nco.step\[14\]
rlabel metal1 27922 37298 27922 37298 0 gps_channel0.ca_nco.step\[15\]
rlabel metal1 32338 39304 32338 39304 0 gps_channel0.ca_nco.step\[16\]
rlabel metal2 32154 31008 32154 31008 0 gps_channel0.ca_nco.step\[1\]
rlabel metal2 28566 29070 28566 29070 0 gps_channel0.ca_nco.step\[2\]
rlabel metal2 18906 32572 18906 32572 0 gps_channel0.ca_nco.step\[3\]
rlabel metal2 13754 35360 13754 35360 0 gps_channel0.ca_nco.step\[4\]
rlabel metal1 15410 33524 15410 33524 0 gps_channel0.ca_nco.step\[5\]
rlabel metal2 17250 26758 17250 26758 0 gps_channel0.ca_nco.step\[6\]
rlabel metal2 13662 27438 13662 27438 0 gps_channel0.ca_nco.step\[7\]
rlabel metal2 17066 30804 17066 30804 0 gps_channel0.ca_nco.step\[8\]
rlabel metal1 13248 30022 13248 30022 0 gps_channel0.ca_nco.step\[9\]
rlabel metal1 22034 4012 22034 4012 0 gps_channel0.lo_i
rlabel metal1 40848 23698 40848 23698 0 gps_channel0.lo_nco.accumulator\[0\]
rlabel via1 28732 14382 28732 14382 0 gps_channel0.lo_nco.accumulator\[10\]
rlabel metal1 24932 16082 24932 16082 0 gps_channel0.lo_nco.accumulator\[11\]
rlabel metal2 27554 11594 27554 11594 0 gps_channel0.lo_nco.accumulator\[12\]
rlabel metal1 27646 10234 27646 10234 0 gps_channel0.lo_nco.accumulator\[13\]
rlabel metal1 31464 10710 31464 10710 0 gps_channel0.lo_nco.accumulator\[14\]
rlabel metal1 34914 12614 34914 12614 0 gps_channel0.lo_nco.accumulator\[15\]
rlabel metal2 38042 13668 38042 13668 0 gps_channel0.lo_nco.accumulator\[16\]
rlabel metal1 38778 10438 38778 10438 0 gps_channel0.lo_nco.accumulator\[17\]
rlabel metal1 39054 9350 39054 9350 0 gps_channel0.lo_nco.accumulator\[18\]
rlabel metal1 39192 10642 39192 10642 0 gps_channel0.lo_nco.accumulator\[19\]
rlabel metal1 38502 21964 38502 21964 0 gps_channel0.lo_nco.accumulator\[1\]
rlabel metal2 45494 13668 45494 13668 0 gps_channel0.lo_nco.accumulator\[20\]
rlabel metal1 43930 14994 43930 14994 0 gps_channel0.lo_nco.accumulator\[21\]
rlabel metal2 44942 10812 44942 10812 0 gps_channel0.lo_nco.accumulator\[22\]
rlabel metal2 43930 10642 43930 10642 0 gps_channel0.lo_nco.accumulator\[23\]
rlabel metal2 40802 14178 40802 14178 0 gps_channel0.lo_nco.accumulator\[24\]
rlabel metal1 41285 15946 41285 15946 0 gps_channel0.lo_nco.accumulator\[25\]
rlabel metal1 43746 18326 43746 18326 0 gps_channel0.lo_nco.accumulator\[26\]
rlabel metal2 43470 17510 43470 17510 0 gps_channel0.lo_nco.accumulator\[27\]
rlabel metal1 45310 22406 45310 22406 0 gps_channel0.lo_nco.accumulator\[28\]
rlabel metal1 45862 21658 45862 21658 0 gps_channel0.lo_nco.accumulator\[29\]
rlabel metal1 37168 21862 37168 21862 0 gps_channel0.lo_nco.accumulator\[2\]
rlabel metal1 21390 18360 21390 18360 0 gps_channel0.lo_nco.accumulator\[30\]
rlabel metal2 34638 26316 34638 26316 0 gps_channel0.lo_nco.accumulator\[3\]
rlabel metal1 31924 21862 31924 21862 0 gps_channel0.lo_nco.accumulator\[4\]
rlabel metal2 37490 19550 37490 19550 0 gps_channel0.lo_nco.accumulator\[5\]
rlabel metal1 36662 17034 36662 17034 0 gps_channel0.lo_nco.accumulator\[6\]
rlabel metal1 34914 16456 34914 16456 0 gps_channel0.lo_nco.accumulator\[7\]
rlabel metal1 28980 20434 28980 20434 0 gps_channel0.lo_nco.accumulator\[8\]
rlabel metal1 26910 19210 26910 19210 0 gps_channel0.lo_nco.accumulator\[9\]
rlabel metal1 36754 24310 36754 24310 0 gps_channel0.lo_nco.phase_in\[0\]
rlabel metal1 28750 14042 28750 14042 0 gps_channel0.lo_nco.phase_in\[10\]
rlabel metal1 22995 16082 22995 16082 0 gps_channel0.lo_nco.phase_in\[11\]
rlabel metal2 22126 11968 22126 11968 0 gps_channel0.lo_nco.phase_in\[12\]
rlabel metal1 23230 13906 23230 13906 0 gps_channel0.lo_nco.phase_in\[13\]
rlabel metal1 31372 14042 31372 14042 0 gps_channel0.lo_nco.phase_in\[14\]
rlabel metal2 33810 13498 33810 13498 0 gps_channel0.lo_nco.phase_in\[15\]
rlabel metal1 34730 21998 34730 21998 0 gps_channel0.lo_nco.phase_in\[1\]
rlabel metal1 35282 23494 35282 23494 0 gps_channel0.lo_nco.phase_in\[2\]
rlabel metal2 32522 25704 32522 25704 0 gps_channel0.lo_nco.phase_in\[3\]
rlabel metal1 31004 22406 31004 22406 0 gps_channel0.lo_nco.phase_in\[4\]
rlabel metal1 32384 19686 32384 19686 0 gps_channel0.lo_nco.phase_in\[5\]
rlabel metal1 32384 18122 32384 18122 0 gps_channel0.lo_nco.phase_in\[6\]
rlabel metal1 33718 15980 33718 15980 0 gps_channel0.lo_nco.phase_in\[7\]
rlabel metal1 28474 21522 28474 21522 0 gps_channel0.lo_nco.phase_in\[8\]
rlabel metal1 24932 18938 24932 18938 0 gps_channel0.lo_nco.phase_in\[9\]
rlabel metal2 25898 21726 25898 21726 0 gps_channel0.lo_nco.phase_sync
rlabel metal2 40710 26180 40710 26180 0 gps_channel0.lo_nco.step\[0\]
rlabel metal1 26910 14382 26910 14382 0 gps_channel0.lo_nco.step\[10\]
rlabel metal1 23874 15334 23874 15334 0 gps_channel0.lo_nco.step\[11\]
rlabel metal2 23322 10778 23322 10778 0 gps_channel0.lo_nco.step\[12\]
rlabel metal2 23230 9724 23230 9724 0 gps_channel0.lo_nco.step\[13\]
rlabel metal1 25346 10744 25346 10744 0 gps_channel0.lo_nco.step\[14\]
rlabel metal1 33350 11084 33350 11084 0 gps_channel0.lo_nco.step\[15\]
rlabel metal1 38088 14382 38088 14382 0 gps_channel0.lo_nco.step\[16\]
rlabel metal1 38962 21998 38962 21998 0 gps_channel0.lo_nco.step\[1\]
rlabel metal1 36064 25942 36064 25942 0 gps_channel0.lo_nco.step\[2\]
rlabel metal1 32384 27302 32384 27302 0 gps_channel0.lo_nco.step\[3\]
rlabel metal1 31786 22644 31786 22644 0 gps_channel0.lo_nco.step\[4\]
rlabel metal2 38226 20060 38226 20060 0 gps_channel0.lo_nco.step\[5\]
rlabel metal1 39330 17850 39330 17850 0 gps_channel0.lo_nco.step\[6\]
rlabel metal1 33442 16422 33442 16422 0 gps_channel0.lo_nco.step\[7\]
rlabel metal1 28474 20502 28474 20502 0 gps_channel0.lo_nco.step\[8\]
rlabel metal1 27002 18258 27002 18258 0 gps_channel0.lo_nco.step\[9\]
rlabel metal2 10074 20094 10074 20094 0 gps_channel0.prompt_i
rlabel metal1 10304 19278 10304 19278 0 gps_channel0.prompt_q
rlabel metal1 9108 47090 9108 47090 0 io_in[23]
rlabel metal2 26450 2166 26450 2166 0 io_oeb[0]
rlabel metal2 2806 16847 2806 16847 0 io_oeb[10]
rlabel metal3 48814 28628 48814 28628 0 io_oeb[11]
rlabel metal3 48814 15028 48814 15028 0 io_oeb[12]
rlabel metal3 48814 13668 48814 13668 0 io_oeb[13]
rlabel metal3 1832 4828 1832 4828 0 io_oeb[14]
rlabel metal1 14490 47090 14490 47090 0 io_oeb[15]
rlabel metal3 48124 2108 48124 2108 0 io_oeb[16]
rlabel metal2 13570 1860 13570 1860 0 io_oeb[17]
rlabel metal2 36110 47644 36110 47644 0 io_oeb[18]
rlabel metal2 14858 47882 14858 47882 0 io_oeb[19]
rlabel metal1 39698 3638 39698 3638 0 io_oeb[1]
rlabel metal3 48814 21828 48814 21828 0 io_oeb[20]
rlabel metal2 2346 47889 2346 47889 0 io_oeb[21]
rlabel metal2 5198 1860 5198 1860 0 io_oeb[22]
rlabel metal1 25852 45866 25852 45866 0 io_oeb[23]
rlabel metal2 25806 47882 25806 47882 0 io_oeb[24]
rlabel metal1 47472 4046 47472 4046 0 io_oeb[25]
rlabel metal3 48814 39508 48814 39508 0 io_oeb[26]
rlabel metal2 29670 47882 29670 47882 0 io_oeb[27]
rlabel metal1 42504 2890 42504 2890 0 io_oeb[28]
rlabel metal3 48860 32708 48860 32708 0 io_oeb[29]
rlabel metal1 43102 46444 43102 46444 0 io_oeb[2]
rlabel metal1 4324 46614 4324 46614 0 io_oeb[30]
rlabel metal2 41262 2200 41262 2200 0 io_oeb[31]
rlabel metal2 2806 25279 2806 25279 0 io_oeb[32]
rlabel metal1 21482 2924 21482 2924 0 io_oeb[33]
rlabel metal2 11086 45227 11086 45227 0 io_oeb[34]
rlabel metal2 2806 21641 2806 21641 0 io_oeb[35]
rlabel metal3 1740 11628 1740 11628 0 io_oeb[36]
rlabel metal2 2806 18309 2806 18309 0 io_oeb[37]
rlabel metal2 25806 1860 25806 1860 0 io_oeb[3]
rlabel metal3 48860 68 48860 68 0 io_oeb[4]
rlabel metal2 2806 32521 2806 32521 0 io_oeb[5]
rlabel metal3 48814 17748 48814 17748 0 io_oeb[6]
rlabel metal2 12926 47882 12926 47882 0 io_oeb[7]
rlabel metal2 4554 1622 4554 1622 0 io_oeb[8]
rlabel metal2 10994 2166 10994 2166 0 io_oeb[9]
rlabel metal3 48814 46988 48814 46988 0 io_out[0]
rlabel metal3 48814 27948 48814 27948 0 io_out[10]
rlabel metal3 1740 2788 1740 2788 0 io_out[11]
rlabel metal2 2806 7429 2806 7429 0 io_out[12]
rlabel metal2 40618 1860 40618 1860 0 io_out[13]
rlabel metal3 48860 40188 48860 40188 0 io_out[14]
rlabel metal2 2806 41293 2806 41293 0 io_out[15]
rlabel metal3 48814 26588 48814 26588 0 io_out[16]
rlabel metal1 46690 46886 46690 46886 0 io_out[17]
rlabel metal2 47058 2166 47058 2166 0 io_out[18]
rlabel metal2 11086 23324 11086 23324 0 io_out[19]
rlabel metal2 33534 47882 33534 47882 0 io_out[1]
rlabel metal2 40618 47644 40618 47644 0 io_out[20]
rlabel metal3 2108 40868 2108 40868 0 io_out[21]
rlabel metal1 32522 2958 32522 2958 0 io_out[22]
rlabel metal2 46598 22321 46598 22321 0 io_out[23]
rlabel metal2 27738 1860 27738 1860 0 io_out[24]
rlabel metal1 37950 46444 37950 46444 0 io_out[25]
rlabel metal3 2108 5508 2108 5508 0 io_out[26]
rlabel metal2 38686 47848 38686 47848 0 io_out[27]
rlabel metal2 17434 2166 17434 2166 0 io_out[28]
rlabel metal3 48308 1428 48308 1428 0 io_out[29]
rlabel metal2 7130 1622 7130 1622 0 io_out[2]
rlabel via2 2806 6851 2806 6851 0 io_out[30]
rlabel metal3 1740 14348 1740 14348 0 io_out[31]
rlabel metal3 1832 47668 1832 47668 0 io_out[32]
rlabel metal3 48814 6868 48814 6868 0 io_out[33]
rlabel metal3 48814 41548 48814 41548 0 io_out[34]
rlabel metal3 48814 38148 48814 38148 0 io_out[35]
rlabel metal2 15502 47644 15502 47644 0 io_out[36]
rlabel metal3 48814 44948 48814 44948 0 io_out[37]
rlabel metal3 1740 43588 1740 43588 0 io_out[3]
rlabel metal3 48860 29308 48860 29308 0 io_out[4]
rlabel metal2 23230 47882 23230 47882 0 io_out[5]
rlabel metal2 48346 47950 48346 47950 0 io_out[6]
rlabel metal3 1832 20468 1832 20468 0 io_out[7]
rlabel metal2 19366 1860 19366 1860 0 io_out[8]
rlabel metal3 1740 15028 1740 15028 0 io_out[9]
rlabel metal2 47886 8347 47886 8347 0 la1_data_in[0]
rlabel metal2 31786 47073 31786 47073 0 la1_data_in[16]
rlabel metal1 24288 47022 24288 47022 0 la1_data_in[17]
rlabel metal2 43838 1554 43838 1554 0 la1_data_in[18]
rlabel metal1 17480 47022 17480 47022 0 la1_data_in[19]
rlabel metal2 20010 1588 20010 1588 0 la1_data_in[1]
rlabel metal3 1142 36788 1142 36788 0 la1_data_in[20]
rlabel metal1 48484 47022 48484 47022 0 la1_data_in[21]
rlabel via2 47978 8891 47978 8891 0 la1_data_in[22]
rlabel metal3 1740 748 1740 748 0 la1_data_in[23]
rlabel metal2 14214 1588 14214 1588 0 la1_data_in[24]
rlabel metal3 1142 38828 1142 38828 0 la1_data_in[25]
rlabel metal2 48070 3247 48070 3247 0 la1_data_in[26]
rlabel metal2 29026 1554 29026 1554 0 la1_data_in[27]
rlabel metal3 1142 34068 1142 34068 0 la1_data_in[28]
rlabel metal1 828 44846 828 44846 0 la1_data_in[29]
rlabel metal2 11638 1588 11638 1588 0 la1_data_in[2]
rlabel metal2 1334 1554 1334 1554 0 la1_data_in[30]
rlabel metal2 38686 1588 38686 1588 0 la1_data_in[31]
rlabel metal3 1142 32028 1142 32028 0 la1_data_in[3]
rlabel metal1 42596 47022 42596 47022 0 la1_data_in[4]
rlabel metal1 48208 24786 48208 24786 0 la1_data_in[5]
rlabel metal1 19458 47022 19458 47022 0 la1_data_in[6]
rlabel metal2 7774 1860 7774 1860 0 la1_data_out[0]
rlabel metal3 48722 12308 48722 12308 0 la1_data_out[10]
rlabel metal2 22586 2404 22586 2404 0 la1_data_out[11]
rlabel metal2 46598 46053 46598 46053 0 la1_data_out[12]
rlabel metal1 5244 45866 5244 45866 0 la1_data_out[13]
rlabel metal1 24656 43826 24656 43826 0 la1_data_out[14]
rlabel metal3 1786 1428 1786 1428 0 la1_data_out[15]
rlabel metal3 48124 17068 48124 17068 0 la1_data_out[16]
rlabel metal3 48814 36108 48814 36108 0 la1_data_out[17]
rlabel metal2 5842 47644 5842 47644 0 la1_data_out[18]
rlabel metal3 48814 25908 48814 25908 0 la1_data_out[19]
rlabel metal3 1740 45628 1740 45628 0 la1_data_out[1]
rlabel metal3 1924 10268 1924 10268 0 la1_data_out[20]
rlabel metal3 48814 42908 48814 42908 0 la1_data_out[21]
rlabel metal1 30958 45866 30958 45866 0 la1_data_out[22]
rlabel metal2 12926 2234 12926 2234 0 la1_data_out[23]
rlabel metal3 48814 19108 48814 19108 0 la1_data_out[24]
rlabel metal3 1740 3468 1740 3468 0 la1_data_out[25]
rlabel metal3 48814 5508 48814 5508 0 la1_data_out[26]
rlabel metal2 2806 47175 2806 47175 0 la1_data_out[27]
rlabel metal1 45402 2890 45402 2890 0 la1_data_out[28]
rlabel metal2 6486 2166 6486 2166 0 la1_data_out[29]
rlabel metal2 20654 2166 20654 2166 0 la1_data_out[2]
rlabel metal3 48814 12988 48814 12988 0 la1_data_out[30]
rlabel metal3 48308 49028 48308 49028 0 la1_data_out[31]
rlabel metal3 1740 9588 1740 9588 0 la1_data_out[3]
rlabel metal2 45770 1860 45770 1860 0 la1_data_out[4]
rlabel metal2 3266 2370 3266 2370 0 la1_data_out[5]
rlabel metal3 48814 20468 48814 20468 0 la1_data_out[6]
rlabel metal2 230 18157 230 18157 0 la1_data_out[7]
rlabel metal3 48032 37468 48032 37468 0 la1_data_out[8]
rlabel metal2 47341 49300 47341 49300 0 la1_data_out[9]
rlabel metal1 1886 42534 1886 42534 0 net1
rlabel metal1 17250 19176 17250 19176 0 net10
rlabel metal2 47978 15266 47978 15266 0 net100
rlabel metal1 46506 13396 46506 13396 0 net101
rlabel metal1 2024 5134 2024 5134 0 net102
rlabel metal1 14030 47022 14030 47022 0 net103
rlabel metal1 45034 2482 45034 2482 0 net104
rlabel metal2 13018 3468 13018 3468 0 net105
rlabel metal2 35466 46172 35466 46172 0 net106
rlabel metal1 14398 45458 14398 45458 0 net107
rlabel metal1 46506 21012 46506 21012 0 net108
rlabel metal1 1886 46444 1886 46444 0 net109
rlabel metal1 39146 18190 39146 18190 0 net11
rlabel metal1 4600 2958 4600 2958 0 net110
rlabel metal1 24380 45934 24380 45934 0 net111
rlabel metal1 24794 46580 24794 46580 0 net112
rlabel metal1 46690 3978 46690 3978 0 net113
rlabel metal2 46506 39644 46506 39644 0 net114
rlabel metal1 28796 46478 28796 46478 0 net115
rlabel metal2 42642 3264 42642 3264 0 net116
rlabel metal1 47242 32946 47242 32946 0 net117
rlabel metal2 4186 46818 4186 46818 0 net118
rlabel metal2 40802 3740 40802 3740 0 net119
rlabel metal2 2898 2142 2898 2142 0 net12
rlabel metal1 1932 24786 1932 24786 0 net120
rlabel metal1 19642 3060 19642 3060 0 net121
rlabel metal2 10534 45084 10534 45084 0 net122
rlabel metal2 2070 21760 2070 21760 0 net123
rlabel metal2 2070 11968 2070 11968 0 net124
rlabel metal2 2070 18496 2070 18496 0 net125
rlabel metal1 16054 2618 16054 2618 0 net13
rlabel metal1 1840 38726 1840 38726 0 net14
rlabel metal1 27692 14382 27692 14382 0 net15
rlabel metal1 26910 2278 26910 2278 0 net16
rlabel metal2 1794 34272 1794 34272 0 net17
rlabel metal2 1794 40800 1794 40800 0 net18
rlabel metal2 17756 16560 17756 16560 0 net19
rlabel metal1 9154 47022 9154 47022 0 net2
rlabel metal1 20286 2516 20286 2516 0 net20
rlabel metal1 35926 2278 35926 2278 0 net21
rlabel metal1 4278 31790 4278 31790 0 net22
rlabel metal1 42872 47158 42872 47158 0 net23
rlabel metal2 46966 24174 46966 24174 0 net24
rlabel metal3 19941 46988 19941 46988 0 net25
rlabel metal1 4232 15062 4232 15062 0 net26
rlabel metal1 11914 21386 11914 21386 0 net27
rlabel metal1 19964 38862 19964 38862 0 net28
rlabel metal2 7314 3468 7314 3468 0 net29
rlabel metal1 32292 25874 32292 25874 0 net3
rlabel metal2 3082 43486 3082 43486 0 net30
rlabel metal2 19734 3808 19734 3808 0 net31
rlabel metal2 2070 9792 2070 9792 0 net32
rlabel metal2 44942 3264 44942 3264 0 net33
rlabel metal1 2898 3706 2898 3706 0 net34
rlabel metal1 46506 19924 46506 19924 0 net35
rlabel metal1 47196 16014 47196 16014 0 net36
rlabel metal2 46506 36380 46506 36380 0 net37
rlabel metal2 5290 46172 5290 46172 0 net38
rlabel metal2 46506 25500 46506 25500 0 net39
rlabel metal2 31878 26554 31878 26554 0 net4
rlabel metal1 2898 10574 2898 10574 0 net40
rlabel metal1 46874 42738 46874 42738 0 net41
rlabel metal2 29762 46478 29762 46478 0 net42
rlabel metal1 12512 10574 12512 10574 0 net43
rlabel metal1 46506 18836 46506 18836 0 net44
rlabel metal1 1610 4692 1610 4692 0 net45
rlabel metal1 46874 5746 46874 5746 0 net46
rlabel metal1 1610 46036 1610 46036 0 net47
rlabel metal1 44758 4658 44758 4658 0 net48
rlabel metal1 5796 3502 5796 3502 0 net49
rlabel metal2 21666 21760 21666 21760 0 net5
rlabel metal1 47242 12342 47242 12342 0 net50
rlabel metal2 45448 46580 45448 46580 0 net51
rlabel metal2 46506 45696 46506 45696 0 net52
rlabel metal1 32890 46580 32890 46580 0 net53
rlabel metal1 6762 2482 6762 2482 0 net54
rlabel metal1 1748 43282 1748 43282 0 net55
rlabel metal2 46506 29852 46506 29852 0 net56
rlabel metal2 22494 46784 22494 46784 0 net57
rlabel metal2 45402 46308 45402 46308 0 net58
rlabel metal2 4186 20672 4186 20672 0 net59
rlabel metal1 41906 2550 41906 2550 0 net6
rlabel metal2 17342 3468 17342 3468 0 net60
rlabel metal1 1978 14994 1978 14994 0 net61
rlabel metal1 46874 27506 46874 27506 0 net62
rlabel metal2 1886 4352 1886 4352 0 net63
rlabel metal2 2070 7616 2070 7616 0 net64
rlabel metal2 39974 3264 39974 3264 0 net65
rlabel metal2 46506 40732 46506 40732 0 net66
rlabel metal2 2070 41344 2070 41344 0 net67
rlabel metal2 46506 26588 46506 26588 0 net68
rlabel metal1 45402 41140 45402 41140 0 net69
rlabel metal1 18262 33422 18262 33422 0 net7
rlabel metal1 44988 3570 44988 3570 0 net70
rlabel metal1 40158 46002 40158 46002 0 net71
rlabel metal2 32338 3264 32338 3264 0 net72
rlabel metal1 41446 22066 41446 22066 0 net73
rlabel metal2 27186 3468 27186 3468 0 net74
rlabel metal1 36984 46478 36984 46478 0 net75
rlabel metal1 9844 4658 9844 4658 0 net76
rlabel metal2 39790 46784 39790 46784 0 net77
rlabel metal2 16790 3740 16790 3740 0 net78
rlabel metal1 45724 5134 45724 5134 0 net79
rlabel metal1 23230 2482 23230 2482 0 net8
rlabel metal1 1978 6290 1978 6290 0 net80
rlabel metal1 1978 13906 1978 13906 0 net81
rlabel metal1 2162 45356 2162 45356 0 net82
rlabel metal1 47242 6834 47242 6834 0 net83
rlabel metal2 46506 41820 46506 41820 0 net84
rlabel metal1 46506 37162 46506 37162 0 net85
rlabel metal2 15042 46172 15042 46172 0 net86
rlabel metal2 46506 45084 46506 45084 0 net87
rlabel metal2 25990 3740 25990 3740 0 net88
rlabel metal2 39054 5440 39054 5440 0 net89
rlabel metal1 4347 37094 4347 37094 0 net9
rlabel metal1 42044 46546 42044 46546 0 net90
rlabel metal2 24794 3468 24794 3468 0 net91
rlabel metal2 43102 5100 43102 5100 0 net92
rlabel metal2 2162 32640 2162 32640 0 net93
rlabel metal2 46506 16796 46506 16796 0 net94
rlabel metal1 12006 46580 12006 46580 0 net95
rlabel metal1 4002 2516 4002 2516 0 net96
rlabel metal1 10626 3026 10626 3026 0 net97
rlabel metal2 1610 16796 1610 16796 0 net98
rlabel metal1 46874 28594 46874 28594 0 net99
rlabel metal2 46874 24259 46874 24259 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
